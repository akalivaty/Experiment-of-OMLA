//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n445, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n548, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT69), .Z(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(G567), .B2(new_n457), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT70), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT71), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT3), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(G137), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n470), .A2(new_n472), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT72), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n472), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n483), .A2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n490), .A2(G124), .B1(G136), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n484), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(G162));
  AND2_X1   g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n470), .A2(new_n484), .A3(new_n472), .A4(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n472), .A2(new_n477), .A3(G138), .A4(new_n484), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n476), .A2(G2105), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(new_n499), .B1(G102), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(G114), .A2(G2104), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n487), .B2(G126), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n497), .B(new_n501), .C1(new_n504), .C2(new_n484), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT73), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n518), .B(new_n520), .C1(new_n507), .C2(new_n508), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n513), .A2(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(new_n511), .A2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(new_n520), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n528), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n524), .B(new_n526), .C1(new_n527), .C2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n516), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n528), .A2(G543), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT74), .B(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n534), .A2(new_n535), .B1(new_n521), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n516), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT75), .B(G81), .Z(new_n542));
  OAI22_X1  g117(.A1(new_n534), .A2(new_n541), .B1(new_n521), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT76), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n511), .A2(G53), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n514), .A2(G65), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n516), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n521), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n514), .A2(new_n528), .A3(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n556), .B1(new_n560), .B2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n553), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n563));
  XNOR2_X1  g138(.A(G171), .B(new_n563), .ZN(G301));
  OR2_X1    g139(.A1(new_n513), .A2(new_n522), .ZN(G303));
  INV_X1    g140(.A(G74), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n516), .B1(new_n527), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n528), .A2(G49), .A3(G543), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  AOI211_X1 g144(.A(new_n567), .B(new_n569), .C1(new_n560), .C2(G87), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n527), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(new_n511), .B2(G48), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n560), .B2(G86), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  AOI211_X1 g153(.A(KEYINPUT79), .B(new_n578), .C1(new_n558), .C2(new_n559), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n516), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT81), .B(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n534), .A2(new_n585), .B1(new_n521), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n560), .A2(G92), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n527), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n511), .B2(G54), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n560), .A2(new_n597), .A3(G92), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n592), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n590), .B1(G868), .B2(new_n600), .ZN(G284));
  OAI21_X1  g176(.A(new_n590), .B1(G868), .B2(new_n600), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  INV_X1    g183(.A(new_n544), .ZN(new_n609));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n599), .A2(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g189(.A1(new_n478), .A2(new_n464), .A3(G2105), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n490), .A2(G123), .B1(G135), .B2(new_n491), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n484), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2430), .ZN(new_n626));
  INV_X1    g201(.A(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT16), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n633), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n634), .B2(new_n638), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OR3_X1    g217(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT83), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2084), .B(G2090), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT82), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n653), .B(new_n656), .C1(new_n652), .C2(new_n647), .ZN(new_n657));
  OR3_X1    g232(.A1(new_n650), .A2(new_n652), .A3(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n651), .A3(new_n647), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G2096), .ZN(new_n662));
  NAND4_X1  g237(.A1(new_n657), .A2(new_n660), .A3(new_n623), .A4(new_n658), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G2100), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(G2100), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT85), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n676), .B2(new_n677), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n672), .A2(new_n679), .A3(new_n675), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n685), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n686), .B2(new_n689), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n670), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n694), .A2(new_n690), .A3(new_n669), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NAND3_X1  g272(.A1(new_n619), .A2(G29), .A3(new_n621), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT95), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G5), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G171), .B2(new_n701), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(KEYINPUT98), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(KEYINPUT98), .ZN(new_n705));
  OAI21_X1  g280(.A(G1961), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(G16), .A2(G21), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G286), .B2(new_n701), .ZN(new_n708));
  INV_X1    g283(.A(G1966), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G11), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT96), .B(G28), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT30), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n711), .B1(new_n713), .B2(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(new_n709), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT97), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n708), .A2(KEYINPUT97), .A3(new_n709), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n700), .A2(new_n706), .A3(new_n710), .A4(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT99), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n544), .A2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G16), .B2(G19), .ZN(new_n724));
  INV_X1    g299(.A(G1341), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G27), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n727), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2078), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n704), .A2(new_n705), .A3(G1961), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n724), .A2(new_n725), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n701), .A2(G4), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n600), .B2(new_n701), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1348), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n701), .A2(G20), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n604), .B2(new_n701), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1956), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n722), .A2(new_n726), .A3(new_n733), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n727), .A2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n490), .A2(G129), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT92), .Z(new_n746));
  INV_X1    g321(.A(new_n464), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n487), .A2(G141), .B1(G105), .B2(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n746), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n744), .B1(new_n754), .B2(new_n727), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT94), .Z(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n755), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G162), .A2(new_n727), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n727), .B2(G35), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT29), .B(G2090), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n761), .B(new_n762), .Z(new_n763));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n764));
  INV_X1    g339(.A(G26), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G29), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(G29), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n490), .A2(G128), .B1(G140), .B2(new_n491), .ZN(new_n768));
  OR2_X1    g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(G2104), .C1(G116), .C2(new_n484), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n767), .B1(new_n771), .B2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n766), .B1(new_n772), .B2(new_n764), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2067), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(KEYINPUT24), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(KEYINPUT24), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n727), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G160), .B2(new_n727), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G2084), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT91), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n743), .A2(new_n759), .A3(new_n763), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n779), .A2(G2084), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT100), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n490), .A2(G119), .B1(G131), .B2(new_n491), .ZN(new_n786));
  OR2_X1    g361(.A1(G95), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G107), .C2(new_n484), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n727), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G25), .B2(new_n727), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT35), .B(G1991), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n701), .A2(G24), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n588), .B2(new_n701), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1986), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n799));
  INV_X1    g374(.A(new_n575), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n560), .A2(G86), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT79), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n576), .A3(G86), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(new_n581), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G16), .ZN(new_n808));
  NOR2_X1   g383(.A1(G6), .A2(G16), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n799), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n701), .B1(new_n805), .B2(new_n806), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n812), .A2(KEYINPUT32), .A3(new_n809), .ZN(new_n813));
  OAI21_X1  g388(.A(G1981), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n808), .A2(new_n799), .A3(new_n810), .ZN(new_n815));
  INV_X1    g390(.A(G1981), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT32), .B1(new_n812), .B2(new_n809), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT86), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G16), .B2(G23), .ZN(new_n821));
  OR3_X1    g396(.A1(new_n820), .A2(G16), .A3(G23), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n821), .B(new_n822), .C1(G288), .C2(new_n701), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT33), .B(G1976), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(G166), .A2(G16), .ZN(new_n826));
  NOR2_X1   g401(.A1(G16), .A2(G22), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT87), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT87), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G1971), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(G1971), .A3(new_n832), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n825), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n819), .A2(KEYINPUT34), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT34), .B1(new_n819), .B2(new_n837), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n794), .B(new_n798), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n783), .B(new_n785), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n841), .ZN(new_n843));
  NOR2_X1   g418(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n727), .A2(G33), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n491), .A2(G139), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT89), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n491), .A2(KEYINPUT89), .A3(G139), .ZN(new_n851));
  NAND2_X1  g426(.A1(G115), .A2(G2104), .ZN(new_n852));
  INV_X1    g427(.A(G127), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n478), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n850), .A2(new_n851), .B1(G2105), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n500), .A2(G103), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT25), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n847), .B1(new_n858), .B2(G29), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT90), .B(G2072), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n842), .A2(new_n846), .A3(new_n861), .ZN(G311));
  INV_X1    g437(.A(new_n743), .ZN(new_n863));
  INV_X1    g438(.A(new_n759), .ZN(new_n864));
  INV_X1    g439(.A(new_n763), .ZN(new_n865));
  INV_X1    g440(.A(new_n782), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n840), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n843), .ZN(new_n869));
  INV_X1    g444(.A(new_n861), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n840), .A2(new_n845), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n785), .ZN(G150));
  INV_X1    g447(.A(G55), .ZN(new_n873));
  INV_X1    g448(.A(G93), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n534), .A2(new_n873), .B1(new_n521), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n516), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(G860), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT37), .Z(new_n882));
  NOR2_X1   g457(.A1(new_n599), .A2(new_n607), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT38), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT39), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n877), .A2(KEYINPUT103), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n544), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT103), .B1(new_n877), .B2(new_n879), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n544), .A3(new_n886), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n885), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n882), .B1(new_n894), .B2(G860), .ZN(G145));
  XOR2_X1   g470(.A(new_n771), .B(new_n616), .Z(new_n896));
  NAND2_X1  g471(.A1(new_n858), .A2(G164), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n855), .A2(new_n505), .A3(new_n857), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n771), .B(new_n616), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(new_n897), .A3(new_n898), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n490), .A2(G130), .B1(G142), .B2(new_n491), .ZN(new_n903));
  NOR2_X1   g478(.A1(G106), .A2(G2105), .ZN(new_n904));
  OAI21_X1  g479(.A(G2104), .B1(new_n484), .B2(G118), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n790), .B(new_n906), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n900), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n900), .B2(new_n902), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n492), .A2(new_n494), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n914));
  OAI21_X1  g489(.A(G160), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n622), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n917));
  INV_X1    g492(.A(G160), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n912), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n916), .B1(new_n915), .B2(new_n919), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n921), .A2(new_n922), .A3(new_n754), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n915), .A2(new_n919), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n622), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n753), .B1(new_n925), .B2(new_n920), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n910), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n754), .B1(new_n921), .B2(new_n922), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n753), .A3(new_n920), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n928), .B(new_n929), .C1(new_n908), .C2(new_n909), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g508(.A1(new_n600), .A2(new_n604), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n599), .A2(G299), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT41), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(KEYINPUT105), .A3(new_n939), .ZN(new_n940));
  OR3_X1    g515(.A1(new_n936), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n893), .A2(new_n612), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n889), .B(new_n892), .C1(G559), .C2(new_n599), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n936), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(new_n945), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n807), .A2(G288), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n570), .B1(new_n805), .B2(new_n806), .ZN(new_n950));
  OAI21_X1  g525(.A(G166), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  NAND2_X1  g527(.A1(G305), .A2(new_n570), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(G303), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n588), .B(KEYINPUT106), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n951), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n951), .B2(new_n954), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT42), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n951), .A2(new_n954), .ZN(new_n959));
  INV_X1    g534(.A(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n951), .A2(new_n954), .A3(new_n955), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n948), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n948), .B1(new_n958), .B2(new_n964), .ZN(new_n967));
  OAI21_X1  g542(.A(G868), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n880), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(G868), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(G295));
  NAND2_X1  g547(.A1(new_n958), .A2(new_n964), .ZN(new_n973));
  INV_X1    g548(.A(new_n948), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n610), .B1(new_n975), .B2(new_n965), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT107), .B1(new_n976), .B2(new_n970), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n968), .A2(new_n978), .A3(new_n971), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(G331));
  AND2_X1   g555(.A1(G171), .A2(G286), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(G301), .B2(G168), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n887), .A2(new_n888), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n969), .A2(KEYINPUT103), .A3(new_n544), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(G301), .A2(G168), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n889), .B(new_n892), .C1(new_n986), .C2(new_n981), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(new_n941), .A3(new_n940), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n987), .A3(new_n947), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n956), .A2(new_n957), .ZN(new_n992));
  AOI21_X1  g567(.A(G37), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n939), .A2(KEYINPUT108), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n937), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n939), .A2(KEYINPUT108), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n988), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n990), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n985), .A2(new_n987), .A3(KEYINPUT109), .A4(new_n947), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n961), .A2(new_n963), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n993), .A2(KEYINPUT43), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n989), .A2(new_n990), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT43), .B1(new_n993), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT44), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n993), .A2(new_n1009), .A3(new_n1003), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1009), .B1(new_n993), .B2(new_n1006), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1008), .B1(new_n1013), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n505), .A2(new_n1016), .A3(KEYINPUT45), .A4(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n470), .A2(G126), .A3(new_n472), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n484), .B1(new_n1019), .B2(new_n502), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n498), .A2(new_n499), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n500), .A2(G102), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n497), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT45), .B(new_n1017), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT111), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1018), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n480), .A2(G2105), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT110), .B(G40), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n466), .B1(new_n487), .B2(G137), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1027), .B(new_n1029), .C1(new_n1030), .C2(G2105), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1017), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1971), .B1(new_n1026), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(new_n1032), .B2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n505), .A2(new_n1037), .A3(new_n1038), .A4(new_n1017), .ZN(new_n1039));
  INV_X1    g614(.A(G2090), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1038), .B(new_n1017), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT116), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1015), .B1(new_n1035), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n474), .A2(new_n481), .A3(new_n1028), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n1025), .B2(new_n1018), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT117), .B(new_n1043), .C1(new_n1049), .C2(G1971), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1045), .A2(new_n1050), .A3(G8), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052));
  XOR2_X1   g627(.A(new_n1052), .B(KEYINPUT55), .Z(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT114), .B(G1981), .Z(new_n1057));
  OAI211_X1 g632(.A(new_n575), .B(new_n1057), .C1(new_n577), .C2(new_n579), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n514), .A2(new_n528), .A3(G86), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n816), .B1(new_n575), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1056), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT49), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1032), .A2(new_n1031), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1056), .B(new_n1067), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT113), .B1(new_n570), .B2(G1976), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1047), .A2(new_n505), .A3(new_n1017), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(G8), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n570), .A2(G1976), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1073), .A3(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1066), .B(new_n1070), .C1(KEYINPUT52), .C2(new_n1073), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1069), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1083));
  OAI221_X1 g658(.A(new_n1082), .B1(G2090), .B2(new_n1083), .C1(new_n1049), .C2(G1971), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(G2090), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT112), .B1(new_n1035), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1084), .A2(new_n1053), .A3(G8), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1069), .A2(new_n1078), .A3(KEYINPUT118), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1055), .A2(new_n1081), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  INV_X1    g665(.A(G2078), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1024), .A2(KEYINPUT111), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1024), .A2(KEYINPUT111), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1091), .B(new_n1034), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1961), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G40), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1091), .A2(KEYINPUT124), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1091), .A2(KEYINPUT124), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1095), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1100), .A2(G160), .A3(new_n1046), .A4(new_n1103), .ZN(new_n1104));
  AND4_X1   g679(.A1(G301), .A2(new_n1096), .A3(new_n1098), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1097), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1034), .A2(KEYINPUT53), .A3(new_n1091), .A4(new_n1024), .ZN(new_n1107));
  AOI21_X1  g682(.A(G301), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1090), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1096), .A2(new_n1104), .A3(new_n1098), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G171), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1106), .A2(G301), .A3(new_n1107), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(KEYINPUT54), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1046), .A2(new_n1047), .A3(new_n1024), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n709), .ZN(new_n1116));
  INV_X1    g691(.A(G2084), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1036), .A2(new_n1117), .A3(new_n1041), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1065), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT51), .B1(new_n1119), .B2(KEYINPUT123), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1116), .A2(G168), .A3(new_n1118), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(G8), .A3(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1036), .A2(new_n1117), .A3(new_n1041), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1966), .B1(new_n1034), .B2(new_n1024), .ZN(new_n1124));
  OAI21_X1  g699(.A(G286), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(new_n1121), .A3(G8), .ZN(new_n1126));
  OAI21_X1  g701(.A(G8), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(KEYINPUT51), .A3(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1122), .A2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1089), .A2(new_n1114), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G299), .B(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1036), .A2(new_n1042), .A3(new_n1039), .ZN(new_n1135));
  INV_X1    g710(.A(G1956), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1026), .A2(new_n1034), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1134), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1137), .A2(new_n1134), .A3(new_n1139), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n599), .ZN(new_n1142));
  INV_X1    g717(.A(G1348), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1083), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(G2067), .B2(new_n1071), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1140), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1141), .B2(new_n1140), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1137), .A2(new_n1134), .A3(new_n1139), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(KEYINPUT122), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1144), .B(new_n600), .C1(G2067), .C2(new_n1071), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1145), .A2(new_n599), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(KEYINPUT60), .A3(new_n1153), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1150), .B1(new_n1141), .B2(new_n1140), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1152), .A2(new_n1154), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(G1996), .ZN(new_n1164));
  INV_X1    g739(.A(G1996), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1026), .A2(KEYINPUT119), .A3(new_n1165), .A4(new_n1034), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1071), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT120), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1071), .A2(new_n1171), .A3(new_n1168), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n544), .B(new_n1161), .C1(new_n1167), .C2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1161), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1175), .B(new_n1176), .C1(new_n1177), .C2(new_n609), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1146), .B1(new_n1158), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1132), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(G1976), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1069), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1059), .B1(new_n1183), .B2(new_n570), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1066), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1184), .A2(new_n1185), .B1(new_n1087), .B2(new_n1079), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1089), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1122), .A2(new_n1130), .A3(new_n1187), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1190), .A2(new_n1108), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1186), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1127), .A2(G286), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1193), .B1(new_n1089), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1084), .A2(G8), .A3(new_n1086), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1079), .B1(new_n1197), .B2(new_n1054), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1198), .A2(KEYINPUT63), .A3(new_n1087), .A4(new_n1194), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1181), .A2(new_n1192), .A3(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1046), .A2(new_n1031), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n754), .A2(new_n1165), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n789), .A2(new_n793), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n771), .A2(G2067), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n771), .A2(G2067), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n753), .A2(G1996), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1203), .A2(new_n1204), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1209), .B1(new_n793), .B2(new_n789), .ZN(new_n1210));
  INV_X1    g785(.A(G1986), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1210), .B1(new_n1211), .B2(new_n588), .ZN(new_n1212));
  NOR2_X1   g787(.A1(G290), .A2(G1986), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1202), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1201), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1202), .A2(new_n1165), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT46), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1217), .A2(KEYINPUT125), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1216), .B(new_n1218), .ZN(new_n1219));
  AND2_X1   g794(.A1(new_n754), .A2(new_n1207), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1202), .ZN(new_n1221));
  OAI221_X1 g796(.A(new_n1219), .B1(KEYINPUT125), .B2(new_n1217), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT47), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1203), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1205), .B1(new_n1224), .B2(new_n1204), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n1202), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1202), .A2(new_n1213), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1227), .B(KEYINPUT48), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1228), .B1(new_n1210), .B2(new_n1221), .ZN(new_n1229));
  AND3_X1   g804(.A1(new_n1223), .A2(new_n1226), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1215), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1233));
  NAND3_X1  g807(.A1(new_n666), .A2(new_n1233), .A3(new_n462), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n662), .A2(new_n663), .ZN(new_n1235));
  INV_X1    g809(.A(G2100), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g811(.A1(new_n662), .A2(G2100), .A3(new_n663), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n1237), .A2(new_n462), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n1239), .A2(KEYINPUT126), .ZN(new_n1240));
  NAND2_X1  g814(.A1(new_n1234), .A2(new_n1240), .ZN(new_n1241));
  AND3_X1   g815(.A1(new_n693), .A2(new_n695), .A3(new_n645), .ZN(new_n1242));
  AOI21_X1  g816(.A(KEYINPUT127), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g817(.A(new_n1233), .B1(new_n666), .B2(new_n462), .ZN(new_n1244));
  AND4_X1   g818(.A1(new_n1233), .A2(new_n1237), .A3(new_n462), .A4(new_n1238), .ZN(new_n1245));
  OAI211_X1 g819(.A(new_n1242), .B(KEYINPUT127), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g820(.A1(new_n1246), .A2(new_n932), .ZN(new_n1247));
  NAND2_X1  g821(.A1(new_n993), .A2(new_n1006), .ZN(new_n1248));
  NAND2_X1  g822(.A1(new_n1248), .A2(KEYINPUT43), .ZN(new_n1249));
  AOI211_X1 g823(.A(new_n1243), .B(new_n1247), .C1(new_n1249), .C2(new_n1010), .ZN(G308));
  AOI21_X1  g824(.A(new_n1243), .B1(new_n1249), .B2(new_n1010), .ZN(new_n1251));
  NAND3_X1  g825(.A1(new_n1251), .A2(new_n932), .A3(new_n1246), .ZN(G225));
endmodule


