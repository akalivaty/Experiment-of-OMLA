//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT64), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n468), .B1(new_n470), .B2(G101), .ZN(new_n471));
  AND4_X1   g046(.A1(new_n468), .A2(new_n465), .A3(G101), .A4(G2104), .ZN(new_n472));
  OAI22_X1  g047(.A1(new_n466), .A2(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT69), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(G113), .A3(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g060(.A(KEYINPUT70), .B(G2105), .C1(new_n477), .C2(new_n482), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n473), .B1(new_n485), .B2(new_n486), .ZN(G160));
  AND2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(new_n465), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n494));
  INV_X1    g069(.A(G136), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n492), .B(new_n494), .C1(new_n495), .C2(new_n466), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  OAI211_X1 g072(.A(G138), .B(new_n465), .C1(new_n488), .C2(new_n489), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .A4(new_n465), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n510), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n507), .A2(new_n515), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n508), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(KEYINPUT74), .A3(new_n518), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n514), .A2(new_n519), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  XOR2_X1   g108(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n531), .A2(new_n533), .A3(new_n536), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n514), .A2(new_n519), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n529), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n507), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  AND2_X1   g121(.A1(new_n514), .A2(G56), .ZN(new_n547));
  AND2_X1   g122(.A1(G68), .A2(G543), .ZN(new_n548));
  OAI21_X1  g123(.A(G651), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n530), .A2(G43), .B1(new_n532), .B2(G81), .ZN(new_n552));
  OAI211_X1 g127(.A(KEYINPUT76), .B(G651), .C1(new_n547), .C2(new_n548), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(KEYINPUT77), .A2(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n529), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(new_n561), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n527), .A2(new_n563), .A3(new_n528), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n532), .A2(KEYINPUT78), .A3(G91), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n542), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n562), .A2(new_n565), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n514), .A2(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n514), .A2(KEYINPUT79), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g149(.A1(G78), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n570), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  AND2_X1   g153(.A1(new_n523), .A2(new_n524), .ZN(G303));
  NAND2_X1  g154(.A1(new_n530), .A2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n532), .A2(G87), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(new_n511), .A2(new_n513), .ZN(new_n584));
  INV_X1    g159(.A(new_n509), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(G61), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n507), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n512), .B1(KEYINPUT5), .B2(new_n508), .ZN(new_n589));
  NOR3_X1   g164(.A1(new_n510), .A2(KEYINPUT72), .A3(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(G86), .B(new_n585), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G48), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n520), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  XOR2_X1   g170(.A(KEYINPUT80), .B(G47), .Z(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT81), .B(G85), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n529), .A2(new_n596), .B1(new_n542), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n507), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n530), .A2(KEYINPUT82), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n529), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n532), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n542), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n604), .A2(new_n607), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n572), .B2(new_n573), .ZN(new_n614));
  AND2_X1   g189(.A1(G79), .A2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(G651), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n603), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n603), .B1(new_n618), .B2(G868), .ZN(G321));
  MUX2_X1   g195(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g196(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n618), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n464), .A2(new_n470), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  INV_X1    g209(.A(new_n466), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n491), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n465), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n633), .A2(new_n634), .A3(new_n641), .ZN(G156));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT84), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n655), .A2(new_n657), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT17), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n670), .B(new_n667), .C1(new_n663), .C2(new_n665), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n663), .A3(new_n665), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(KEYINPUT87), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT19), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(KEYINPUT87), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  INV_X1    g260(.A(new_n682), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n677), .A2(new_n678), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n686), .A2(new_n679), .A3(new_n688), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n685), .B(new_n689), .C1(new_n686), .C2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  NAND3_X1  g271(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT25), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n464), .A2(G127), .ZN(new_n699));
  NAND2_X1  g274(.A1(G115), .A2(G2104), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n465), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI211_X1 g276(.A(new_n698), .B(new_n701), .C1(G139), .C2(new_n635), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(G33), .ZN(new_n705));
  OR3_X1    g280(.A1(new_n704), .A2(G2072), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(G2072), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n703), .A2(G32), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n635), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT26), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G129), .B2(new_n491), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n708), .B1(new_n714), .B2(new_n703), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT27), .B(G1996), .Z(new_n716));
  OAI211_X1 g291(.A(new_n706), .B(new_n707), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT24), .ZN(new_n718));
  INV_X1    g293(.A(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n718), .B2(new_n719), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G160), .B2(new_n703), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n717), .B1(G2084), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT95), .ZN(new_n724));
  NOR2_X1   g299(.A1(G4), .A2(G16), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n618), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT92), .B(G1348), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n722), .A2(G2084), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT96), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n703), .A2(G26), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n635), .A2(G140), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT94), .Z(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G116), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n491), .B2(G128), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(G29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2067), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G21), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G168), .B2(new_n743), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G1966), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(G1966), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n742), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n743), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n743), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1961), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n703), .A2(G27), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT97), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n505), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT30), .B(G28), .ZN(new_n757));
  OR2_X1    g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  NAND2_X1  g333(.A1(KEYINPUT31), .A2(G11), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n757), .A2(new_n703), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n640), .B2(new_n703), .ZN(new_n761));
  NAND2_X1  g336(.A1(G162), .A2(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G29), .B2(G35), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT29), .B(G2090), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n715), .A2(new_n716), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(new_n764), .C2(new_n765), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n748), .A2(new_n751), .A3(new_n756), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G19), .ZN(new_n770));
  OR3_X1    g345(.A1(new_n770), .A2(KEYINPUT93), .A3(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(KEYINPUT93), .B1(new_n770), .B2(G16), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n771), .B(new_n772), .C1(new_n555), .C2(new_n743), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1341), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n743), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n724), .A2(new_n731), .A3(new_n769), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n743), .A2(G23), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n743), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT33), .B(G1976), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n743), .A2(G22), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n743), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n787), .B1(new_n789), .B2(G1971), .ZN(new_n790));
  NOR2_X1   g365(.A1(G6), .A2(G16), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n594), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  INV_X1    g368(.A(G1981), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n789), .A2(G1971), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n790), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NOR2_X1   g375(.A1(G25), .A2(G29), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n635), .A2(G131), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT88), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  INV_X1    g380(.A(G107), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(G2105), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n491), .B2(G119), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT89), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n802), .B1(new_n810), .B2(new_n703), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n743), .A2(G24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n601), .B2(new_n743), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1986), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n799), .A2(new_n800), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n819), .A2(KEYINPUT90), .A3(KEYINPUT36), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(KEYINPUT90), .B1(new_n819), .B2(KEYINPUT36), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n799), .A2(new_n824), .A3(new_n800), .A4(new_n818), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT91), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n782), .B1(new_n823), .B2(new_n827), .ZN(G311));
  INV_X1    g403(.A(new_n822), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n825), .A2(KEYINPUT91), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(KEYINPUT91), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n820), .ZN(new_n832));
  INV_X1    g407(.A(new_n782), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(G150));
  NOR2_X1   g409(.A1(new_n617), .A2(new_n623), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n529), .A2(new_n837), .B1(new_n838), .B2(new_n542), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n507), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n554), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n842), .A2(new_n553), .A3(new_n551), .A4(new_n552), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n836), .B(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n842), .A2(new_n849), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT100), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(G145));
  NAND2_X1  g431(.A1(new_n491), .A2(G130), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n465), .A2(G118), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(G142), .B2(new_n635), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n630), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n810), .B(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n502), .A2(new_n504), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n501), .A4(new_n500), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n505), .A2(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n863), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n702), .B(new_n713), .ZN(new_n870));
  INV_X1    g445(.A(new_n740), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(G160), .B(KEYINPUT101), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n640), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  INV_X1    g455(.A(new_n878), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n873), .A2(new_n881), .A3(new_n874), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g459(.A(new_n625), .B(new_n846), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n617), .A2(G299), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n612), .A2(new_n570), .A3(new_n576), .A4(new_n616), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT41), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n888), .B2(new_n885), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(G303), .A2(G288), .ZN(new_n898));
  NAND2_X1  g473(.A1(G166), .A2(new_n784), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n601), .B(new_n594), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n896), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n897), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n897), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(G868), .B2(new_n842), .ZN(G295));
  OAI21_X1  g485(.A(new_n909), .B1(G868), .B2(new_n842), .ZN(G331));
  NAND2_X1  g486(.A1(G168), .A2(G301), .ZN(new_n912));
  NAND2_X1  g487(.A1(G286), .A2(G171), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n846), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n912), .A2(new_n844), .A3(new_n845), .A4(new_n913), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n890), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n889), .A2(new_n892), .A3(new_n916), .A4(new_n915), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n905), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n880), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n918), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n905), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n919), .A2(new_n918), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT104), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n903), .A2(new_n904), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n921), .B1(new_n930), .B2(new_n922), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n929), .B(KEYINPUT44), .C1(new_n928), .C2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n925), .B2(new_n905), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n922), .A2(new_n930), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n928), .A4(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n935), .A2(new_n928), .A3(new_n920), .A4(new_n880), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT105), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n936), .B(new_n938), .C1(new_n927), .C2(new_n928), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n932), .B1(new_n942), .B2(new_n943), .ZN(G397));
  INV_X1    g519(.A(new_n473), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n479), .B(new_n481), .C1(new_n490), .C2(new_n474), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT70), .B1(new_n946), .B2(G2105), .ZN(new_n947));
  INV_X1    g522(.A(new_n486), .ZN(new_n948));
  OAI211_X1 g523(.A(G40), .B(new_n945), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n866), .A2(new_n867), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(KEYINPUT107), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(KEYINPUT107), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(G1996), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT46), .Z(new_n959));
  XNOR2_X1  g534(.A(new_n957), .B(KEYINPUT109), .ZN(new_n960));
  INV_X1    g535(.A(G2067), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n740), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n714), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n959), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n959), .B2(new_n964), .ZN(new_n967));
  INV_X1    g542(.A(new_n812), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n810), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n810), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n960), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n962), .B1(new_n972), .B2(new_n714), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n960), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT108), .B1(new_n958), .B2(new_n714), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n958), .A2(KEYINPUT108), .A3(new_n714), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n971), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n957), .A2(G1986), .A3(G290), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT48), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n966), .A2(new_n967), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n974), .B(new_n970), .C1(new_n975), .C2(new_n976), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(G2067), .B2(new_n740), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n960), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT111), .B(G8), .ZN(new_n984));
  NOR2_X1   g559(.A1(G168), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(KEYINPUT51), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n505), .A2(new_n952), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n505), .B2(new_n952), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n990), .A2(new_n949), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G2084), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n951), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(G40), .A3(G160), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1966), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n993), .A2(new_n994), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n986), .B1(new_n999), .B2(new_n984), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n998), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n949), .A2(new_n992), .ZN(new_n1003));
  INV_X1    g578(.A(new_n990), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n994), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1001), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT51), .B1(new_n1006), .B2(new_n985), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n999), .A2(G168), .A3(new_n984), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1000), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT119), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1011), .B(new_n1000), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n523), .A2(G8), .A3(new_n524), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT55), .Z(new_n1016));
  NAND4_X1  g591(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT45), .A4(new_n952), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n950), .A2(new_n1017), .A3(new_n995), .ZN(new_n1018));
  INV_X1    g593(.A(G1971), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G2090), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n993), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1001), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n987), .A2(new_n989), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n505), .A2(new_n991), .A3(new_n952), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(G40), .A3(G160), .A4(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1027), .A2(G2090), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n984), .B1(new_n1028), .B2(new_n1020), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1024), .B1(new_n1016), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n949), .A2(new_n987), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n984), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n784), .A2(G1976), .ZN(new_n1033));
  INV_X1    g608(.A(G1976), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n586), .A2(new_n587), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G651), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n591), .A2(new_n592), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n519), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1043), .A3(new_n794), .ZN(new_n1044));
  OAI21_X1  g619(.A(G1981), .B1(new_n588), .B2(new_n593), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n984), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n949), .B2(new_n987), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n1053));
  AOI211_X1 g628(.A(new_n1053), .B(KEYINPUT49), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1049), .B(KEYINPUT113), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n794), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n588), .A2(new_n593), .A3(G1981), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1051), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1053), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1050), .A2(KEYINPUT112), .A3(new_n1051), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT113), .B1(new_n1062), .B2(new_n1049), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1039), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT115), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1066), .B(new_n1039), .C1(new_n1056), .C2(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1030), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n997), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n755), .A2(KEYINPUT53), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1071));
  INV_X1    g646(.A(G1961), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1069), .A2(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n950), .A2(new_n1017), .A3(new_n755), .A4(new_n995), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G301), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1010), .A2(new_n1079), .A3(new_n1012), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1014), .A2(new_n1068), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1034), .B(new_n784), .C1(new_n1056), .C2(new_n1063), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1048), .B1(new_n1082), .B2(new_n1044), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1064), .A2(KEYINPUT114), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1039), .C1(new_n1056), .C2(new_n1063), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1024), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1083), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n570), .A2(new_n576), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n570), .B2(new_n576), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n950), .A2(new_n1017), .A3(new_n995), .A4(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1027), .A2(KEYINPUT118), .A3(new_n778), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT118), .B1(new_n1027), .B2(new_n778), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1093), .B(new_n1095), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1348), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n949), .A2(G2067), .A3(new_n987), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n618), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1093), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(KEYINPUT61), .A3(new_n1099), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1101), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n617), .C1(new_n993), .C2(G1348), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1102), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n617), .A2(KEYINPUT60), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1112), .A2(KEYINPUT60), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1018), .A2(G1996), .B1(new_n1031), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n555), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1120), .A3(new_n555), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1109), .A2(new_n1115), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT61), .B1(new_n1107), .B2(new_n1099), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1108), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1078), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n993), .B2(G1961), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1071), .A2(KEYINPUT121), .A3(new_n1072), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1128), .A2(new_n1129), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n945), .A2(G40), .A3(new_n483), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n953), .B2(new_n951), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1017), .A2(new_n1070), .ZN(new_n1137));
  NOR4_X1   g712(.A1(new_n1135), .A2(new_n1136), .A3(KEYINPUT123), .A4(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1132), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1137), .B1(new_n1140), .B2(KEYINPUT122), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1141), .B2(new_n1134), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1130), .B(G301), .C1(new_n1138), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1126), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1125), .A2(new_n1146), .A3(new_n1068), .A4(new_n1013), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1130), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G171), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1145), .B1(new_n1077), .B2(G301), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1081), .B(new_n1089), .C1(new_n1147), .C2(new_n1154), .ZN(new_n1155));
  OR3_X1    g730(.A1(new_n999), .A2(G286), .A3(new_n984), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n1068), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1157), .A2(new_n1024), .A3(KEYINPUT63), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT116), .B1(new_n1087), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT116), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1163), .B(new_n1160), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1159), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1158), .B1(new_n1165), .B2(KEYINPUT117), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(new_n1159), .C1(new_n1162), .C2(new_n1164), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1155), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n977), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n601), .B(G1986), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n957), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n983), .B1(new_n1169), .B2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g748(.A1(G227), .A2(new_n462), .ZN(new_n1175));
  XOR2_X1   g749(.A(new_n1175), .B(KEYINPUT126), .Z(new_n1176));
  NOR2_X1   g750(.A1(G229), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g751(.A1(new_n883), .A2(new_n661), .A3(new_n939), .A4(new_n1177), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


