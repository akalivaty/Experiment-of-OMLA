

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771;

  NOR2_X1 U366 ( .A1(n755), .A2(n625), .ZN(n416) );
  OR2_X1 U367 ( .A1(n650), .A2(n624), .ZN(n625) );
  NOR2_X1 U368 ( .A1(n740), .A2(n704), .ZN(n622) );
  AND2_X1 U369 ( .A1(n604), .A2(n344), .ZN(n612) );
  NOR2_X1 U370 ( .A1(n345), .A2(n607), .ZN(n344) );
  INV_X1 U371 ( .A(n605), .ZN(n345) );
  XNOR2_X1 U372 ( .A(n761), .B(G146), .ZN(n507) );
  XNOR2_X1 U373 ( .A(G143), .B(G128), .ZN(n406) );
  INV_X1 U374 ( .A(G125), .ZN(n480) );
  NAND2_X2 U375 ( .A1(n522), .A2(G214), .ZN(n698) );
  NOR2_X2 U376 ( .A1(n596), .A2(n527), .ZN(n528) );
  XNOR2_X1 U377 ( .A(n507), .B(n477), .ZN(n654) );
  XNOR2_X2 U378 ( .A(n476), .B(n474), .ZN(n372) );
  XNOR2_X2 U379 ( .A(n472), .B(n473), .ZN(n761) );
  XNOR2_X2 U380 ( .A(n491), .B(n490), .ZN(n657) );
  XNOR2_X2 U381 ( .A(n518), .B(n461), .ZN(n759) );
  XNOR2_X2 U382 ( .A(n378), .B(n434), .ZN(n562) );
  XNOR2_X2 U383 ( .A(n615), .B(n376), .ZN(n745) );
  XNOR2_X2 U384 ( .A(n523), .B(KEYINPUT82), .ZN(n615) );
  INV_X2 U385 ( .A(KEYINPUT64), .ZN(n471) );
  NOR2_X2 U386 ( .A1(n560), .A2(n411), .ZN(n561) );
  INV_X1 U387 ( .A(G953), .ZN(n762) );
  BUF_X1 U388 ( .A(G113), .Z(n368) );
  XOR2_X1 U389 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n346) );
  XOR2_X1 U390 ( .A(n682), .B(n681), .Z(n347) );
  OR2_X1 U391 ( .A1(n762), .A2(G952), .ZN(n348) );
  XOR2_X1 U392 ( .A(KEYINPUT36), .B(n617), .Z(n349) );
  AND2_X2 U393 ( .A1(n462), .A2(n456), .ZN(n429) );
  NOR2_X2 U394 ( .A1(n577), .A2(n649), .ZN(n578) );
  INV_X2 U395 ( .A(n600), .ZN(n748) );
  INV_X1 U396 ( .A(G902), .ZN(n554) );
  INV_X1 U397 ( .A(G110), .ZN(n474) );
  XNOR2_X1 U398 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n514) );
  XNOR2_X1 U399 ( .A(G143), .B(G128), .ZN(n515) );
  NOR2_X1 U400 ( .A1(n443), .A2(n441), .ZN(n440) );
  AND2_X1 U401 ( .A1(n442), .A2(KEYINPUT39), .ZN(n441) );
  BUF_X1 U402 ( .A(n657), .Z(n658) );
  BUF_X1 U403 ( .A(n759), .Z(n403) );
  INV_X1 U404 ( .A(n552), .ZN(n472) );
  XNOR2_X1 U405 ( .A(n371), .B(n402), .ZN(n370) );
  XNOR2_X1 U406 ( .A(n515), .B(n514), .ZN(n371) );
  XNOR2_X1 U407 ( .A(n375), .B(G140), .ZN(n531) );
  INV_X1 U408 ( .A(KEYINPUT90), .ZN(n386) );
  INV_X1 U409 ( .A(G131), .ZN(n375) );
  INV_X1 U410 ( .A(KEYINPUT19), .ZN(n376) );
  INV_X1 U411 ( .A(KEYINPUT124), .ZN(n354) );
  BUF_X1 U412 ( .A(G119), .Z(n431) );
  INV_X1 U413 ( .A(KEYINPUT56), .ZN(n351) );
  NOR2_X1 U414 ( .A1(n771), .A2(n770), .ZN(n418) );
  NAND2_X1 U415 ( .A1(n440), .A2(n438), .ZN(n412) );
  NOR2_X1 U416 ( .A1(n720), .A2(n455), .ZN(n564) );
  AND2_X1 U417 ( .A1(n447), .A2(n446), .ZN(n445) );
  INV_X1 U418 ( .A(n676), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n556), .B(n555), .ZN(n570) );
  XNOR2_X1 U420 ( .A(n669), .B(n369), .ZN(n687) );
  XNOR2_X1 U421 ( .A(n675), .B(KEYINPUT123), .ZN(n676) );
  XNOR2_X1 U422 ( .A(n519), .B(n370), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n531), .B(n435), .ZN(n758) );
  XNOR2_X1 U424 ( .A(G107), .B(G104), .ZN(n475) );
  XNOR2_X1 U425 ( .A(G902), .B(KEYINPUT84), .ZN(n492) );
  XNOR2_X1 U426 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n461) );
  XNOR2_X1 U427 ( .A(G101), .B(G131), .ZN(n503) );
  XNOR2_X1 U428 ( .A(G128), .B(G137), .ZN(n481) );
  BUF_X1 U429 ( .A(KEYINPUT125), .Z(n660) );
  INV_X2 U430 ( .A(n679), .ZN(n684) );
  XNOR2_X1 U431 ( .A(n350), .B(n660), .ZN(G66) );
  NAND2_X1 U432 ( .A1(n367), .A2(n348), .ZN(n350) );
  XNOR2_X1 U433 ( .A(n352), .B(n351), .ZN(G51) );
  NAND2_X1 U434 ( .A1(n365), .A2(n348), .ZN(n352) );
  NAND2_X1 U435 ( .A1(n353), .A2(n348), .ZN(n358) );
  XNOR2_X1 U436 ( .A(n683), .B(n347), .ZN(n353) );
  XNOR2_X1 U437 ( .A(n355), .B(n354), .ZN(G63) );
  NAND2_X1 U438 ( .A1(n363), .A2(n348), .ZN(n355) );
  XNOR2_X1 U439 ( .A(n356), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U440 ( .A1(n361), .A2(n348), .ZN(n356) );
  XNOR2_X1 U441 ( .A(n357), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U442 ( .A1(n359), .A2(n348), .ZN(n357) );
  XNOR2_X1 U443 ( .A(n358), .B(n346), .ZN(G60) );
  XNOR2_X1 U444 ( .A(n645), .B(n360), .ZN(n359) );
  INV_X1 U445 ( .A(n644), .ZN(n360) );
  XNOR2_X1 U446 ( .A(n656), .B(n362), .ZN(n361) );
  INV_X1 U447 ( .A(n655), .ZN(n362) );
  XNOR2_X1 U448 ( .A(n677), .B(n364), .ZN(n363) );
  BUF_X1 U449 ( .A(n582), .Z(n430) );
  XNOR2_X1 U450 ( .A(n689), .B(n366), .ZN(n365) );
  INV_X1 U451 ( .A(n688), .ZN(n366) );
  XNOR2_X1 U452 ( .A(n659), .B(n658), .ZN(n367) );
  XNOR2_X1 U453 ( .A(n530), .B(n529), .ZN(n421) );
  NAND2_X1 U454 ( .A1(n421), .A2(n619), .ZN(n557) );
  XNOR2_X2 U455 ( .A(n373), .B(n513), .ZN(n669) );
  XNOR2_X2 U456 ( .A(n372), .B(n475), .ZN(n513) );
  XNOR2_X2 U457 ( .A(n420), .B(n374), .ZN(n373) );
  XNOR2_X1 U458 ( .A(n512), .B(G122), .ZN(n374) );
  XNOR2_X2 U459 ( .A(n466), .B(n465), .ZN(n420) );
  XNOR2_X2 U460 ( .A(n377), .B(KEYINPUT33), .ZN(n459) );
  NAND2_X1 U461 ( .A1(n562), .A2(n511), .ZN(n377) );
  NOR2_X2 U462 ( .A1(n711), .A2(n712), .ZN(n378) );
  XNOR2_X2 U463 ( .A(n576), .B(KEYINPUT107), .ZN(n649) );
  NAND2_X1 U464 ( .A1(n582), .A2(n468), .ZN(n379) );
  NAND2_X1 U465 ( .A1(n582), .A2(n468), .ZN(n581) );
  BUF_X1 U466 ( .A(n654), .Z(n380) );
  XNOR2_X1 U467 ( .A(n467), .B(KEYINPUT0), .ZN(n381) );
  XNOR2_X1 U468 ( .A(n467), .B(KEYINPUT0), .ZN(n457) );
  XNOR2_X1 U469 ( .A(n758), .B(n382), .ZN(n419) );
  NAND2_X1 U470 ( .A1(G227), .A2(n762), .ZN(n382) );
  XNOR2_X1 U471 ( .A(n507), .B(n449), .ZN(n643) );
  XNOR2_X1 U472 ( .A(n609), .B(n479), .ZN(n711) );
  BUF_X1 U473 ( .A(n711), .Z(n424) );
  XNOR2_X1 U474 ( .A(n453), .B(n452), .ZN(n451) );
  NAND2_X1 U475 ( .A1(n451), .A2(n389), .ZN(n450) );
  XNOR2_X1 U476 ( .A(n379), .B(KEYINPUT32), .ZN(n383) );
  XNOR2_X1 U477 ( .A(n450), .B(KEYINPUT45), .ZN(n384) );
  XNOR2_X1 U478 ( .A(n581), .B(KEYINPUT32), .ZN(n661) );
  XNOR2_X1 U479 ( .A(n450), .B(KEYINPUT45), .ZN(n662) );
  INV_X1 U480 ( .A(n679), .ZN(n385) );
  NAND2_X2 U481 ( .A1(n642), .A2(n695), .ZN(n679) );
  XNOR2_X1 U482 ( .A(n386), .B(n497), .ZN(n498) );
  BUF_X1 U483 ( .A(n687), .Z(n387) );
  XNOR2_X2 U484 ( .A(n408), .B(n409), .ZN(n598) );
  XNOR2_X1 U485 ( .A(n454), .B(KEYINPUT110), .ZN(n592) );
  INV_X1 U486 ( .A(KEYINPUT65), .ZN(n463) );
  INV_X1 U487 ( .A(KEYINPUT88), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n460), .B(n485), .ZN(n486) );
  XNOR2_X1 U489 ( .A(n759), .B(KEYINPUT75), .ZN(n460) );
  XOR2_X1 U490 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n483) );
  XNOR2_X1 U491 ( .A(n508), .B(G472), .ZN(n716) );
  XOR2_X1 U492 ( .A(G107), .B(G122), .Z(n551) );
  INV_X1 U493 ( .A(KEYINPUT9), .ZN(n428) );
  OR2_X1 U494 ( .A1(n571), .A2(n565), .ZN(n600) );
  INV_X1 U495 ( .A(KEYINPUT80), .ZN(n452) );
  XOR2_X1 U496 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n494) );
  XOR2_X1 U497 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n504) );
  XNOR2_X1 U498 ( .A(n368), .B(G143), .ZN(n536) );
  XNOR2_X1 U499 ( .A(G104), .B(G122), .ZN(n532) );
  NAND2_X1 U500 ( .A1(n401), .A2(KEYINPUT86), .ZN(n400) );
  INV_X1 U501 ( .A(G224), .ZN(n401) );
  NAND2_X1 U502 ( .A1(KEYINPUT86), .A2(G953), .ZN(n399) );
  NAND2_X1 U503 ( .A1(G237), .A2(G234), .ZN(n524) );
  NOR2_X1 U504 ( .A1(n614), .A2(n613), .ZN(n626) );
  INV_X1 U505 ( .A(KEYINPUT71), .ZN(n434) );
  XNOR2_X1 U506 ( .A(G110), .B(n431), .ZN(n488) );
  NAND2_X1 U507 ( .A1(n398), .A2(n397), .ZN(n517) );
  NAND2_X1 U508 ( .A1(n396), .A2(G224), .ZN(n397) );
  AND2_X1 U509 ( .A1(n400), .A2(n399), .ZN(n398) );
  NOR2_X1 U510 ( .A1(KEYINPUT86), .A2(G953), .ZN(n396) );
  XNOR2_X1 U511 ( .A(n546), .B(n545), .ZN(n571) );
  XNOR2_X1 U512 ( .A(n544), .B(n678), .ZN(n545) );
  BUF_X1 U513 ( .A(n716), .Z(n411) );
  XNOR2_X1 U514 ( .A(n559), .B(KEYINPUT93), .ZN(n454) );
  XOR2_X1 U515 ( .A(KEYINPUT62), .B(n643), .Z(n644) );
  INV_X1 U516 ( .A(n765), .ZN(n437) );
  XNOR2_X1 U517 ( .A(n550), .B(n427), .ZN(n675) );
  XNOR2_X1 U518 ( .A(n553), .B(n428), .ZN(n427) );
  XOR2_X1 U519 ( .A(G116), .B(KEYINPUT7), .Z(n549) );
  INV_X1 U520 ( .A(n729), .ZN(n458) );
  XNOR2_X1 U521 ( .A(n422), .B(n601), .ZN(n771) );
  AND2_X1 U522 ( .A1(n580), .A2(n614), .ZN(n468) );
  AND2_X1 U523 ( .A1(n413), .A2(n693), .ZN(n388) );
  XOR2_X1 U524 ( .A(n588), .B(KEYINPUT69), .Z(n389) );
  OR2_X1 U525 ( .A1(n706), .A2(n705), .ZN(n390) );
  AND2_X1 U526 ( .A1(n430), .A2(n614), .ZN(n391) );
  AND2_X1 U527 ( .A1(n444), .A2(n439), .ZN(n392) );
  INV_X1 U528 ( .A(n663), .ZN(n426) );
  AND2_X1 U529 ( .A1(n424), .A2(n584), .ZN(n393) );
  NOR2_X1 U530 ( .A1(n701), .A2(n707), .ZN(n394) );
  NOR2_X1 U531 ( .A1(n607), .A2(n448), .ZN(n395) );
  XNOR2_X1 U532 ( .A(n471), .B(KEYINPUT4), .ZN(n402) );
  XNOR2_X1 U533 ( .A(n494), .B(n493), .ZN(n404) );
  BUF_X1 U534 ( .A(n381), .Z(n405) );
  XNOR2_X1 U535 ( .A(n380), .B(n653), .ZN(n655) );
  BUF_X1 U536 ( .A(n413), .Z(n407) );
  NOR2_X2 U537 ( .A1(n687), .A2(n636), .ZN(n408) );
  NAND2_X1 U538 ( .A1(n522), .A2(G210), .ZN(n409) );
  NAND2_X1 U539 ( .A1(n383), .A2(n647), .ZN(n410) );
  NAND2_X1 U540 ( .A1(n661), .A2(n647), .ZN(n585) );
  BUF_X1 U541 ( .A(n745), .Z(n432) );
  NAND2_X1 U542 ( .A1(n412), .A2(n748), .ZN(n422) );
  AND2_X1 U543 ( .A1(n412), .A2(n752), .ZN(n757) );
  NAND2_X1 U544 ( .A1(n413), .A2(n663), .ZN(n691) );
  NAND2_X1 U545 ( .A1(n635), .A2(n413), .ZN(n638) );
  XNOR2_X1 U546 ( .A(n407), .B(n437), .ZN(n763) );
  XNOR2_X2 U547 ( .A(n639), .B(KEYINPUT79), .ZN(n413) );
  XNOR2_X1 U548 ( .A(n414), .B(n436), .ZN(n634) );
  NAND2_X1 U549 ( .A1(n415), .A2(n417), .ZN(n414) );
  XNOR2_X1 U550 ( .A(n416), .B(KEYINPUT68), .ZN(n415) );
  XNOR2_X1 U551 ( .A(n418), .B(KEYINPUT46), .ZN(n417) );
  XNOR2_X1 U552 ( .A(n419), .B(n513), .ZN(n477) );
  XNOR2_X1 U553 ( .A(n420), .B(n506), .ZN(n449) );
  NAND2_X1 U554 ( .A1(n652), .A2(KEYINPUT44), .ZN(n456) );
  NOR2_X1 U555 ( .A1(n445), .A2(n599), .ZN(n443) );
  NAND2_X2 U556 ( .A1(n430), .A2(n393), .ZN(n647) );
  NAND2_X1 U557 ( .A1(n423), .A2(n395), .ZN(n444) );
  INV_X1 U558 ( .A(n597), .ZN(n423) );
  NAND2_X1 U559 ( .A1(n592), .A2(n591), .ZN(n597) );
  NAND2_X1 U560 ( .A1(n694), .A2(n425), .ZN(n696) );
  NAND2_X1 U561 ( .A1(n388), .A2(n426), .ZN(n425) );
  NAND2_X1 U562 ( .A1(n585), .A2(KEYINPUT44), .ZN(n464) );
  NAND2_X1 U563 ( .A1(n429), .A2(n578), .ZN(n453) );
  XNOR2_X2 U564 ( .A(n641), .B(KEYINPUT72), .ZN(n695) );
  XNOR2_X1 U565 ( .A(n464), .B(n463), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n433), .B(KEYINPUT94), .ZN(n560) );
  NAND2_X1 U567 ( .A1(n381), .A2(n454), .ZN(n433) );
  INV_X1 U568 ( .A(KEYINPUT48), .ZN(n436) );
  NAND2_X1 U569 ( .A1(n445), .A2(n444), .ZN(n618) );
  NAND2_X1 U570 ( .A1(n445), .A2(n392), .ZN(n438) );
  NOR2_X1 U571 ( .A1(n602), .A2(KEYINPUT39), .ZN(n439) );
  NAND2_X1 U572 ( .A1(n444), .A2(n699), .ZN(n442) );
  NAND2_X1 U573 ( .A1(n607), .A2(n448), .ZN(n446) );
  NAND2_X1 U574 ( .A1(n597), .A2(n448), .ZN(n447) );
  INV_X1 U575 ( .A(KEYINPUT73), .ZN(n448) );
  NOR2_X2 U576 ( .A1(n424), .A2(n349), .ZN(n755) );
  NAND2_X1 U577 ( .A1(n457), .A2(n394), .ZN(n573) );
  INV_X1 U578 ( .A(n405), .ZN(n455) );
  XNOR2_X2 U579 ( .A(n557), .B(KEYINPUT35), .ZN(n652) );
  NAND2_X1 U580 ( .A1(n459), .A2(n405), .ZN(n530) );
  AND2_X1 U581 ( .A1(n459), .A2(n390), .ZN(n725) );
  NAND2_X1 U582 ( .A1(n459), .A2(n458), .ZN(n730) );
  XNOR2_X2 U583 ( .A(G119), .B(KEYINPUT3), .ZN(n465) );
  XNOR2_X2 U584 ( .A(G116), .B(G113), .ZN(n466) );
  NOR2_X2 U585 ( .A1(n745), .A2(n528), .ZN(n467) );
  NAND2_X1 U586 ( .A1(n391), .A2(n575), .ZN(n576) );
  BUF_X1 U587 ( .A(n598), .Z(n631) );
  AND2_X1 U588 ( .A1(n533), .A2(G210), .ZN(n469) );
  AND2_X1 U589 ( .A1(n533), .A2(G214), .ZN(n470) );
  XNOR2_X1 U590 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U591 ( .A(n505), .B(n469), .ZN(n506) );
  XNOR2_X1 U592 ( .A(n534), .B(n470), .ZN(n535) );
  INV_X1 U593 ( .A(KEYINPUT34), .ZN(n529) );
  INV_X1 U594 ( .A(KEYINPUT39), .ZN(n599) );
  XNOR2_X1 U595 ( .A(n471), .B(KEYINPUT4), .ZN(n516) );
  XNOR2_X1 U596 ( .A(G137), .B(n516), .ZN(n473) );
  XNOR2_X1 U597 ( .A(n406), .B(G134), .ZN(n552) );
  XNOR2_X2 U598 ( .A(G101), .B(KEYINPUT85), .ZN(n476) );
  NAND2_X1 U599 ( .A1(n654), .A2(n554), .ZN(n478) );
  XNOR2_X2 U600 ( .A(n478), .B(G469), .ZN(n609) );
  INV_X1 U601 ( .A(KEYINPUT1), .ZN(n479) );
  XNOR2_X2 U602 ( .A(n480), .B(G146), .ZN(n518) );
  XOR2_X1 U603 ( .A(KEYINPUT89), .B(G140), .Z(n482) );
  XNOR2_X1 U604 ( .A(n482), .B(n481), .ZN(n484) );
  INV_X1 U605 ( .A(n486), .ZN(n491) );
  NAND2_X1 U606 ( .A1(G234), .A2(n762), .ZN(n487) );
  XOR2_X1 U607 ( .A(KEYINPUT8), .B(n487), .Z(n547) );
  NAND2_X1 U608 ( .A1(n547), .A2(G221), .ZN(n489) );
  XNOR2_X1 U609 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U610 ( .A1(n657), .A2(n554), .ZN(n499) );
  XOR2_X1 U611 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n496) );
  XNOR2_X1 U612 ( .A(n492), .B(KEYINPUT15), .ZN(n520) );
  NAND2_X1 U613 ( .A1(n520), .A2(G234), .ZN(n493) );
  XNOR2_X1 U614 ( .A(n494), .B(n493), .ZN(n500) );
  NAND2_X1 U615 ( .A1(n500), .A2(G217), .ZN(n495) );
  XNOR2_X1 U616 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U617 ( .A(n499), .B(n498), .ZN(n574) );
  NAND2_X1 U618 ( .A1(n404), .A2(G221), .ZN(n502) );
  XNOR2_X1 U619 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n501) );
  XNOR2_X1 U620 ( .A(n502), .B(n501), .ZN(n707) );
  OR2_X1 U621 ( .A1(n574), .A2(n707), .ZN(n712) );
  XNOR2_X1 U622 ( .A(n504), .B(n503), .ZN(n505) );
  NOR2_X1 U623 ( .A1(G953), .A2(G237), .ZN(n533) );
  NAND2_X1 U624 ( .A1(n643), .A2(n554), .ZN(n508) );
  INV_X1 U625 ( .A(KEYINPUT105), .ZN(n509) );
  XNOR2_X1 U626 ( .A(n509), .B(KEYINPUT6), .ZN(n510) );
  XNOR2_X1 U627 ( .A(n716), .B(n510), .ZN(n614) );
  INV_X1 U628 ( .A(n614), .ZN(n511) );
  XNOR2_X2 U629 ( .A(KEYINPUT70), .B(KEYINPUT16), .ZN(n512) );
  XNOR2_X1 U630 ( .A(n518), .B(n517), .ZN(n519) );
  INV_X1 U631 ( .A(n520), .ZN(n636) );
  INV_X1 U632 ( .A(G237), .ZN(n521) );
  NAND2_X1 U633 ( .A1(n554), .A2(n521), .ZN(n522) );
  NAND2_X1 U634 ( .A1(n598), .A2(n698), .ZN(n523) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n525) );
  XNOR2_X1 U636 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U637 ( .A1(G952), .A2(n526), .ZN(n727) );
  NOR2_X1 U638 ( .A1(n727), .A2(G953), .ZN(n596) );
  NAND2_X1 U639 ( .A1(G902), .A2(n526), .ZN(n593) );
  INV_X1 U640 ( .A(G898), .ZN(n666) );
  NAND2_X1 U641 ( .A1(G953), .A2(n666), .ZN(n671) );
  NOR2_X1 U642 ( .A1(n593), .A2(n671), .ZN(n527) );
  XNOR2_X1 U643 ( .A(n531), .B(n532), .ZN(n534) );
  XNOR2_X1 U644 ( .A(n403), .B(n535), .ZN(n543) );
  XOR2_X1 U645 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n537) );
  XNOR2_X1 U646 ( .A(n537), .B(n536), .ZN(n541) );
  XOR2_X1 U647 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n539) );
  XNOR2_X1 U648 ( .A(KEYINPUT11), .B(KEYINPUT101), .ZN(n538) );
  XNOR2_X1 U649 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U650 ( .A(n541), .B(n540), .Z(n542) );
  XNOR2_X1 U651 ( .A(n543), .B(n542), .ZN(n682) );
  NOR2_X1 U652 ( .A1(G902), .A2(n682), .ZN(n546) );
  XNOR2_X1 U653 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n544) );
  INV_X1 U654 ( .A(G475), .ZN(n678) );
  NAND2_X1 U655 ( .A1(G217), .A2(n547), .ZN(n548) );
  XNOR2_X1 U656 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U657 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U658 ( .A1(n675), .A2(n554), .ZN(n556) );
  XNOR2_X1 U659 ( .A(KEYINPUT103), .B(G478), .ZN(n555) );
  NOR2_X1 U660 ( .A1(n571), .A2(n570), .ZN(n619) );
  NOR2_X1 U661 ( .A1(n574), .A2(n707), .ZN(n558) );
  NAND2_X1 U662 ( .A1(n558), .A2(n609), .ZN(n559) );
  XNOR2_X1 U663 ( .A(n561), .B(KEYINPUT96), .ZN(n736) );
  NAND2_X1 U664 ( .A1(n562), .A2(n411), .ZN(n720) );
  XNOR2_X1 U665 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n563) );
  XNOR2_X1 U666 ( .A(n564), .B(n563), .ZN(n753) );
  NOR2_X1 U667 ( .A1(n736), .A2(n753), .ZN(n569) );
  INV_X1 U668 ( .A(n570), .ZN(n565) );
  AND2_X1 U669 ( .A1(n571), .A2(n565), .ZN(n752) );
  INV_X1 U670 ( .A(n752), .ZN(n566) );
  NAND2_X1 U671 ( .A1(n566), .A2(n600), .ZN(n568) );
  INV_X1 U672 ( .A(KEYINPUT104), .ZN(n567) );
  XNOR2_X1 U673 ( .A(n568), .B(n567), .ZN(n704) );
  NOR2_X1 U674 ( .A1(n569), .A2(n704), .ZN(n577) );
  NAND2_X1 U675 ( .A1(n571), .A2(n570), .ZN(n701) );
  INV_X1 U676 ( .A(KEYINPUT22), .ZN(n572) );
  XNOR2_X2 U677 ( .A(n573), .B(n572), .ZN(n582) );
  INV_X1 U678 ( .A(n424), .ZN(n579) );
  BUF_X1 U679 ( .A(n574), .Z(n604) );
  XNOR2_X1 U680 ( .A(n604), .B(KEYINPUT106), .ZN(n708) );
  NOR2_X1 U681 ( .A1(n579), .A2(n708), .ZN(n575) );
  AND2_X1 U682 ( .A1(n579), .A2(n708), .ZN(n580) );
  INV_X1 U683 ( .A(n604), .ZN(n583) );
  NOR2_X1 U684 ( .A1(n411), .A2(n583), .ZN(n584) );
  NOR2_X1 U685 ( .A1(n652), .A2(KEYINPUT44), .ZN(n587) );
  XNOR2_X1 U686 ( .A(n410), .B(KEYINPUT81), .ZN(n586) );
  NAND2_X1 U687 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U688 ( .A1(n662), .A2(n636), .ZN(n589) );
  XNOR2_X1 U689 ( .A(n589), .B(KEYINPUT77), .ZN(n635) );
  XNOR2_X1 U690 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n601) );
  NAND2_X1 U691 ( .A1(n716), .A2(n698), .ZN(n590) );
  XOR2_X1 U692 ( .A(KEYINPUT30), .B(n590), .Z(n591) );
  OR2_X1 U693 ( .A1(n762), .A2(n593), .ZN(n594) );
  NOR2_X1 U694 ( .A1(G900), .A2(n594), .ZN(n595) );
  NOR2_X1 U695 ( .A1(n596), .A2(n595), .ZN(n607) );
  XNOR2_X1 U696 ( .A(n631), .B(KEYINPUT38), .ZN(n602) );
  INV_X1 U697 ( .A(n602), .ZN(n699) );
  NAND2_X1 U698 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U699 ( .A1(n703), .A2(n701), .ZN(n603) );
  XNOR2_X1 U700 ( .A(KEYINPUT41), .B(n603), .ZN(n729) );
  INV_X1 U701 ( .A(n707), .ZN(n605) );
  AND2_X1 U702 ( .A1(n411), .A2(n612), .ZN(n608) );
  XNOR2_X1 U703 ( .A(KEYINPUT28), .B(n608), .ZN(n610) );
  NAND2_X1 U704 ( .A1(n610), .A2(n609), .ZN(n740) );
  NOR2_X1 U705 ( .A1(n729), .A2(n740), .ZN(n611) );
  XNOR2_X1 U706 ( .A(n611), .B(KEYINPUT42), .ZN(n770) );
  NAND2_X1 U707 ( .A1(n748), .A2(n612), .ZN(n613) );
  XOR2_X1 U708 ( .A(n626), .B(KEYINPUT112), .Z(n616) );
  NOR2_X1 U709 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U710 ( .A1(n619), .A2(n631), .ZN(n620) );
  NOR2_X1 U711 ( .A1(n618), .A2(n620), .ZN(n650) );
  INV_X1 U712 ( .A(n432), .ZN(n621) );
  NAND2_X1 U713 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U714 ( .A(n623), .B(KEYINPUT47), .ZN(n624) );
  XOR2_X1 U715 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n630) );
  NAND2_X1 U716 ( .A1(n626), .A2(n698), .ZN(n627) );
  XOR2_X1 U717 ( .A(KEYINPUT108), .B(n627), .Z(n628) );
  NAND2_X1 U718 ( .A1(n628), .A2(n424), .ZN(n629) );
  XOR2_X1 U719 ( .A(n630), .B(n629), .Z(n632) );
  NOR2_X1 U720 ( .A1(n632), .A2(n631), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n757), .A2(n651), .ZN(n633) );
  NAND2_X1 U722 ( .A1(n634), .A2(n633), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n636), .A2(KEYINPUT2), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n642) );
  INV_X1 U725 ( .A(KEYINPUT2), .ZN(n690) );
  NOR2_X1 U726 ( .A1(n639), .A2(n690), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n640), .A2(n384), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n385), .A2(G472), .ZN(n645) );
  XOR2_X1 U729 ( .A(G110), .B(KEYINPUT113), .Z(n646) );
  XNOR2_X1 U730 ( .A(n647), .B(n646), .ZN(G12) );
  NAND2_X1 U731 ( .A1(n736), .A2(n748), .ZN(n648) );
  XNOR2_X1 U732 ( .A(n648), .B(G104), .ZN(G6) );
  XOR2_X1 U733 ( .A(G101), .B(n649), .Z(G3) );
  XOR2_X1 U734 ( .A(G143), .B(n650), .Z(G45) );
  XOR2_X1 U735 ( .A(n651), .B(G140), .Z(G42) );
  XOR2_X1 U736 ( .A(n652), .B(G122), .Z(G24) );
  NAND2_X1 U737 ( .A1(n684), .A2(G469), .ZN(n656) );
  XNOR2_X1 U738 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n653) );
  NAND2_X1 U739 ( .A1(n684), .A2(G217), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n383), .B(n431), .ZN(G21) );
  BUF_X1 U741 ( .A(n384), .Z(n663) );
  NOR2_X1 U742 ( .A1(n426), .A2(G953), .ZN(n668) );
  NAND2_X1 U743 ( .A1(G953), .A2(G224), .ZN(n664) );
  XOR2_X1 U744 ( .A(KEYINPUT61), .B(n664), .Z(n665) );
  NOR2_X1 U745 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n674) );
  BUF_X1 U747 ( .A(n669), .Z(n670) );
  INV_X1 U748 ( .A(n670), .ZN(n672) );
  NAND2_X1 U749 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U750 ( .A(n674), .B(n673), .ZN(G69) );
  NAND2_X1 U751 ( .A1(n684), .A2(G478), .ZN(n677) );
  NOR2_X1 U752 ( .A1(n679), .A2(n678), .ZN(n683) );
  XNOR2_X1 U753 ( .A(KEYINPUT66), .B(KEYINPUT83), .ZN(n680) );
  XOR2_X1 U754 ( .A(n680), .B(KEYINPUT59), .Z(n681) );
  NAND2_X1 U755 ( .A1(n385), .A2(G210), .ZN(n689) );
  XOR2_X1 U756 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n685) );
  XNOR2_X1 U757 ( .A(n685), .B(KEYINPUT55), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n387), .B(n686), .ZN(n688) );
  NAND2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n692), .A2(KEYINPUT76), .ZN(n694) );
  NOR2_X1 U761 ( .A1(KEYINPUT2), .A2(KEYINPUT76), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U763 ( .A(n697), .B(KEYINPUT78), .ZN(n734) );
  NOR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U766 ( .A(KEYINPUT119), .B(n702), .Z(n706) );
  NOR2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U768 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n710) );
  NAND2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U770 ( .A(n710), .B(n709), .ZN(n718) );
  NAND2_X1 U771 ( .A1(n712), .A2(n424), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT117), .ZN(n714) );
  XNOR2_X1 U773 ( .A(KEYINPUT50), .B(n714), .ZN(n715) );
  NOR2_X1 U774 ( .A1(n411), .A2(n715), .ZN(n717) );
  NAND2_X1 U775 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U777 ( .A(KEYINPUT51), .B(n721), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n729), .A2(n722), .ZN(n723) );
  XNOR2_X1 U779 ( .A(n723), .B(KEYINPUT118), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U781 ( .A(n726), .B(KEYINPUT52), .ZN(n728) );
  NOR2_X1 U782 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U783 ( .A1(n730), .A2(n762), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U786 ( .A(KEYINPUT53), .B(n735), .Z(G75) );
  NAND2_X1 U787 ( .A1(n736), .A2(n752), .ZN(n738) );
  XOR2_X1 U788 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n737) );
  XNOR2_X1 U789 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U790 ( .A(G107), .B(n739), .ZN(G9) );
  INV_X1 U791 ( .A(n740), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(n752), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n741), .A2(n432), .ZN(n743) );
  XNOR2_X1 U794 ( .A(G128), .B(KEYINPUT29), .ZN(n742) );
  XNOR2_X1 U795 ( .A(n743), .B(n742), .ZN(G30) );
  NAND2_X1 U796 ( .A1(n744), .A2(n748), .ZN(n746) );
  NOR2_X1 U797 ( .A1(n746), .A2(n432), .ZN(n747) );
  XOR2_X1 U798 ( .A(G146), .B(n747), .Z(G48) );
  XOR2_X1 U799 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n750) );
  NAND2_X1 U800 ( .A1(n753), .A2(n748), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U802 ( .A(n368), .B(n751), .ZN(G15) );
  NAND2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U804 ( .A(n754), .B(G116), .ZN(G18) );
  XNOR2_X1 U805 ( .A(G125), .B(n755), .ZN(n756) );
  XNOR2_X1 U806 ( .A(n756), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U807 ( .A(G134), .B(n757), .Z(G36) );
  XOR2_X1 U808 ( .A(n758), .B(n403), .Z(n760) );
  XNOR2_X1 U809 ( .A(n761), .B(n760), .ZN(n765) );
  NAND2_X1 U810 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U811 ( .A(n764), .B(KEYINPUT126), .ZN(n769) );
  XNOR2_X1 U812 ( .A(G227), .B(n765), .ZN(n766) );
  NAND2_X1 U813 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U814 ( .A1(n767), .A2(G953), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n769), .A2(n768), .ZN(G72) );
  XOR2_X1 U816 ( .A(G137), .B(n770), .Z(G39) );
  XOR2_X1 U817 ( .A(n771), .B(G131), .Z(G33) );
endmodule

