//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT79), .B(G104), .ZN(new_n190));
  AOI21_X1  g004(.A(KEYINPUT80), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT79), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT79), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  AND4_X1   g009(.A1(KEYINPUT80), .A2(new_n193), .A3(new_n195), .A4(G107), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n192), .A2(KEYINPUT3), .A3(G107), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(G107), .B1(new_n193), .B2(new_n195), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G101), .B1(new_n197), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n194), .A2(G104), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n192), .A2(KEYINPUT79), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n198), .B1(new_n207), .B2(KEYINPUT3), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n193), .A2(new_n195), .A3(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n190), .A2(KEYINPUT80), .A3(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n203), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G119), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n220), .A3(G116), .ZN(new_n221));
  INV_X1    g035(.A(G116), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G119), .ZN(new_n223));
  INV_X1    g037(.A(G113), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n221), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n221), .B2(new_n223), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI211_X1 g046(.A(KEYINPUT67), .B(new_n228), .C1(new_n221), .C2(new_n223), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n214), .B1(new_n208), .B2(new_n213), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n216), .A2(new_n234), .A3(KEYINPUT85), .A4(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n204), .A2(G104), .ZN(new_n240));
  OAI21_X1  g054(.A(G101), .B1(new_n200), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n215), .A2(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n221), .A2(KEYINPUT5), .A3(new_n223), .ZN(new_n243));
  OAI21_X1  g057(.A(G113), .B1(new_n221), .B2(KEYINPUT5), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n229), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  AOI211_X1 g061(.A(new_n214), .B(new_n236), .C1(new_n208), .C2(new_n213), .ZN(new_n248));
  INV_X1    g062(.A(new_n231), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT67), .A3(new_n229), .ZN(new_n250));
  INV_X1    g064(.A(new_n233), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT85), .B1(new_n253), .B2(new_n216), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n189), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n216), .A2(new_n238), .A3(new_n234), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n258), .A2(new_n188), .A3(new_n246), .A4(new_n239), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(KEYINPUT6), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  INV_X1    g076(.A(G146), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT64), .B1(new_n263), .B2(G143), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n261), .A3(G146), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n263), .A2(G143), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(G146), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n267), .A2(new_n269), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G125), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n264), .A2(new_n266), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G128), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n272), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G128), .B1(new_n262), .B2(new_n279), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n274), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(G125), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G224), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G953), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n286), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n290), .B(new_n189), .C1(new_n247), .C2(new_n254), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n260), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n286), .B1(KEYINPUT86), .B2(new_n288), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n288), .ZN(new_n295));
  INV_X1    g109(.A(new_n288), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n286), .A2(KEYINPUT86), .A3(KEYINPUT7), .A4(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n242), .B(new_n245), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n188), .B(KEYINPUT8), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n295), .A2(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n300), .B2(new_n259), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n292), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n292), .B2(new_n301), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n187), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  INV_X1    g121(.A(G128), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n282), .B1(new_n267), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n215), .A2(new_n241), .A3(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n215), .A2(new_n241), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(new_n285), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT65), .ZN(new_n314));
  INV_X1    g128(.A(G137), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT11), .A2(G134), .ZN(new_n317));
  NAND2_X1  g131(.A1(KEYINPUT65), .A2(G137), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT11), .A2(G134), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT11), .A2(G134), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(G137), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G131), .ZN(new_n324));
  INV_X1    g138(.A(G131), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT12), .B1(new_n313), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n215), .A2(new_n241), .A3(new_n310), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n285), .B1(new_n215), .B2(new_n241), .ZN(new_n330));
  OAI211_X1 g144(.A(KEYINPUT12), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n276), .B1(new_n235), .B2(new_n237), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n334), .A2(new_n216), .B1(new_n335), .B2(new_n311), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n282), .B2(new_n284), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n215), .A2(new_n241), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT82), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n215), .A2(KEYINPUT82), .A3(new_n241), .A4(new_n337), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n327), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G110), .B(G140), .ZN(new_n345));
  INV_X1    g159(.A(G227), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n333), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n336), .A2(new_n342), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n327), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n349), .B1(new_n353), .B2(new_n344), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n306), .B(new_n307), .C1(new_n351), .C2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n306), .A2(new_n307), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n344), .B1(new_n328), .B2(new_n332), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n348), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n344), .A2(new_n360), .A3(new_n349), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n353), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n360), .B1(new_n344), .B2(new_n349), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n359), .B(G469), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G221), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(new_n368), .B2(new_n307), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT84), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n365), .A2(new_n373), .A3(new_n370), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n305), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT92), .ZN(new_n376));
  INV_X1    g190(.A(G237), .ZN(new_n377));
  INV_X1    g191(.A(G953), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G214), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(G143), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n380), .A2(new_n325), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n325), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT17), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G140), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT16), .B1(new_n385), .B2(G125), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT77), .A2(G125), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(G140), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(KEYINPUT16), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n389), .A2(new_n263), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n263), .ZN(new_n391));
  OR3_X1    g205(.A1(new_n380), .A2(new_n383), .A3(new_n325), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n384), .A2(new_n390), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n380), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(new_n325), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n380), .A2(new_n394), .A3(KEYINPUT18), .A4(G131), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n388), .A2(G146), .ZN(new_n400));
  XNOR2_X1  g214(.A(G125), .B(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n263), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT89), .B(G104), .Z(new_n405));
  XNOR2_X1  g219(.A(G113), .B(G122), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n393), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n393), .B2(new_n404), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n307), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT90), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT90), .B(new_n307), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(G475), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n416));
  NOR2_X1   g230(.A1(G475), .A2(G902), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n381), .A2(new_n382), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n401), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(KEYINPUT19), .B2(new_n388), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n263), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n422), .A3(new_n390), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n407), .B1(new_n404), .B2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n416), .B(new_n417), .C1(new_n409), .C2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n417), .ZN(new_n426));
  INV_X1    g240(.A(new_n424), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n408), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n429));
  OAI21_X1  g243(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n415), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n307), .B(new_n378), .C1(G234), .C2(G237), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(G898), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n378), .A2(G952), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(G234), .B2(G237), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n308), .A2(G143), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n261), .A2(G128), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G134), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G116), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(new_n204), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT13), .B1(new_n261), .B2(G128), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n441), .B1(KEYINPUT13), .B2(new_n440), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n444), .B(new_n446), .C1(new_n451), .C2(new_n443), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n442), .B(new_n443), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n222), .A2(KEYINPUT14), .A3(G122), .ZN(new_n454));
  INV_X1    g268(.A(new_n445), .ZN(new_n455));
  OAI211_X1 g269(.A(G107), .B(new_n454), .C1(new_n455), .C2(KEYINPUT14), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n453), .B(new_n456), .C1(G107), .C2(new_n455), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT74), .B(G217), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n367), .A2(new_n459), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n452), .A2(new_n457), .A3(new_n460), .ZN(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G478), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(KEYINPUT15), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n464), .B(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n432), .A2(new_n439), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n375), .A2(new_n376), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n187), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n292), .A2(new_n301), .ZN(new_n471));
  INV_X1    g285(.A(new_n302), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n292), .A2(new_n301), .A3(new_n302), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n374), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n373), .B1(new_n365), .B2(new_n370), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n475), .B(new_n468), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT92), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n459), .B1(G234), .B2(new_n307), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT24), .B(G110), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n308), .A2(G119), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT75), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT75), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n308), .A3(G119), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT76), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT66), .B(G119), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G128), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n488), .B1(new_n487), .B2(new_n490), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n482), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT23), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n483), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(G128), .B2(new_n489), .ZN(new_n496));
  INV_X1    g310(.A(G110), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n489), .B2(G128), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n496), .A2(KEYINPUT78), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT78), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n498), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(G110), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n390), .A2(new_n402), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n390), .A2(new_n391), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(G110), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n491), .A2(new_n492), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n482), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT22), .B(G137), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n378), .A2(G221), .A3(G234), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n511), .B(new_n512), .Z(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n505), .A2(new_n509), .A3(new_n513), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n307), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT25), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n515), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n516), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n481), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n516), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n513), .B1(new_n505), .B2(new_n509), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n480), .A2(G902), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n377), .A2(new_n378), .A3(G210), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT27), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(G101), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n267), .A2(new_n269), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n271), .A2(new_n274), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n319), .A2(new_n325), .A3(new_n322), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n325), .B1(new_n319), .B2(new_n322), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n316), .A2(new_n443), .A3(new_n318), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n325), .B1(G134), .B2(G137), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n280), .B(new_n262), .C1(new_n264), .C2(new_n266), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n272), .A2(new_n273), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(new_n309), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n326), .B(new_n539), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n536), .B(new_n543), .C1(new_n232), .C2(new_n233), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT68), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n326), .A2(new_n539), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n327), .A2(new_n275), .B1(new_n547), .B2(new_n285), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n548), .B2(new_n252), .ZN(new_n549));
  OAI211_X1 g363(.A(KEYINPUT69), .B(new_n531), .C1(new_n545), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n536), .A2(new_n543), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT30), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT30), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n536), .A2(new_n543), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n252), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n531), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n544), .A2(KEYINPUT68), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n252), .A2(new_n546), .A3(new_n543), .A4(new_n536), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(KEYINPUT69), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT31), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n551), .A2(KEYINPUT71), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n252), .B1(new_n551), .B2(KEYINPUT71), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n559), .A2(new_n560), .B1(new_n234), .B2(new_n551), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(new_n564), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n558), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n555), .B1(new_n561), .B2(KEYINPUT69), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n531), .B1(new_n545), .B2(new_n549), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT69), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT31), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT70), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT70), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n572), .A2(new_n575), .A3(new_n579), .A4(new_n576), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n571), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(G472), .A2(G902), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(KEYINPUT72), .Z(new_n583));
  OAI21_X1  g397(.A(KEYINPUT32), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(new_n580), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n572), .A2(new_n575), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n586), .A2(KEYINPUT31), .B1(new_n558), .B2(new_n569), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  INV_X1    g403(.A(new_n583), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n531), .B(new_n567), .C1(new_n568), .C2(new_n564), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT29), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n307), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n595), .A2(KEYINPUT73), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n556), .B1(new_n545), .B2(new_n549), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n558), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n594), .A3(new_n593), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(KEYINPUT73), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G472), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n527), .B1(new_n592), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n469), .A2(new_n479), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NOR2_X1   g419(.A1(new_n476), .A2(new_n477), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n588), .A2(new_n590), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n585), .B2(new_n587), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n606), .A2(new_n610), .A3(new_n527), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT93), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n187), .B(new_n439), .C1(new_n303), .C2(new_n304), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n462), .A2(new_n463), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT33), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n462), .A2(new_n616), .A3(new_n463), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(G478), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(G478), .A2(G902), .ZN(new_n619));
  INV_X1    g433(.A(new_n464), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n618), .B(new_n619), .C1(G478), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n431), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n612), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT96), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  OR2_X1    g444(.A1(new_n428), .A2(new_n429), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n428), .A2(new_n429), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n467), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n415), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n413), .A2(KEYINPUT97), .A3(G475), .A4(new_n414), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT98), .B1(new_n613), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n637), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n475), .A2(new_n639), .A3(new_n640), .A4(new_n439), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n612), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NAND2_X1  g459(.A1(new_n519), .A2(new_n520), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n480), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n514), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n510), .B(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n649), .A2(G902), .A3(new_n480), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n647), .A2(KEYINPUT99), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n521), .B2(new_n650), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n610), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n479), .A2(new_n469), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AOI21_X1  g473(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n660));
  AOI211_X1 g474(.A(KEYINPUT32), .B(new_n583), .C1(new_n585), .C2(new_n587), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n602), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n652), .A2(new_n654), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n433), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n438), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n637), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n375), .A2(new_n662), .A3(new_n663), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n666), .B(KEYINPUT39), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n671), .B(new_n672), .C1(new_n476), .C2(new_n477), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n663), .A2(new_n470), .A3(new_n432), .A4(new_n467), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT38), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n303), .B2(new_n304), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n473), .A2(KEYINPUT38), .A3(new_n474), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n568), .A2(new_n531), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n572), .B2(new_n575), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n681), .B2(G902), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n660), .B2(new_n661), .ZN(new_n683));
  AND4_X1   g497(.A1(new_n673), .A2(new_n674), .A3(new_n679), .A4(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n606), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n685), .A2(new_n672), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n684), .B1(new_n686), .B2(new_n671), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  NOR2_X1   g502(.A1(new_n623), .A2(new_n667), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n375), .A2(new_n662), .A3(new_n663), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  OAI21_X1  g505(.A(new_n307), .B1(new_n351), .B2(new_n354), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n370), .A3(new_n355), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n603), .A2(new_n624), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND3_X1  g512(.A1(new_n642), .A2(new_n603), .A3(new_n695), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  AOI21_X1  g514(.A(new_n655), .B1(new_n592), .B2(new_n602), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n305), .A2(new_n694), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n468), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  AOI21_X1  g518(.A(new_n467), .B1(new_n415), .B2(new_n430), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n475), .A2(new_n695), .A3(new_n439), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n609), .B2(new_n608), .ZN(new_n708));
  OAI211_X1 g522(.A(KEYINPUT100), .B(G472), .C1(new_n581), .C2(G902), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n607), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n706), .A2(new_n710), .A3(new_n526), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  NAND4_X1  g526(.A1(new_n710), .A2(new_n663), .A3(new_n689), .A4(new_n702), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  NAND2_X1  g528(.A1(new_n662), .A2(new_n526), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n473), .A2(new_n187), .A3(new_n474), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n362), .B2(new_n363), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n350), .A2(KEYINPUT83), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(KEYINPUT101), .A3(new_n353), .A4(new_n361), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(G469), .A3(new_n359), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n355), .A2(new_n357), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n369), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n473), .A2(KEYINPUT102), .A3(new_n187), .A4(new_n474), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n718), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n689), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n718), .A2(new_n728), .A3(new_n727), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n603), .A3(new_n689), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT103), .B(G131), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G33));
  NAND3_X1  g552(.A1(new_n732), .A2(new_n603), .A3(new_n668), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  XNOR2_X1  g554(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n431), .B2(new_n621), .ZN(new_n742));
  NOR2_X1   g556(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n622), .A2(new_n415), .A3(new_n430), .A4(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n742), .A2(new_n745), .B1(new_n652), .B2(new_n654), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n610), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n718), .A2(new_n728), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n746), .A2(new_n610), .A3(KEYINPUT44), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n718), .A2(new_n753), .A3(new_n728), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n749), .A2(new_n751), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n355), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  INV_X1    g571(.A(new_n359), .ZN(new_n758));
  AOI211_X1 g572(.A(new_n757), .B(new_n758), .C1(new_n720), .C2(new_n722), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n757), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(G469), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n357), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n756), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n723), .A2(KEYINPUT45), .A3(new_n359), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n306), .B1(new_n760), .B2(new_n757), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n356), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n369), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(KEYINPUT104), .A3(new_n672), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n355), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n763), .A2(new_n764), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n370), .B(new_n672), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n755), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n315), .ZN(G39));
  NAND2_X1  g592(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n370), .B1(new_n772), .B2(new_n773), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n750), .ZN(new_n784));
  INV_X1    g598(.A(new_n689), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n662), .A2(new_n526), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  OR2_X1    g602(.A1(G952), .A2(G953), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n306), .B(new_n758), .C1(new_n720), .C2(new_n722), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n370), .B1(new_n790), .B2(new_n725), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n705), .B(new_n187), .C1(new_n303), .C2(new_n304), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n666), .B(KEYINPUT109), .Z(new_n794));
  NAND3_X1  g608(.A1(new_n647), .A2(new_n651), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AND4_X1   g610(.A1(KEYINPUT110), .A2(new_n793), .A3(new_n683), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n795), .B1(new_n592), .B2(new_n682), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT110), .B1(new_n798), .B2(new_n793), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n701), .B(new_n375), .C1(new_n668), .C2(new_n689), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n713), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT52), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n793), .A2(new_n683), .A3(new_n796), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n798), .A2(KEYINPUT110), .A3(new_n793), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n713), .A4(new_n801), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n696), .A2(new_n699), .A3(new_n703), .A4(new_n711), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n736), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n708), .A2(new_n709), .A3(new_n607), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n814), .A2(new_n655), .A3(new_n785), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n730), .A2(new_n668), .B1(new_n815), .B2(new_n732), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT107), .ZN(new_n817));
  INV_X1    g631(.A(new_n467), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n432), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n613), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n817), .B1(new_n613), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n623), .B2(new_n613), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n611), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n479), .B(new_n469), .C1(new_n603), .C2(new_n656), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n467), .A2(new_n666), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n631), .B2(new_n632), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n826), .A2(new_n635), .A3(new_n636), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n718), .A2(new_n728), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT108), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT108), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n718), .A2(new_n827), .A3(new_n830), .A4(new_n728), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n829), .A2(new_n685), .A3(new_n701), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n816), .A2(new_n823), .A3(new_n824), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n813), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n811), .A2(new_n834), .A3(KEYINPUT53), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n824), .A2(new_n823), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n815), .A2(new_n732), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n832), .A2(new_n739), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n839), .A3(new_n736), .A4(new_n812), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n803), .A2(new_n810), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n835), .A2(new_n842), .A3(KEYINPUT111), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n844), .B(new_n836), .C1(new_n840), .C2(new_n841), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(KEYINPUT54), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n833), .A2(new_n836), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n812), .A2(new_n736), .A3(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n731), .A2(new_n735), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n699), .A2(new_n696), .A3(new_n703), .A4(new_n711), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT112), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n811), .A2(new_n847), .A3(new_n849), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n842), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT113), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n853), .A2(new_n857), .A3(new_n842), .A4(new_n854), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n846), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n784), .A2(new_n695), .ZN(new_n860));
  INV_X1    g674(.A(new_n683), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n437), .A3(new_n526), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n860), .A2(new_n862), .A3(new_n431), .A4(new_n622), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n678), .A2(new_n470), .A3(new_n695), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT114), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT50), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n438), .B1(new_n742), .B2(new_n745), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n710), .A2(new_n526), .A3(new_n867), .ZN(new_n868));
  OR3_X1    g682(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n865), .B2(new_n868), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n784), .A2(new_n695), .A3(new_n867), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT115), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(KEYINPUT115), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n663), .A3(new_n710), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n871), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n693), .A2(new_n355), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n779), .B(new_n782), .C1(new_n370), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n751), .A2(new_n754), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n868), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n878), .A2(KEYINPUT51), .A3(new_n880), .A4(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n860), .A2(new_n862), .A3(new_n623), .ZN(new_n887));
  INV_X1    g701(.A(new_n868), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n436), .B(new_n887), .C1(new_n702), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT48), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n875), .B2(new_n603), .ZN(new_n891));
  AOI211_X1 g705(.A(KEYINPUT48), .B(new_n715), .C1(new_n873), .C2(new_n874), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n871), .A2(new_n885), .A3(new_n876), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n789), .B1(new_n859), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n881), .A2(KEYINPUT49), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n526), .A2(new_n370), .A3(new_n187), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n881), .A2(KEYINPUT49), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n432), .A2(new_n622), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n678), .A3(new_n861), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n898), .A2(new_n904), .ZN(G75));
  NAND2_X1  g719(.A1(new_n260), .A2(new_n291), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n289), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT55), .Z(new_n908));
  INV_X1    g722(.A(G210), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n909), .B(new_n307), .C1(new_n853), .C2(new_n842), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(KEYINPUT56), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n378), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n910), .A2(KEYINPUT56), .A3(new_n908), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(G51));
  AOI21_X1  g730(.A(new_n307), .B1(new_n853), .B2(new_n842), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n759), .A2(new_n762), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n917), .A2(KEYINPUT117), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT117), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n356), .B(KEYINPUT57), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n853), .A2(new_n854), .A3(new_n842), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n854), .B1(new_n853), .B2(new_n842), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n351), .A2(new_n354), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n912), .B1(new_n921), .B2(new_n927), .ZN(G54));
  NAND2_X1  g742(.A1(new_n427), .A2(new_n408), .ZN(new_n929));
  AND2_X1   g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n917), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n917), .B2(new_n930), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n912), .ZN(G60));
  AND2_X1   g747(.A1(new_n615), .A2(new_n617), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n619), .B(KEYINPUT59), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n923), .B2(new_n924), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n913), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n859), .A2(new_n936), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n934), .ZN(G63));
  XNOR2_X1  g755(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n853), .A2(new_n842), .ZN(new_n944));
  INV_X1    g758(.A(new_n649), .ZN(new_n945));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT118), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT60), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n913), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n524), .B(KEYINPUT119), .Z(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n944), .B2(new_n948), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n943), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n953), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(new_n913), .A3(new_n949), .A4(new_n942), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(G66));
  OAI21_X1  g771(.A(G953), .B1(new_n434), .B2(new_n287), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n837), .A2(new_n812), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n960), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n906), .B1(G898), .B2(new_n378), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  OAI21_X1  g777(.A(G953), .B1(new_n346), .B2(new_n664), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT124), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n552), .A2(new_n554), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT121), .Z(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(new_n421), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(G900), .B2(G953), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n715), .A2(new_n792), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT104), .B1(new_n770), .B2(new_n672), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n774), .A2(new_n775), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g789(.A1(new_n731), .A2(new_n735), .B1(new_n668), .B2(new_n730), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n787), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT122), .ZN(new_n978));
  AND4_X1   g792(.A1(new_n978), .A2(new_n713), .A3(new_n669), .A4(new_n690), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n801), .B2(new_n713), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT125), .B1(new_n981), .B2(new_n777), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n802), .A2(KEYINPUT122), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n801), .A2(new_n978), .A3(new_n713), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n755), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n973), .B2(new_n974), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n977), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n971), .B1(new_n990), .B2(new_n378), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n992));
  INV_X1    g806(.A(new_n787), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n687), .B1(new_n979), .B2(new_n980), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n687), .B(KEYINPUT62), .C1(new_n979), .C2(new_n980), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT123), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n819), .A2(new_n623), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n686), .A2(new_n603), .A3(new_n784), .A4(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n987), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1001), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT123), .B1(new_n777), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(G953), .B1(new_n998), .B2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g820(.A1(new_n991), .A2(new_n992), .B1(new_n1006), .B2(new_n968), .ZN(new_n1007));
  AOI211_X1 g821(.A(KEYINPUT127), .B(new_n971), .C1(new_n990), .C2(new_n378), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n965), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n996), .A2(new_n997), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n1005), .A3(new_n787), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n378), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n965), .B1(new_n1013), .B2(new_n969), .ZN(new_n1014));
  INV_X1    g828(.A(new_n991), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n968), .B1(new_n1012), .B2(new_n378), .ZN(new_n1017));
  NOR4_X1   g831(.A1(new_n1017), .A2(new_n991), .A3(KEYINPUT126), .A4(new_n965), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1009), .B1(new_n1016), .B2(new_n1018), .ZN(G72));
  NAND2_X1  g833(.A1(new_n990), .A2(new_n960), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  AOI211_X1 g836(.A(new_n531), .B(new_n597), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n598), .A2(new_n586), .ZN(new_n1024));
  AND4_X1   g838(.A1(new_n845), .A2(new_n843), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n597), .A2(new_n531), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n998), .A2(new_n960), .A3(new_n1005), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1026), .B1(new_n1027), .B2(new_n1022), .ZN(new_n1028));
  NOR4_X1   g842(.A1(new_n1023), .A2(new_n1025), .A3(new_n912), .A4(new_n1028), .ZN(G57));
endmodule


