//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G58), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  OR3_X1    g0017(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n218));
  OAI21_X1  g0018(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT65), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n225), .A2(G1), .A3(G13), .ZN(new_n226));
  AND2_X1   g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n201), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n217), .B(new_n222), .C1(new_n229), .C2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n245), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(KEYINPUT67), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n227), .A2(KEYINPUT68), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(KEYINPUT68), .B1(new_n227), .B2(new_n257), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G50), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT69), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(new_n208), .A3(KEYINPUT8), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n228), .A2(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n260), .A2(new_n275), .B1(new_n202), .B2(new_n263), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n266), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT9), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  AND2_X1   g0079(.A1(G1), .A2(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(new_n280), .B2(new_n281), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(G226), .B2(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n224), .A2(new_n226), .B1(G33), .B2(G41), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G222), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G223), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(G77), .B2(new_n292), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n289), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(G200), .B2(new_n298), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n278), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT10), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n298), .A2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(new_n298), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n277), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n267), .A2(G50), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n247), .A2(G20), .ZN(new_n309));
  INV_X1    g0109(.A(G77), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n308), .B(new_n309), .C1(new_n310), .C2(new_n274), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n260), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n313));
  XOR2_X1   g0113(.A(new_n312), .B(new_n313), .Z(new_n314));
  XNOR2_X1  g0114(.A(new_n262), .B(KEYINPUT70), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n260), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(G68), .A3(new_n265), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT12), .B1(new_n315), .B2(G68), .ZN(new_n319));
  INV_X1    g0119(.A(G13), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G1), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT12), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n319), .B1(new_n309), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n314), .B1(KEYINPUT75), .B2(new_n325), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n325), .A2(KEYINPUT75), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n288), .A2(G238), .B1(new_n285), .B2(new_n282), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G33), .A3(G97), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n294), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n209), .A2(G1698), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n337), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT73), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n335), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n290), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n335), .B2(new_n343), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n330), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n330), .C1(new_n346), .C2(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n299), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(G200), .B2(new_n352), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n329), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n317), .A2(G77), .A3(new_n265), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT71), .ZN(new_n357));
  INV_X1    g0157(.A(new_n269), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT15), .B(G87), .Z(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n274), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n260), .A2(new_n362), .B1(new_n310), .B2(new_n316), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n288), .A2(G244), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n292), .A2(G232), .A3(new_n294), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n292), .A2(G238), .A3(G1698), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n292), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n287), .B(new_n365), .C1(new_n369), .C2(new_n290), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G169), .B2(new_n370), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n364), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n357), .A2(new_n363), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n370), .A2(G190), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n370), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n303), .A2(new_n307), .A3(new_n355), .A4(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n273), .B1(new_n261), .B2(G20), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT68), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n255), .A2(new_n256), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n224), .A2(new_n226), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n227), .A2(KEYINPUT68), .A3(new_n257), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n382), .A2(new_n388), .A3(new_n262), .ZN(new_n389));
  INV_X1    g0189(.A(new_n273), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n262), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n208), .A2(new_n247), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n392), .A2(new_n201), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(G20), .B1(G159), .B2(new_n267), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n228), .A2(KEYINPUT7), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n337), .B2(new_n341), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n340), .A2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n228), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT78), .B1(new_n402), .B2(new_n247), .ZN(new_n403));
  AOI21_X1  g0203(.A(G20), .B1(new_n337), .B2(new_n341), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n404), .A2(KEYINPUT7), .B1(new_n396), .B2(new_n292), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT78), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(G68), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n395), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n388), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT79), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n340), .B2(G33), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n336), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n341), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT80), .ZN(new_n414));
  INV_X1    g0214(.A(new_n396), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n401), .B1(new_n292), .B2(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n419));
  OAI21_X1  g0219(.A(G68), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT16), .B1(new_n420), .B2(new_n394), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n391), .B1(new_n409), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n287), .B1(G232), .B2(new_n288), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n338), .A2(G1698), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G223), .B2(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n337), .A2(new_n341), .ZN(new_n427));
  INV_X1    g0227(.A(G87), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n426), .A2(new_n427), .B1(new_n336), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n290), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n424), .A2(G179), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n305), .B1(new_n424), .B2(new_n430), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT18), .B1(new_n423), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n264), .A2(new_n382), .B1(new_n263), .B2(new_n273), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n427), .A2(new_n415), .ZN(new_n436));
  AOI211_X1 g0236(.A(KEYINPUT78), .B(new_n247), .C1(new_n417), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n406), .B1(new_n405), .B2(G68), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT16), .B(new_n394), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n260), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n435), .B1(new_n440), .B2(new_n421), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  INV_X1    g0242(.A(new_n433), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n424), .A2(new_n299), .A3(new_n430), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n288), .A2(G232), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n430), .A2(new_n286), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(G200), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n435), .B(new_n448), .C1(new_n440), .C2(new_n421), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n419), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n417), .A3(new_n416), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n395), .B1(new_n453), .B2(G68), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n439), .B(new_n260), .C1(new_n454), .C2(KEYINPUT16), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n435), .A4(new_n448), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n434), .A2(new_n444), .A3(new_n451), .A4(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n349), .A2(G179), .A3(new_n351), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT76), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT76), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n349), .A2(new_n460), .A3(G179), .A4(new_n351), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n352), .A2(G169), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT14), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT14), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n352), .A2(new_n465), .A3(G169), .ZN(new_n466));
  AND4_X1   g0266(.A1(KEYINPUT77), .A2(new_n462), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n352), .B2(G169), .ZN(new_n468));
  AOI211_X1 g0268(.A(KEYINPUT14), .B(new_n305), .C1(new_n349), .C2(new_n351), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT77), .B1(new_n470), .B2(new_n462), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n328), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n381), .A2(new_n457), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n337), .A2(new_n341), .A3(G244), .A4(new_n294), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n294), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n290), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n280), .A2(new_n281), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n261), .B(G45), .C1(new_n283), .C2(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT5), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G41), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT82), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n485), .B2(G41), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n283), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n284), .A2(G1), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(G41), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n483), .A2(G274), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n487), .A2(new_n211), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n482), .A2(new_n299), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n481), .B2(new_n290), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(G200), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n262), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n261), .A2(G33), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT81), .ZN(new_n502));
  AOI211_X1 g0302(.A(new_n263), .B(new_n502), .C1(new_n386), .C2(new_n387), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n503), .B2(G97), .ZN(new_n504));
  OAI21_X1  g0304(.A(G107), .B1(new_n418), .B2(new_n419), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n368), .A2(KEYINPUT6), .A3(G97), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n210), .A2(new_n368), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n260), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n499), .A2(new_n504), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n211), .A2(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G250), .B2(G1698), .ZN(new_n516));
  INV_X1    g0316(.A(G294), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n516), .A2(new_n427), .B1(new_n336), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n290), .ZN(new_n519));
  INV_X1    g0319(.A(new_n484), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n520), .A2(new_n282), .A3(new_n489), .A4(new_n490), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n483), .B(G264), .C1(new_n484), .C2(new_n486), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n519), .A2(G190), .A3(new_n521), .A4(new_n522), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n337), .A2(new_n341), .A3(new_n228), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n292), .A2(new_n529), .A3(new_n228), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g0331(.A(KEYINPUT86), .B(KEYINPUT24), .Z(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G116), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G20), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n228), .B2(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n368), .A2(KEYINPUT23), .A3(G20), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n532), .B1(new_n531), .B2(new_n538), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n260), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n503), .A2(G107), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n262), .A2(G107), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n544), .B(KEYINPUT25), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n526), .A2(new_n542), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT83), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n482), .A2(new_n496), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(G179), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n498), .A2(KEYINPUT83), .A3(new_n371), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n388), .B1(new_n505), .B2(new_n511), .ZN(new_n552));
  INV_X1    g0352(.A(new_n500), .ZN(new_n553));
  INV_X1    g0353(.A(new_n502), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n262), .B(new_n554), .C1(new_n258), .C2(new_n259), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(new_n210), .ZN(new_n556));
  OAI22_X1  g0356(.A1(new_n552), .A2(new_n556), .B1(G169), .B2(new_n498), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n514), .B(new_n546), .C1(new_n551), .C2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G257), .A2(G1698), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n294), .A2(G264), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n292), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G303), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n427), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n290), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n483), .B(G270), .C1(new_n484), .C2(new_n486), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n521), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G169), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n315), .A2(G116), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT20), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n385), .B1(new_n255), .B2(new_n256), .ZN(new_n571));
  AOI21_X1  g0371(.A(G20), .B1(G33), .B2(G283), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n336), .A2(G97), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n572), .A2(new_n573), .B1(G20), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n570), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT20), .B(new_n575), .C1(new_n384), .C2(new_n385), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n502), .A2(new_n574), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n388), .A2(new_n315), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n568), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT85), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(KEYINPUT21), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n579), .A2(new_n581), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n567), .A2(new_n371), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n582), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n568), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n584), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n567), .A2(new_n299), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n567), .A2(G200), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n592), .A2(new_n579), .A3(new_n581), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n588), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n523), .A2(G169), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT87), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n519), .A2(G179), .A3(new_n521), .A4(new_n522), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n598), .A2(new_n597), .ZN(new_n600));
  INV_X1    g0400(.A(new_n541), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n388), .B1(new_n601), .B2(new_n539), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n545), .B1(new_n555), .B2(new_n368), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n599), .B(new_n600), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n491), .A2(new_n279), .ZN(new_n605));
  INV_X1    g0405(.A(G250), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n284), .B2(G1), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n483), .A3(new_n607), .ZN(new_n608));
  MUX2_X1   g0408(.A(G238), .B(G244), .S(G1698), .Z(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(new_n292), .B1(G33), .B2(G116), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n610), .B2(new_n291), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(new_n299), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n315), .A2(new_n360), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n508), .A2(new_n428), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT19), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n332), .B2(new_n334), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n617), .B2(G20), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n274), .B2(new_n210), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(KEYINPUT84), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n292), .A2(new_n228), .A3(G68), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(KEYINPUT84), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n618), .A2(new_n620), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n614), .B1(new_n260), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n611), .A2(G200), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n388), .A2(G87), .A3(new_n262), .A4(new_n554), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n613), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n624), .B1(new_n361), .B2(new_n555), .ZN(new_n628));
  INV_X1    g0428(.A(new_n608), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n609), .A2(new_n292), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n533), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n629), .B1(new_n631), .B2(new_n290), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n371), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n611), .A2(new_n305), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n604), .A2(new_n627), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n595), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n474), .A2(new_n559), .A3(new_n639), .ZN(G372));
  AND2_X1   g0440(.A1(new_n451), .A2(new_n456), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n375), .B(new_n372), .C1(G169), .C2(new_n370), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n329), .B2(new_n354), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n473), .B2(new_n643), .ZN(new_n644));
  AOI211_X1 g0444(.A(KEYINPUT18), .B(new_n433), .C1(new_n455), .C2(new_n435), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n442), .B1(new_n441), .B2(new_n443), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n303), .B1(new_n277), .B2(new_n306), .ZN(new_n649));
  INV_X1    g0449(.A(new_n474), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n503), .A2(new_n360), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n635), .B1(new_n651), .B2(new_n624), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT88), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n612), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n624), .A2(new_n626), .A3(KEYINPUT88), .A4(new_n625), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n551), .A2(new_n557), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n504), .A2(new_n513), .B1(new_n305), .B2(new_n548), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n549), .A2(new_n550), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n637), .A2(new_n627), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT26), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n660), .A2(new_n637), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n588), .A2(new_n591), .A3(new_n604), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n558), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT89), .B1(new_n669), .B2(new_n657), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n552), .A2(new_n556), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n661), .A2(new_n662), .B1(new_n671), .B2(new_n499), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n588), .A2(new_n591), .A3(new_n604), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(new_n657), .A3(new_n546), .A4(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n667), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n649), .B1(new_n650), .B2(new_n678), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n321), .A2(new_n228), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(G213), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n586), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n588), .B2(new_n591), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n588), .A2(new_n591), .A3(new_n594), .A4(new_n686), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT91), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT91), .B1(new_n690), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n604), .A2(new_n685), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n685), .B1(new_n602), .B2(new_n603), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n546), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n695), .B1(new_n697), .B2(new_n604), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n694), .A2(G330), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n685), .B1(new_n588), .B2(new_n591), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n695), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n220), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n508), .A2(new_n428), .A3(new_n574), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n261), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n232), .B2(new_n705), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  INV_X1    g0509(.A(new_n685), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n677), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT96), .ZN(new_n714));
  INV_X1    g0514(.A(new_n657), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT26), .B1(new_n715), .B2(new_n663), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n659), .A2(new_n658), .A3(new_n627), .A4(new_n637), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n652), .B(KEYINPUT97), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(new_n674), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .A3(new_n710), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT96), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n711), .A2(new_n721), .A3(new_n712), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n714), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n587), .A2(new_n498), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT92), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n632), .A2(new_n725), .A3(new_n522), .A4(new_n519), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n519), .A2(new_n522), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT92), .B1(new_n727), .B2(new_n611), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n724), .A2(new_n729), .A3(KEYINPUT30), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n632), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n548), .A3(new_n523), .A4(new_n567), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT93), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n587), .A2(new_n498), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n726), .B2(new_n728), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT30), .B1(new_n724), .B2(new_n729), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT93), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n733), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n740), .A2(new_n685), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT94), .B1(new_n741), .B2(KEYINPUT31), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT31), .B1(new_n740), .B2(new_n685), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT94), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n733), .B1(KEYINPUT30), .B2(new_n736), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n742), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n639), .A2(new_n559), .A3(new_n710), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT95), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT95), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n639), .A2(new_n559), .A3(new_n751), .A4(new_n710), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(G330), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n723), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n709), .B1(new_n756), .B2(G1), .ZN(G364));
  NAND2_X1  g0557(.A1(new_n694), .A2(G330), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT98), .Z(new_n759));
  NOR2_X1   g0559(.A1(new_n320), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n261), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n759), .B1(G330), .B2(new_n694), .C1(new_n705), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n705), .A2(new_n762), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT99), .Z(new_n765));
  NOR2_X1   g0565(.A1(new_n704), .A2(new_n292), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n232), .A2(new_n284), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n766), .B(new_n767), .C1(new_n284), .C2(new_n251), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n220), .A2(G355), .A3(new_n292), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n768), .B(new_n769), .C1(G116), .C2(new_n220), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(KEYINPUT100), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n227), .B1(G20), .B2(new_n305), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n770), .B2(KEYINPUT100), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n765), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n228), .A2(G179), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G190), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n228), .A2(new_n371), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n780), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n377), .A2(G190), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n779), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n310), .B1(new_n789), .B2(new_n368), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G87), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n299), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n228), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n210), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n786), .A2(G190), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G200), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(G58), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n786), .A2(new_n788), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n292), .B1(new_n800), .B2(new_n247), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n797), .A2(new_n377), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G50), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n785), .A2(new_n793), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n802), .ZN(new_n805));
  INV_X1    g0605(.A(G326), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n805), .A2(new_n806), .B1(new_n517), .B2(new_n795), .ZN(new_n807));
  INV_X1    g0607(.A(new_n787), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n807), .A2(KEYINPUT102), .B1(G311), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(KEYINPUT102), .B2(new_n807), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT103), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n427), .B1(new_n791), .B2(new_n563), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT104), .Z(new_n813));
  NAND2_X1  g0613(.A1(new_n798), .A2(G322), .ZN(new_n814));
  INV_X1    g0614(.A(new_n781), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(new_n800), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT33), .B(G317), .ZN(new_n818));
  INV_X1    g0618(.A(new_n789), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n817), .A2(new_n818), .B1(new_n819), .B2(G283), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n804), .B1(new_n811), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n778), .B1(new_n822), .B2(new_n772), .ZN(new_n823));
  INV_X1    g0623(.A(new_n775), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n694), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n763), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n368), .A2(new_n791), .B1(new_n800), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n292), .B(new_n829), .C1(G116), .C2(new_n808), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n789), .A2(new_n428), .B1(new_n781), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT105), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n798), .A2(G294), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n796), .B1(G303), .B2(new_n802), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n830), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G150), .A2(new_n817), .B1(new_n808), .B2(G159), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n798), .A2(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n805), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n791), .A2(new_n202), .B1(new_n781), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n789), .A2(new_n247), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n844), .A2(new_n427), .A3(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n842), .B(new_n846), .C1(new_n208), .C2(new_n795), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n840), .A2(new_n841), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n836), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n772), .ZN(new_n850));
  INV_X1    g0650(.A(new_n765), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n772), .A2(new_n773), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(new_n310), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n364), .A2(new_n710), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n642), .B1(new_n854), .B2(new_n379), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n374), .A2(new_n710), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n850), .B(new_n853), .C1(new_n858), .C2(new_n774), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n374), .A2(new_n379), .A3(new_n685), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n677), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n858), .B1(new_n677), .B2(new_n710), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n863), .A2(KEYINPUT106), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(KEYINPUT106), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n754), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n866), .A2(new_n867), .B1(new_n705), .B2(new_n762), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n859), .B1(new_n868), .B2(new_n869), .ZN(G384));
  OR2_X1    g0670(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n871), .A2(G116), .A3(new_n229), .A4(new_n872), .ZN(new_n873));
  XOR2_X1   g0673(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n874));
  XNOR2_X1  g0674(.A(new_n873), .B(new_n874), .ZN(new_n875));
  OR3_X1    g0675(.A1(new_n231), .A2(new_n310), .A3(new_n392), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n261), .B(G13), .C1(new_n876), .C2(new_n246), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT108), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n472), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT77), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n464), .A2(new_n466), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n459), .A2(new_n461), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n470), .A2(KEYINPUT77), .A3(new_n462), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(KEYINPUT108), .A3(new_n328), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n685), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT109), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n394), .B1(new_n437), .B2(new_n438), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT16), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n391), .B1(new_n409), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n449), .B1(new_n894), .B2(new_n683), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n433), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n441), .A2(new_n443), .ZN(new_n898));
  INV_X1    g0698(.A(new_n683), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n441), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n898), .A2(new_n900), .A3(new_n901), .A4(new_n449), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n894), .A2(new_n683), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n457), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n903), .A2(new_n905), .A3(KEYINPUT38), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n890), .B(KEYINPUT39), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n898), .A2(new_n900), .A3(new_n449), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n902), .ZN(new_n911));
  INV_X1    g0711(.A(new_n900), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n457), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n903), .A2(new_n905), .A3(KEYINPUT38), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n908), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n403), .A2(new_n407), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT16), .B1(new_n921), .B2(new_n394), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n435), .B1(new_n440), .B2(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n423), .A2(new_n448), .B1(new_n923), .B2(new_n899), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n443), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n901), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND4_X1   g0726(.A1(new_n901), .A2(new_n898), .A3(new_n900), .A4(new_n449), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n904), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n647), .B2(new_n641), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n915), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n918), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n890), .B1(new_n932), .B2(KEYINPUT39), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n889), .B1(new_n920), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n647), .A2(new_n899), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n710), .B1(new_n326), .B2(new_n327), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n329), .B2(new_n354), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n880), .A2(new_n887), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n886), .A2(new_n936), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n861), .A2(new_n856), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n935), .B1(new_n940), .B2(new_n932), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n934), .A2(KEYINPUT110), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT110), .B1(new_n934), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n714), .A2(new_n474), .A3(new_n720), .A4(new_n722), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n649), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n938), .A2(new_n939), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n750), .A2(new_n752), .ZN(new_n949));
  INV_X1    g0749(.A(new_n739), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n730), .B(new_n732), .C1(new_n738), .C2(KEYINPUT93), .ZN(new_n951));
  OAI211_X1 g0751(.A(KEYINPUT31), .B(new_n685), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n743), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n948), .A2(new_n858), .A3(new_n932), .A4(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(new_n916), .B2(new_n918), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n959), .A2(new_n948), .A3(new_n858), .A4(new_n955), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n474), .A2(new_n955), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(G330), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n947), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n261), .B2(new_n760), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n947), .A2(new_n965), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n878), .B1(new_n967), .B2(new_n968), .ZN(G367));
  OAI21_X1  g0769(.A(new_n685), .B1(new_n552), .B2(new_n556), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n672), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(new_n604), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n685), .B1(new_n972), .B2(new_n663), .ZN(new_n973));
  INV_X1    g0773(.A(new_n971), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n659), .B2(new_n685), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n701), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n973), .B1(new_n977), .B2(KEYINPUT42), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(KEYINPUT42), .B2(new_n977), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT43), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n710), .B1(new_n624), .B2(new_n626), .ZN(new_n981));
  MUX2_X1   g0781(.A(new_n715), .B(new_n637), .S(new_n981), .Z(new_n982));
  OAI21_X1  g0782(.A(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n980), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n699), .A2(new_n975), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n985), .B(new_n986), .Z(new_n987));
  INV_X1    g0787(.A(KEYINPUT112), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n975), .A2(new_n701), .A3(new_n695), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n976), .A2(KEYINPUT45), .A3(new_n702), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n976), .B2(new_n702), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n975), .B(KEYINPUT44), .C1(new_n695), .C2(new_n701), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n990), .A2(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT111), .B1(new_n995), .B2(new_n699), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n699), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n995), .A2(KEYINPUT111), .A3(new_n699), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n698), .B(new_n700), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n758), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n759), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n756), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n988), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n998), .A2(new_n999), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1006), .A2(KEYINPUT112), .A3(new_n756), .A4(new_n1003), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n755), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n705), .B(KEYINPUT41), .Z(new_n1009));
  OAI21_X1  g0809(.A(KEYINPUT113), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n761), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1008), .A2(KEYINPUT113), .A3(new_n1009), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n987), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n766), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n237), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n776), .B1(new_n220), .B2(new_n361), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n765), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n795), .A2(new_n247), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n427), .B(new_n1018), .C1(G159), .C2(new_n817), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G50), .A2(new_n808), .B1(new_n815), .B2(G137), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n792), .A2(G58), .B1(new_n819), .B2(G77), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G143), .A2(new_n802), .B1(new_n798), .B2(G150), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n792), .A2(G116), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT46), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n368), .B2(new_n795), .C1(new_n831), .C2(new_n805), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n427), .B1(new_n789), .B2(new_n210), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G303), .B2(new_n798), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G283), .A2(new_n808), .B1(new_n817), .B2(G294), .ZN(new_n1029));
  INV_X1    g0829(.A(G317), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1028), .B(new_n1029), .C1(new_n1030), .C2(new_n781), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1023), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1017), .B1(new_n1033), .B2(new_n772), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT114), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n982), .A2(new_n775), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1013), .A2(new_n1038), .ZN(G387));
  INV_X1    g0839(.A(new_n705), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1003), .B2(new_n756), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT116), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT116), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n756), .C2(new_n1003), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n241), .A2(new_n284), .A3(new_n292), .ZN(new_n1045));
  OR3_X1    g0845(.A1(new_n269), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT50), .B1(new_n269), .B2(G50), .ZN(new_n1047));
  AOI21_X1  g0847(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n706), .B1(new_n1049), .B2(new_n427), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n220), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n776), .C1(new_n368), .C2(new_n220), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n765), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n698), .A2(new_n824), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n310), .A2(new_n791), .B1(new_n787), .B2(new_n247), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G150), .B2(new_n815), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n292), .B1(new_n789), .B2(new_n210), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G50), .B2(new_n798), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n390), .A2(new_n817), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n795), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n360), .A2(new_n1060), .B1(new_n802), .B2(G159), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n292), .B1(new_n819), .B2(G116), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n795), .A2(new_n828), .B1(new_n791), .B2(new_n517), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G303), .A2(new_n808), .B1(new_n817), .B2(G311), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT115), .B(G322), .Z(new_n1066));
  INV_X1    g0866(.A(new_n798), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1065), .B1(new_n805), .B2(new_n1066), .C1(new_n1030), .C2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1063), .B1(new_n806), .B2(new_n781), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1062), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1053), .B(new_n1054), .C1(new_n772), .C2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1003), .B2(new_n762), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1044), .A2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n995), .B(new_n699), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1040), .B1(new_n1004), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1080), .A2(new_n761), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n975), .A2(new_n775), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1014), .A2(new_n245), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n776), .B1(new_n210), .B2(new_n220), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n765), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G294), .A2(new_n808), .B1(new_n817), .B2(G303), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n574), .B2(new_n795), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT117), .Z(new_n1090));
  AOI22_X1  g0890(.A1(G311), .A2(new_n798), .B1(new_n802), .B2(G317), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT52), .Z(new_n1092));
  OAI22_X1  g0892(.A1(new_n1066), .A2(new_n781), .B1(new_n791), .B2(new_n828), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n292), .B(new_n1093), .C1(G107), .C2(new_n819), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G150), .A2(new_n802), .B1(new_n798), .B2(G159), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n795), .A2(new_n310), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n427), .B(new_n1098), .C1(G87), .C2(new_n819), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n358), .A2(new_n808), .B1(new_n817), .B2(G50), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n792), .A2(G68), .B1(new_n815), .B2(G143), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1095), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT118), .Z(new_n1104));
  AOI21_X1  g0904(.A(new_n1087), .B1(new_n1104), .B2(new_n772), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1083), .B1(new_n1084), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1082), .A2(new_n1106), .ZN(G390));
  OAI211_X1 g0907(.A(G330), .B(new_n858), .C1(new_n748), .C2(new_n753), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n948), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n719), .A2(new_n855), .A3(new_n710), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(new_n856), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n948), .ZN(new_n1113));
  INV_X1    g0913(.A(G330), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n949), .B2(new_n954), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n858), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1110), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1113), .A2(new_n857), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1119), .A2(new_n1115), .B1(new_n1113), .B2(new_n1108), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n861), .A2(new_n856), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1118), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n474), .A2(new_n1115), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n945), .A2(new_n649), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n945), .A2(new_n649), .A3(KEYINPUT119), .A4(new_n1124), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1123), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n889), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT38), .B1(new_n911), .B2(new_n913), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1130), .B1(new_n906), .B2(new_n1131), .C1(new_n1113), .C2(new_n1112), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n917), .B1(new_n931), .B2(new_n918), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n906), .A2(new_n1131), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1133), .A2(new_n890), .B1(new_n1134), .B2(new_n917), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n932), .A2(KEYINPUT39), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT109), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n889), .C2(new_n940), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1132), .A2(new_n1138), .A3(new_n1110), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1119), .A2(new_n1115), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1040), .B1(new_n1129), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1142), .B2(new_n1129), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1141), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1140), .B2(new_n1110), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n762), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n852), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n765), .B1(new_n390), .B2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n787), .A2(new_n210), .B1(new_n781), .B2(new_n517), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n845), .B(new_n1150), .C1(G107), .C2(new_n817), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n292), .B(new_n1098), .C1(G87), .C2(new_n792), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G116), .A2(new_n798), .B1(new_n802), .B2(G283), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n792), .A2(G150), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n815), .A2(G125), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1157), .B1(new_n839), .B2(new_n800), .C1(new_n787), .C2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G159), .A2(new_n1060), .B1(new_n802), .B2(G128), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n843), .C2(new_n1067), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n292), .B1(new_n789), .B2(new_n202), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT120), .Z(new_n1164));
  OAI21_X1  g0964(.A(new_n1154), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1149), .B1(new_n1165), .B2(new_n772), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n920), .A2(new_n933), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n1168), .B2(new_n774), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1144), .A2(new_n1147), .A3(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(KEYINPUT110), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1130), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1121), .A2(new_n932), .A3(new_n948), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n935), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1171), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n934), .A2(new_n941), .A3(KEYINPUT110), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n307), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n277), .A3(new_n899), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n277), .A2(new_n899), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n303), .A2(new_n307), .A3(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n956), .A2(new_n957), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n960), .A2(G330), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI221_X4 g0992(.A(new_n857), .B1(new_n949), .B2(new_n954), .C1(new_n938), .C2(new_n939), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1114), .B1(new_n1193), .B2(new_n959), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n958), .A3(new_n1188), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(KEYINPUT122), .B1(new_n1178), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT123), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1178), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1178), .B2(new_n1196), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT122), .ZN(new_n1202));
  AND4_X1   g1002(.A1(G330), .A2(new_n958), .A3(new_n1188), .A4(new_n960), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1188), .B1(new_n1194), .B2(new_n958), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1202), .B1(new_n1205), .B2(new_n944), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1203), .A2(new_n1204), .B1(new_n942), .B2(new_n943), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT123), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1178), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1201), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1123), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1127), .B(new_n1128), .C1(new_n1142), .C2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1207), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1178), .A2(new_n1196), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1146), .B2(new_n1123), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n705), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1214), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1188), .A2(new_n773), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n764), .B1(new_n1148), .B2(G50), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n817), .A2(G132), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n839), .B2(new_n787), .C1(new_n791), .C2(new_n1158), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G150), .A2(new_n1060), .B1(new_n802), .B2(G125), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(G128), .C2(new_n798), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n336), .B(new_n283), .C1(new_n789), .C2(new_n782), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G124), .B2(new_n815), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G97), .A2(new_n817), .B1(new_n808), .B2(new_n360), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT121), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n427), .A2(new_n283), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n792), .B2(G77), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n208), .B2(new_n789), .C1(new_n828), .C2(new_n781), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1018), .B1(G107), .B2(new_n798), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n574), .B2(new_n805), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1236), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT58), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1237), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1242), .A2(KEYINPUT58), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1234), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1223), .B1(new_n1246), .B2(new_n772), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1222), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1211), .B2(new_n762), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1221), .A2(new_n1250), .ZN(G375));
  XNOR2_X1  g1051(.A(new_n761), .B(KEYINPUT124), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1113), .A2(new_n773), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n765), .B1(G68), .B2(new_n1148), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G116), .A2(new_n817), .B1(new_n815), .B2(G303), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1256), .B1(new_n210), .B2(new_n791), .C1(new_n368), .C2(new_n787), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G283), .A2(new_n798), .B1(new_n802), .B2(G294), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n292), .B1(new_n819), .B2(G77), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(new_n361), .C2(new_n795), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G50), .A2(new_n1060), .B1(new_n798), .B2(G137), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n427), .B1(new_n819), .B2(G58), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n843), .C2(new_n805), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n792), .A2(G159), .B1(new_n815), .B2(G128), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n808), .A2(G150), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n800), .C2(new_n1158), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1257), .A2(new_n1260), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1255), .B1(new_n772), .B2(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1123), .A2(new_n1253), .B1(new_n1254), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1009), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1129), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1123), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1269), .B1(new_n1271), .B2(new_n1272), .ZN(G381));
  INV_X1    g1073(.A(G387), .ZN(new_n1274));
  INV_X1    g1074(.A(G378), .ZN(new_n1275));
  INV_X1    g1075(.A(G375), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1044), .A2(new_n826), .A3(new_n1077), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(G390), .A2(new_n1277), .A3(G384), .A4(G381), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1278), .ZN(G407));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n684), .A3(new_n1275), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G407), .A2(G213), .A3(new_n1280), .ZN(G409));
  AOI21_X1  g1081(.A(new_n826), .B1(new_n1044), .B2(new_n1077), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(G390), .A3(new_n1277), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1277), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1082), .B(new_n1106), .C1(new_n1285), .C2(new_n1282), .ZN(new_n1286));
  AND4_X1   g1086(.A1(new_n1013), .A2(new_n1038), .A3(new_n1284), .A4(new_n1286), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1013), .A2(new_n1038), .B1(new_n1286), .B2(new_n1284), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G378), .B(new_n1250), .C1(new_n1214), .C2(new_n1220), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1009), .B(new_n1219), .C1(new_n1201), .C2(new_n1210), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1253), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1248), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1275), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G213), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(G343), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1272), .B1(KEYINPUT60), .B2(new_n1129), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1218), .A2(new_n1212), .A3(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n705), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1269), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(G384), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G384), .B(new_n1269), .C1(new_n1300), .C2(new_n1302), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1296), .A2(new_n1299), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1298), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1298), .A2(G2897), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1305), .A2(new_n1306), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1311), .B(new_n1312), .C1(new_n1313), .C2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1313), .A2(new_n1320), .A3(new_n1308), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1310), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1318), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1311), .B1(new_n1325), .B2(new_n1312), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1290), .B1(new_n1322), .B2(new_n1326), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1287), .A2(new_n1288), .A3(KEYINPUT61), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1309), .A2(KEYINPUT125), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT63), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1309), .A2(KEYINPUT125), .A3(new_n1331), .ZN(new_n1332));
  OR2_X1    g1132(.A1(new_n1318), .A2(KEYINPUT126), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1318), .A2(KEYINPUT126), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1333), .A2(new_n1323), .A3(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1328), .A2(new_n1330), .A3(new_n1332), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1327), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1275), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1291), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1308), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1338), .A2(new_n1291), .A3(new_n1307), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1290), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1340), .A2(new_n1289), .A3(new_n1341), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(G402));
endmodule


