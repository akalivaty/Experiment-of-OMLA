

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729;

  NOR2_X1 U367 ( .A1(n716), .A2(n605), .ZN(n443) );
  NAND2_X1 U368 ( .A1(n407), .A2(n406), .ZN(n445) );
  NOR2_X1 U369 ( .A1(n577), .A2(n578), .ZN(n456) );
  BUF_X1 U370 ( .A(n538), .Z(n346) );
  NAND2_X1 U371 ( .A1(n538), .A2(n640), .ZN(n551) );
  NOR2_X1 U372 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U373 ( .A(n584), .B(KEYINPUT1), .ZN(n538) );
  BUF_X1 U374 ( .A(n571), .Z(n638) );
  OR2_X1 U375 ( .A1(n685), .A2(G902), .ZN(n392) );
  XNOR2_X1 U376 ( .A(n528), .B(n459), .ZN(n685) );
  XNOR2_X1 U377 ( .A(n528), .B(n452), .ZN(n531) );
  XOR2_X1 U378 ( .A(KEYINPUT69), .B(G131), .Z(n487) );
  XNOR2_X2 U379 ( .A(n604), .B(KEYINPUT84), .ZN(n716) );
  XNOR2_X2 U380 ( .A(n715), .B(G146), .ZN(n528) );
  AND2_X2 U381 ( .A1(n442), .A2(n365), .ZN(n441) );
  XNOR2_X2 U382 ( .A(n345), .B(KEYINPUT75), .ZN(n670) );
  NAND2_X1 U383 ( .A1(n451), .A2(n349), .ZN(n345) );
  INV_X1 U384 ( .A(G953), .ZN(n717) );
  NOR2_X1 U385 ( .A1(n728), .A2(n729), .ZN(n449) );
  NOR2_X2 U386 ( .A1(n673), .A2(n554), .ZN(n400) );
  AND2_X1 U387 ( .A1(n536), .A2(n552), .ZN(n371) );
  XNOR2_X1 U388 ( .A(n503), .B(n360), .ZN(n594) );
  XOR2_X2 U389 ( .A(G122), .B(G104), .Z(n497) );
  XNOR2_X1 U390 ( .A(n551), .B(KEYINPUT107), .ZN(n387) );
  NOR2_X1 U391 ( .A1(n604), .A2(n603), .ZN(n451) );
  NOR2_X1 U392 ( .A1(n726), .A2(n383), .ZN(n382) );
  XNOR2_X1 U393 ( .A(n601), .B(n600), .ZN(n728) );
  XNOR2_X1 U394 ( .A(n435), .B(n434), .ZN(n729) );
  NOR2_X1 U395 ( .A1(n597), .A2(n598), .ZN(n408) );
  XNOR2_X1 U396 ( .A(n371), .B(n363), .ZN(n542) );
  XNOR2_X1 U397 ( .A(n534), .B(n533), .ZN(n673) );
  NAND2_X1 U398 ( .A1(n387), .A2(n568), .ZN(n534) );
  NOR2_X1 U399 ( .A1(n655), .A2(n654), .ZN(n436) );
  XOR2_X1 U400 ( .A(KEYINPUT6), .B(n638), .Z(n568) );
  XNOR2_X1 U401 ( .A(n468), .B(n467), .ZN(n496) );
  XNOR2_X1 U402 ( .A(n414), .B(G146), .ZN(n499) );
  INV_X1 U403 ( .A(KEYINPUT60), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(G60) );
  NAND2_X1 U405 ( .A1(n370), .A2(n369), .ZN(n348) );
  INV_X1 U406 ( .A(n349), .ZN(n704) );
  XNOR2_X2 U407 ( .A(n561), .B(n350), .ZN(n349) );
  XOR2_X1 U408 ( .A(KEYINPUT45), .B(KEYINPUT85), .Z(n350) );
  XOR2_X2 U409 ( .A(KEYINPUT38), .B(n398), .Z(n651) );
  NOR2_X2 U410 ( .A1(n416), .A2(n415), .ZN(n640) );
  XNOR2_X1 U411 ( .A(n656), .B(n374), .ZN(n589) );
  INV_X1 U412 ( .A(KEYINPUT81), .ZN(n374) );
  XNOR2_X1 U413 ( .A(n469), .B(G137), .ZN(n454) );
  XOR2_X1 U414 ( .A(G107), .B(G110), .Z(n524) );
  INV_X1 U415 ( .A(G113), .ZN(n465) );
  INV_X1 U416 ( .A(KEYINPUT44), .ZN(n380) );
  XNOR2_X1 U417 ( .A(G110), .B(KEYINPUT76), .ZN(n511) );
  INV_X1 U418 ( .A(G125), .ZN(n414) );
  XOR2_X1 U419 ( .A(G137), .B(G140), .Z(n530) );
  XNOR2_X1 U420 ( .A(G104), .B(G101), .ZN(n529) );
  XNOR2_X1 U421 ( .A(n399), .B(G472), .ZN(n571) );
  OR2_X1 U422 ( .A1(n531), .A2(G902), .ZN(n399) );
  XNOR2_X1 U423 ( .A(n489), .B(n433), .ZN(n547) );
  XNOR2_X1 U424 ( .A(n490), .B(G475), .ZN(n433) );
  NOR2_X1 U425 ( .A1(G902), .A2(n692), .ZN(n489) );
  AND2_X1 U426 ( .A1(n422), .A2(n421), .ZN(n420) );
  NAND2_X1 U427 ( .A1(n423), .A2(G902), .ZN(n421) );
  OR2_X1 U428 ( .A1(n698), .A2(n418), .ZN(n417) );
  INV_X1 U429 ( .A(G902), .ZN(n419) );
  INV_X1 U430 ( .A(n650), .ZN(n457) );
  XNOR2_X1 U431 ( .A(n436), .B(n595), .ZN(n675) );
  INV_X1 U432 ( .A(KEYINPUT0), .ZN(n506) );
  NAND2_X1 U433 ( .A1(n420), .A2(n417), .ZN(n633) );
  XNOR2_X1 U434 ( .A(n384), .B(n473), .ZN(n476) );
  NOR2_X1 U435 ( .A1(n355), .A2(n351), .ZN(n450) );
  INV_X1 U436 ( .A(KEYINPUT48), .ZN(n440) );
  OR2_X1 U437 ( .A1(G902), .A2(G237), .ZN(n504) );
  INV_X1 U438 ( .A(KEYINPUT25), .ZN(n519) );
  NOR2_X1 U439 ( .A1(G953), .A2(G237), .ZN(n482) );
  NAND2_X1 U440 ( .A1(n386), .A2(n438), .ZN(n604) );
  NOR2_X1 U441 ( .A1(n632), .A2(n439), .ZN(n438) );
  XNOR2_X1 U442 ( .A(n373), .B(n440), .ZN(n386) );
  INV_X1 U443 ( .A(n631), .ZN(n439) );
  NAND2_X1 U444 ( .A1(G224), .A2(n717), .ZN(n502) );
  INV_X1 U445 ( .A(KEYINPUT88), .ZN(n448) );
  XNOR2_X1 U446 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U447 ( .A(KEYINPUT4), .ZN(n462) );
  XNOR2_X1 U448 ( .A(n550), .B(n375), .ZN(n656) );
  INV_X1 U449 ( .A(KEYINPUT103), .ZN(n375) );
  XNOR2_X1 U450 ( .A(n432), .B(KEYINPUT104), .ZN(n654) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n582) );
  INV_X1 U452 ( .A(KEYINPUT70), .ZN(n396) );
  AND2_X1 U453 ( .A1(n633), .A2(n357), .ZN(n397) );
  INV_X1 U454 ( .A(n420), .ZN(n415) );
  XNOR2_X1 U455 ( .A(n496), .B(n453), .ZN(n452) );
  XNOR2_X1 U456 ( .A(n454), .B(n354), .ZN(n453) );
  XNOR2_X1 U457 ( .A(n437), .B(n496), .ZN(n707) );
  XNOR2_X1 U458 ( .A(n378), .B(n524), .ZN(n437) );
  XNOR2_X1 U459 ( .A(n497), .B(n379), .ZN(n378) );
  INV_X1 U460 ( .A(KEYINPUT16), .ZN(n379) );
  XNOR2_X1 U461 ( .A(n508), .B(n530), .ZN(n713) );
  XOR2_X1 U462 ( .A(KEYINPUT97), .B(KEYINPUT24), .Z(n512) );
  XOR2_X1 U463 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n478) );
  XNOR2_X1 U464 ( .A(n472), .B(n385), .ZN(n384) );
  INV_X1 U465 ( .A(G134), .ZN(n385) );
  XNOR2_X1 U466 ( .A(G122), .B(G116), .ZN(n472) );
  XOR2_X1 U467 ( .A(KEYINPUT7), .B(G107), .Z(n473) );
  XNOR2_X1 U468 ( .A(n499), .B(KEYINPUT10), .ZN(n508) );
  XNOR2_X1 U469 ( .A(n527), .B(n460), .ZN(n459) );
  XNOR2_X1 U470 ( .A(n530), .B(n529), .ZN(n460) );
  XNOR2_X1 U471 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U472 ( .A(n446), .B(n707), .ZN(n681) );
  XNOR2_X1 U473 ( .A(n501), .B(n425), .ZN(n446) );
  XNOR2_X1 U474 ( .A(n447), .B(n500), .ZN(n425) );
  XNOR2_X1 U475 ( .A(n502), .B(n448), .ZN(n447) );
  BUF_X1 U476 ( .A(n673), .Z(n391) );
  AND2_X1 U477 ( .A1(n538), .A2(n633), .ZN(n541) );
  INV_X1 U478 ( .A(KEYINPUT78), .ZN(n390) );
  XNOR2_X1 U479 ( .A(n424), .B(KEYINPUT19), .ZN(n586) );
  NAND2_X1 U480 ( .A1(n594), .A2(n650), .ZN(n424) );
  NOR2_X1 U481 ( .A1(n572), .A2(n410), .ZN(n409) );
  INV_X1 U482 ( .A(n573), .ZN(n411) );
  INV_X1 U483 ( .A(n574), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n376), .B(KEYINPUT98), .ZN(n573) );
  NAND2_X1 U485 ( .A1(n584), .A2(n640), .ZN(n376) );
  INV_X1 U486 ( .A(KEYINPUT96), .ZN(n507) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n692) );
  XNOR2_X1 U488 ( .A(n488), .B(n428), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n359), .B(n508), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n485), .B(n483), .ZN(n428) );
  INV_X1 U491 ( .A(KEYINPUT42), .ZN(n434) );
  INV_X1 U492 ( .A(KEYINPUT35), .ZN(n444) );
  XNOR2_X1 U493 ( .A(n430), .B(n372), .ZN(n726) );
  XNOR2_X1 U494 ( .A(n429), .B(n390), .ZN(n372) );
  NOR2_X1 U495 ( .A1(n542), .A2(n431), .ZN(n430) );
  INV_X1 U496 ( .A(KEYINPUT32), .ZN(n429) );
  AND2_X1 U497 ( .A1(n596), .A2(n586), .ZN(n622) );
  XNOR2_X1 U498 ( .A(KEYINPUT106), .B(n540), .ZN(n727) );
  NOR2_X1 U499 ( .A1(n549), .A2(n548), .ZN(n624) );
  XNOR2_X1 U500 ( .A(n694), .B(n402), .ZN(n401) );
  INV_X1 U501 ( .A(n695), .ZN(n402) );
  XNOR2_X1 U502 ( .A(G902), .B(KEYINPUT15), .ZN(n605) );
  XOR2_X1 U503 ( .A(KEYINPUT82), .B(n620), .Z(n351) );
  AND2_X1 U504 ( .A1(n624), .A2(n568), .ZN(n352) );
  XOR2_X1 U505 ( .A(G134), .B(n487), .Z(n353) );
  XNOR2_X1 U506 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n354) );
  AND2_X1 U507 ( .A1(n593), .A2(KEYINPUT47), .ZN(n355) );
  XOR2_X1 U508 ( .A(KEYINPUT71), .B(G469), .Z(n356) );
  AND2_X1 U509 ( .A1(n574), .A2(n566), .ZN(n357) );
  XOR2_X1 U510 ( .A(n541), .B(KEYINPUT105), .Z(n358) );
  XOR2_X1 U511 ( .A(n484), .B(n486), .Z(n359) );
  AND2_X1 U512 ( .A1(G210), .A2(n504), .ZN(n360) );
  NOR2_X1 U513 ( .A1(n582), .A2(n457), .ZN(n361) );
  XOR2_X1 U514 ( .A(KEYINPUT34), .B(KEYINPUT77), .Z(n362) );
  XOR2_X1 U515 ( .A(n537), .B(KEYINPUT65), .Z(n363) );
  XOR2_X1 U516 ( .A(n471), .B(n470), .Z(n364) );
  XNOR2_X1 U517 ( .A(KEYINPUT66), .B(n607), .ZN(n365) );
  XOR2_X1 U518 ( .A(n692), .B(n691), .Z(n366) );
  NOR2_X1 U519 ( .A1(G952), .A2(n717), .ZN(n700) );
  INV_X1 U520 ( .A(n700), .ZN(n369) );
  XOR2_X1 U521 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n367) );
  XOR2_X1 U522 ( .A(KEYINPUT86), .B(KEYINPUT56), .Z(n368) );
  NAND2_X1 U523 ( .A1(n725), .A2(n382), .ZN(n381) );
  XNOR2_X2 U524 ( .A(n445), .B(n444), .ZN(n725) );
  XNOR2_X1 U525 ( .A(n693), .B(n366), .ZN(n370) );
  XNOR2_X1 U526 ( .A(n475), .B(n476), .ZN(n480) );
  XOR2_X1 U527 ( .A(G478), .B(n481), .Z(n549) );
  NAND2_X1 U528 ( .A1(n535), .A2(n547), .ZN(n432) );
  NAND2_X1 U529 ( .A1(n696), .A2(G475), .ZN(n693) );
  NOR2_X4 U530 ( .A1(n441), .A2(n670), .ZN(n696) );
  INV_X1 U531 ( .A(n521), .ZN(n423) );
  NAND2_X1 U532 ( .A1(n521), .A2(n419), .ZN(n418) );
  XNOR2_X1 U533 ( .A(n381), .B(n380), .ZN(n560) );
  XNOR2_X1 U534 ( .A(n394), .B(KEYINPUT30), .ZN(n572) );
  NAND2_X1 U535 ( .A1(n413), .A2(n412), .ZN(n373) );
  AND2_X1 U536 ( .A1(n591), .A2(n450), .ZN(n412) );
  XNOR2_X1 U537 ( .A(n408), .B(n599), .ZN(n602) );
  XNOR2_X2 U538 ( .A(n377), .B(n506), .ZN(n552) );
  NAND2_X1 U539 ( .A1(n586), .A2(n505), .ZN(n377) );
  INV_X1 U540 ( .A(n727), .ZN(n383) );
  NAND2_X1 U541 ( .A1(n596), .A2(n675), .ZN(n435) );
  NAND2_X1 U542 ( .A1(n409), .A2(n411), .ZN(n597) );
  INV_X1 U543 ( .A(n575), .ZN(n406) );
  XNOR2_X1 U544 ( .A(n389), .B(n367), .ZN(G57) );
  NAND2_X1 U545 ( .A1(n395), .A2(n369), .ZN(n389) );
  NOR2_X2 U546 ( .A1(n542), .A2(n346), .ZN(n545) );
  XNOR2_X2 U547 ( .A(n392), .B(n356), .ZN(n584) );
  XNOR2_X1 U548 ( .A(n393), .B(n368), .ZN(G51) );
  NAND2_X1 U549 ( .A1(n684), .A2(n369), .ZN(n393) );
  NAND2_X1 U550 ( .A1(n571), .A2(n650), .ZN(n394) );
  XNOR2_X1 U551 ( .A(n608), .B(n364), .ZN(n395) );
  XNOR2_X1 U552 ( .A(n583), .B(KEYINPUT28), .ZN(n585) );
  BUF_X2 U553 ( .A(n594), .Z(n398) );
  XNOR2_X1 U554 ( .A(n400), .B(n362), .ZN(n407) );
  NAND2_X1 U555 ( .A1(n401), .A2(n369), .ZN(n405) );
  NAND2_X1 U556 ( .A1(n403), .A2(n676), .ZN(n677) );
  NAND2_X1 U557 ( .A1(n671), .A2(n672), .ZN(n403) );
  XNOR2_X1 U558 ( .A(n404), .B(KEYINPUT53), .ZN(G75) );
  AND2_X1 U559 ( .A1(n679), .A2(n717), .ZN(n404) );
  NAND2_X1 U560 ( .A1(n696), .A2(G478), .ZN(n694) );
  XNOR2_X1 U561 ( .A(n405), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U562 ( .A(n449), .B(KEYINPUT46), .ZN(n413) );
  NAND2_X1 U563 ( .A1(n417), .A2(n566), .ZN(n416) );
  NAND2_X1 U564 ( .A1(n698), .A2(n423), .ZN(n422) );
  XNOR2_X1 U565 ( .A(n517), .B(n516), .ZN(n698) );
  XNOR2_X2 U566 ( .A(n474), .B(n462), .ZN(n501) );
  XNOR2_X2 U567 ( .A(n458), .B(G143), .ZN(n474) );
  NAND2_X1 U568 ( .A1(n543), .A2(n358), .ZN(n431) );
  NAND2_X1 U569 ( .A1(n443), .A2(n349), .ZN(n442) );
  INV_X1 U570 ( .A(n398), .ZN(n578) );
  XNOR2_X2 U571 ( .A(n501), .B(n353), .ZN(n715) );
  XNOR2_X1 U572 ( .A(n456), .B(n455), .ZN(n579) );
  INV_X1 U573 ( .A(KEYINPUT36), .ZN(n455) );
  NAND2_X1 U574 ( .A1(n352), .A2(n361), .ZN(n577) );
  XNOR2_X2 U575 ( .A(G128), .B(KEYINPUT64), .ZN(n458) );
  AND2_X1 U576 ( .A1(G221), .A2(n509), .ZN(n461) );
  XNOR2_X1 U577 ( .A(n466), .B(n465), .ZN(n467) );
  INV_X1 U578 ( .A(KEYINPUT23), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n532), .B(KEYINPUT108), .ZN(n533) );
  XNOR2_X1 U580 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n552), .B(n507), .ZN(n554) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n713), .B(n461), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(n521) );
  INV_X1 U585 ( .A(KEYINPUT40), .ZN(n600) );
  XOR2_X1 U586 ( .A(KEYINPUT62), .B(KEYINPUT89), .Z(n471) );
  XOR2_X1 U587 ( .A(G119), .B(KEYINPUT92), .Z(n464) );
  XNOR2_X1 U588 ( .A(KEYINPUT3), .B(KEYINPUT72), .ZN(n463) );
  XNOR2_X1 U589 ( .A(n464), .B(n463), .ZN(n468) );
  XNOR2_X1 U590 ( .A(G116), .B(G101), .ZN(n466) );
  NAND2_X1 U591 ( .A1(n482), .A2(G210), .ZN(n469) );
  XNOR2_X1 U592 ( .A(n531), .B(KEYINPUT110), .ZN(n470) );
  XNOR2_X1 U593 ( .A(n474), .B(KEYINPUT9), .ZN(n475) );
  NAND2_X1 U594 ( .A1(G234), .A2(n717), .ZN(n477) );
  XNOR2_X1 U595 ( .A(n478), .B(n477), .ZN(n509) );
  NAND2_X1 U596 ( .A1(G217), .A2(n509), .ZN(n479) );
  XNOR2_X1 U597 ( .A(n480), .B(n479), .ZN(n695) );
  NOR2_X1 U598 ( .A1(n695), .A2(G902), .ZN(n481) );
  INV_X1 U599 ( .A(n549), .ZN(n535) );
  XNOR2_X1 U600 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n490) );
  XOR2_X1 U601 ( .A(G140), .B(KEYINPUT11), .Z(n484) );
  NAND2_X1 U602 ( .A1(n482), .A2(G214), .ZN(n483) );
  XOR2_X1 U603 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n486) );
  XNOR2_X1 U604 ( .A(G143), .B(G113), .ZN(n485) );
  XNOR2_X1 U605 ( .A(n497), .B(n487), .ZN(n488) );
  OR2_X1 U606 ( .A1(n535), .A2(n547), .ZN(n575) );
  NAND2_X1 U607 ( .A1(G237), .A2(G234), .ZN(n491) );
  XNOR2_X1 U608 ( .A(n491), .B(KEYINPUT14), .ZN(n493) );
  NAND2_X1 U609 ( .A1(G902), .A2(n493), .ZN(n562) );
  XOR2_X1 U610 ( .A(G898), .B(KEYINPUT94), .Z(n703) );
  NAND2_X1 U611 ( .A1(G953), .A2(n703), .ZN(n708) );
  NOR2_X1 U612 ( .A1(n562), .A2(n708), .ZN(n492) );
  XNOR2_X1 U613 ( .A(KEYINPUT95), .B(n492), .ZN(n495) );
  NAND2_X1 U614 ( .A1(G952), .A2(n493), .ZN(n666) );
  NOR2_X1 U615 ( .A1(n666), .A2(G953), .ZN(n494) );
  XNOR2_X1 U616 ( .A(n494), .B(KEYINPUT93), .ZN(n565) );
  NAND2_X1 U617 ( .A1(n495), .A2(n565), .ZN(n505) );
  XOR2_X1 U618 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n498) );
  NAND2_X1 U619 ( .A1(n605), .A2(n681), .ZN(n503) );
  NAND2_X1 U620 ( .A1(G214), .A2(n504), .ZN(n650) );
  XNOR2_X1 U621 ( .A(G128), .B(G119), .ZN(n514) );
  XNOR2_X1 U622 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U623 ( .A1(n605), .A2(G234), .ZN(n518) );
  XNOR2_X1 U624 ( .A(n518), .B(KEYINPUT20), .ZN(n522) );
  NAND2_X1 U625 ( .A1(n522), .A2(G217), .ZN(n520) );
  NAND2_X1 U626 ( .A1(G221), .A2(n522), .ZN(n523) );
  XOR2_X1 U627 ( .A(KEYINPUT21), .B(n523), .Z(n566) );
  INV_X1 U628 ( .A(n566), .ZN(n634) );
  INV_X1 U629 ( .A(n524), .ZN(n526) );
  NAND2_X1 U630 ( .A1(G227), .A2(n717), .ZN(n525) );
  INV_X1 U631 ( .A(KEYINPUT33), .ZN(n532) );
  NOR2_X1 U632 ( .A1(n634), .A2(n654), .ZN(n536) );
  XNOR2_X1 U633 ( .A(KEYINPUT22), .B(KEYINPUT73), .ZN(n537) );
  INV_X1 U634 ( .A(n633), .ZN(n567) );
  NOR2_X1 U635 ( .A1(n567), .A2(n638), .ZN(n539) );
  NAND2_X1 U636 ( .A1(n545), .A2(n539), .ZN(n540) );
  INV_X1 U637 ( .A(n568), .ZN(n544) );
  XOR2_X1 U638 ( .A(n544), .B(KEYINPUT79), .Z(n543) );
  INV_X1 U639 ( .A(n346), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U641 ( .A1(n633), .A2(n546), .ZN(n609) );
  XNOR2_X1 U642 ( .A(KEYINPUT102), .B(n547), .ZN(n548) );
  AND2_X1 U643 ( .A1(n549), .A2(n548), .ZN(n626) );
  NOR2_X1 U644 ( .A1(n626), .A2(n624), .ZN(n550) );
  INV_X1 U645 ( .A(n638), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n581), .A2(n551), .ZN(n646) );
  NAND2_X1 U647 ( .A1(n552), .A2(n646), .ZN(n553) );
  XNOR2_X1 U648 ( .A(n553), .B(KEYINPUT31), .ZN(n627) );
  NOR2_X1 U649 ( .A1(n573), .A2(n554), .ZN(n555) );
  NAND2_X1 U650 ( .A1(n555), .A2(n581), .ZN(n556) );
  XNOR2_X1 U651 ( .A(KEYINPUT99), .B(n556), .ZN(n612) );
  NOR2_X1 U652 ( .A1(n627), .A2(n612), .ZN(n557) );
  NOR2_X1 U653 ( .A1(n589), .A2(n557), .ZN(n558) );
  NOR2_X1 U654 ( .A1(n609), .A2(n558), .ZN(n559) );
  NAND2_X1 U655 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U656 ( .A1(G900), .A2(n562), .ZN(n563) );
  NAND2_X1 U657 ( .A1(G953), .A2(n563), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n565), .A2(n564), .ZN(n574) );
  NOR2_X1 U659 ( .A1(n346), .A2(n577), .ZN(n569) );
  XNOR2_X1 U660 ( .A(n569), .B(KEYINPUT43), .ZN(n570) );
  NOR2_X1 U661 ( .A1(n398), .A2(n570), .ZN(n632) );
  NOR2_X1 U662 ( .A1(n597), .A2(n575), .ZN(n576) );
  NAND2_X1 U663 ( .A1(n398), .A2(n576), .ZN(n620) );
  NOR2_X1 U664 ( .A1(n580), .A2(n579), .ZN(n629) );
  XNOR2_X1 U665 ( .A(KEYINPUT47), .B(KEYINPUT67), .ZN(n587) );
  AND2_X1 U666 ( .A1(n584), .A2(n585), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n587), .A2(n622), .ZN(n588) );
  NOR2_X1 U668 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U669 ( .A1(n629), .A2(n590), .ZN(n591) );
  INV_X1 U670 ( .A(n656), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n592), .A2(n622), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n651), .A2(n650), .ZN(n655) );
  XNOR2_X1 U673 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n595) );
  INV_X1 U674 ( .A(n651), .ZN(n598) );
  XNOR2_X1 U675 ( .A(KEYINPUT87), .B(KEYINPUT39), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n602), .A2(n624), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n626), .ZN(n631) );
  INV_X1 U678 ( .A(KEYINPUT2), .ZN(n603) );
  INV_X1 U679 ( .A(n605), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n606), .A2(KEYINPUT2), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n696), .A2(G472), .ZN(n608) );
  XOR2_X1 U682 ( .A(G101), .B(n609), .Z(G3) );
  XOR2_X1 U683 ( .A(G104), .B(KEYINPUT111), .Z(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n624), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(G6) );
  XOR2_X1 U686 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n614) );
  NAND2_X1 U687 ( .A1(n612), .A2(n626), .ZN(n613) );
  XNOR2_X1 U688 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U689 ( .A(G107), .B(n615), .ZN(G9) );
  XOR2_X1 U690 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n617) );
  NAND2_X1 U691 ( .A1(n622), .A2(n626), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n617), .B(n616), .ZN(n619) );
  XOR2_X1 U693 ( .A(G128), .B(KEYINPUT112), .Z(n618) );
  XNOR2_X1 U694 ( .A(n619), .B(n618), .ZN(G30) );
  XNOR2_X1 U695 ( .A(G143), .B(KEYINPUT114), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n621), .B(n620), .ZN(G45) );
  NAND2_X1 U697 ( .A1(n622), .A2(n624), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(G146), .ZN(G48) );
  NAND2_X1 U699 ( .A1(n627), .A2(n624), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n625), .B(G113), .ZN(G15) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n628), .B(G116), .ZN(G18) );
  XNOR2_X1 U703 ( .A(n629), .B(G125), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U705 ( .A(G134), .B(n631), .ZN(G36) );
  XOR2_X1 U706 ( .A(G140), .B(n632), .Z(G42) );
  XNOR2_X1 U707 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n648) );
  XOR2_X1 U708 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n636) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U712 ( .A(KEYINPUT116), .B(n639), .Z(n644) );
  NOR2_X1 U713 ( .A1(n640), .A2(n346), .ZN(n641) );
  XOR2_X1 U714 ( .A(KEYINPUT117), .B(n641), .Z(n642) );
  XNOR2_X1 U715 ( .A(KEYINPUT50), .B(n642), .ZN(n643) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n649), .A2(n675), .ZN(n662) );
  NOR2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U721 ( .A(KEYINPUT119), .B(n652), .Z(n653) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n658) );
  NOR2_X1 U723 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U725 ( .A1(n391), .A2(n659), .ZN(n660) );
  XOR2_X1 U726 ( .A(KEYINPUT120), .B(n660), .Z(n661) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U728 ( .A(n663), .B(KEYINPUT121), .ZN(n664) );
  XNOR2_X1 U729 ( .A(n664), .B(KEYINPUT52), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n678) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n667) );
  NAND2_X1 U732 ( .A1(n704), .A2(n667), .ZN(n672) );
  NAND2_X1 U733 ( .A1(n716), .A2(n667), .ZN(n668) );
  XNOR2_X1 U734 ( .A(KEYINPUT83), .B(n668), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  INV_X1 U736 ( .A(n391), .ZN(n674) );
  NAND2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U739 ( .A1(n696), .A2(G210), .ZN(n683) );
  XOR2_X1 U740 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n680) );
  XNOR2_X1 U741 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U742 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U743 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n687) );
  XNOR2_X1 U744 ( .A(n685), .B(KEYINPUT57), .ZN(n686) );
  XNOR2_X1 U745 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U746 ( .A1(n696), .A2(G469), .ZN(n688) );
  XOR2_X1 U747 ( .A(n689), .B(n688), .Z(n690) );
  NOR2_X1 U748 ( .A1(n700), .A2(n690), .ZN(G54) );
  XOR2_X1 U749 ( .A(KEYINPUT59), .B(KEYINPUT90), .Z(n691) );
  NAND2_X1 U750 ( .A1(G217), .A2(n696), .ZN(n697) );
  XNOR2_X1 U751 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U752 ( .A1(n700), .A2(n699), .ZN(G66) );
  NAND2_X1 U753 ( .A1(G953), .A2(G224), .ZN(n701) );
  XOR2_X1 U754 ( .A(KEYINPUT61), .B(n701), .Z(n702) );
  NOR2_X1 U755 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U756 ( .A1(G953), .A2(n704), .ZN(n705) );
  NOR2_X1 U757 ( .A1(n706), .A2(n705), .ZN(n712) );
  XNOR2_X1 U758 ( .A(n707), .B(KEYINPUT124), .ZN(n709) );
  NAND2_X1 U759 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U760 ( .A(n710), .B(KEYINPUT125), .ZN(n711) );
  XOR2_X1 U761 ( .A(n712), .B(n711), .Z(G69) );
  XOR2_X1 U762 ( .A(n713), .B(KEYINPUT126), .Z(n714) );
  XNOR2_X1 U763 ( .A(n715), .B(n714), .ZN(n719) );
  XNOR2_X1 U764 ( .A(n716), .B(n719), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n718), .A2(n717), .ZN(n724) );
  XNOR2_X1 U766 ( .A(G227), .B(n719), .ZN(n720) );
  NAND2_X1 U767 ( .A1(n720), .A2(G900), .ZN(n721) );
  NAND2_X1 U768 ( .A1(n721), .A2(G953), .ZN(n722) );
  XOR2_X1 U769 ( .A(KEYINPUT127), .B(n722), .Z(n723) );
  NAND2_X1 U770 ( .A1(n724), .A2(n723), .ZN(G72) );
  XNOR2_X1 U771 ( .A(n725), .B(G122), .ZN(G24) );
  XOR2_X1 U772 ( .A(n726), .B(G119), .Z(G21) );
  XNOR2_X1 U773 ( .A(n727), .B(G110), .ZN(G12) );
  XOR2_X1 U774 ( .A(n728), .B(G131), .Z(G33) );
  XOR2_X1 U775 ( .A(G137), .B(n729), .Z(G39) );
endmodule

