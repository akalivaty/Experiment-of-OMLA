//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G120gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G134gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(G127gat), .ZN(new_n210));
  INV_X1    g009(.A(G127gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n207), .B(new_n209), .C1(KEYINPUT68), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(KEYINPUT70), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT69), .B1(new_n203), .B2(G120gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(new_n205), .A3(G113gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n203), .A2(G120gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n210), .A2(new_n212), .A3(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n215), .A2(new_n220), .A3(new_n202), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n232), .A2(KEYINPUT23), .B1(new_n233), .B2(KEYINPUT65), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G169gat), .A3(G176gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n231), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  INV_X1    g039(.A(G190gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n242), .B(new_n245), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT24), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n240), .A2(new_n241), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n244), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n232), .A2(KEYINPUT23), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n230), .B1(G169gat), .B2(G176gat), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .A4(new_n233), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n238), .A2(new_n250), .B1(new_n258), .B2(new_n226), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT27), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G183gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(new_n241), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT27), .B(G183gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT28), .A3(new_n241), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n232), .A2(KEYINPUT26), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT26), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(G169gat), .B2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n272), .A2(new_n233), .B1(G183gat), .B2(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n225), .B1(new_n259), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT64), .ZN(new_n278));
  INV_X1    g077(.A(new_n255), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n257), .A3(new_n233), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n226), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n242), .A2(new_n244), .A3(new_n243), .ZN(new_n282));
  INV_X1    g081(.A(new_n249), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(new_n247), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n281), .B1(new_n284), .B2(new_n237), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n274), .A3(new_n224), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT33), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G15gat), .B(G43gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT72), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G71gat), .B(G99gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n293), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n293), .B2(new_n297), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n290), .A3(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n287), .B(KEYINPUT32), .C1(new_n289), .C2(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n278), .B1(new_n276), .B2(new_n286), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT34), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI211_X1 g108(.A(KEYINPUT34), .B(new_n278), .C1(new_n276), .C2(new_n286), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n309), .A2(new_n310), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(new_n304), .A3(new_n305), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT36), .ZN(new_n316));
  XNOR2_X1  g115(.A(G1gat), .B(G29gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT0), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n318), .B(KEYINPUT77), .Z(new_n319));
  XOR2_X1   g118(.A(G57gat), .B(G85gat), .Z(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT78), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n319), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT5), .ZN(new_n323));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325));
  XOR2_X1   g124(.A(G155gat), .B(G162gat), .Z(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G141gat), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G148gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n328), .A2(new_n330), .B1(KEYINPUT2), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n326), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(KEYINPUT2), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n329), .A2(G148gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n327), .A2(G141gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G155gat), .B(G162gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n333), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n225), .A2(new_n325), .A3(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n332), .A2(new_n326), .A3(new_n334), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n339), .B2(new_n333), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT4), .B1(new_n346), .B2(new_n224), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT75), .B(KEYINPUT3), .Z(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n344), .B2(new_n345), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n341), .A3(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n224), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n342), .A2(new_n349), .B1(new_n214), .B2(new_n223), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT76), .B1(new_n355), .B2(new_n351), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n324), .B(new_n348), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n224), .B(new_n342), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n324), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n323), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n352), .A2(new_n353), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n355), .A2(KEYINPUT76), .A3(new_n351), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n362), .A2(new_n363), .B1(new_n347), .B2(new_n343), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT5), .B1(new_n364), .B2(new_n324), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n322), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n322), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n323), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n359), .B1(new_n364), .B2(new_n324), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(new_n323), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n366), .A2(new_n370), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n361), .A2(new_n365), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n374), .B(new_n367), .C1(KEYINPUT79), .C2(KEYINPUT6), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G211gat), .A2(G218gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G204gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G197gat), .ZN(new_n381));
  INV_X1    g180(.A(G197gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G204gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(G211gat), .A2(G218gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT73), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n377), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n384), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G226gat), .ZN(new_n389));
  INV_X1    g188(.A(G233gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n285), .A2(new_n274), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n238), .A2(new_n250), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n395), .A2(new_n281), .B1(new_n268), .B2(new_n273), .ZN(new_n396));
  INV_X1    g195(.A(new_n391), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n388), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n396), .B2(KEYINPUT29), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n392), .A2(new_n391), .ZN(new_n401));
  INV_X1    g200(.A(new_n388), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT30), .ZN(new_n404));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n399), .A2(new_n403), .A3(new_n404), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n399), .A2(new_n403), .A3(new_n408), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n399), .B2(new_n403), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n376), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n415));
  INV_X1    g214(.A(new_n349), .ZN(new_n416));
  XOR2_X1   g215(.A(G211gat), .B(G218gat), .Z(new_n417));
  NAND2_X1  g216(.A1(new_n384), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n385), .A2(new_n377), .ZN(new_n419));
  XNOR2_X1  g218(.A(G197gat), .B(G204gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n379), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n416), .B1(new_n422), .B2(new_n393), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n415), .B1(new_n423), .B2(new_n342), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n418), .B2(new_n421), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n346), .B(KEYINPUT81), .C1(new_n416), .C2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n416), .B1(new_n335), .B2(new_n341), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n388), .B1(new_n427), .B2(KEYINPUT29), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G228gat), .A2(G233gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n388), .B2(KEYINPUT29), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n433), .B2(new_n346), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n428), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G22gat), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n431), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT31), .B(G50gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT80), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n429), .A2(new_n430), .B1(new_n428), .B2(new_n434), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT83), .B1(new_n448), .B2(new_n438), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n443), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n436), .B2(G22gat), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n448), .A2(KEYINPUT82), .A3(new_n438), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n445), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n316), .B1(new_n414), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n348), .B1(new_n354), .B2(new_n356), .ZN(new_n458));
  INV_X1    g257(.A(new_n324), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT39), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n358), .B2(new_n324), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n367), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n461), .A3(new_n459), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT40), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n462), .B1(new_n364), .B2(new_n324), .ZN(new_n466));
  AND4_X1   g265(.A1(KEYINPUT40), .A2(new_n466), .A3(new_n464), .A4(new_n322), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n465), .A2(new_n413), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n370), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n357), .A2(new_n360), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT5), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n472), .A2(KEYINPUT84), .A3(new_n367), .A4(new_n368), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT85), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n466), .A2(new_n464), .A3(new_n322), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n412), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(KEYINPUT30), .A3(new_n410), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n466), .A2(new_n464), .A3(KEYINPUT40), .A4(new_n322), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n478), .A2(new_n480), .A3(new_n409), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n470), .A2(new_n473), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT85), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n470), .A2(new_n372), .A3(new_n366), .A4(new_n473), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n374), .A2(KEYINPUT6), .A3(new_n367), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n399), .A2(new_n403), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n407), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n490), .B1(new_n399), .B2(new_n403), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n494), .A2(new_n410), .ZN(new_n495));
  INV_X1    g294(.A(new_n399), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n496), .A2(KEYINPUT86), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n403), .B1(new_n496), .B2(KEYINPUT86), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT37), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n492), .A2(KEYINPUT38), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n455), .B1(new_n489), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n457), .B1(new_n486), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n315), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n455), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT35), .B1(new_n414), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n443), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n439), .A2(new_n446), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n448), .A2(KEYINPUT83), .A3(new_n438), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n436), .A2(new_n451), .A3(G22gat), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT82), .B1(new_n448), .B2(new_n438), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n315), .B1(new_n515), .B2(new_n445), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT35), .B1(new_n480), .B2(new_n409), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n489), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n504), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G190gat), .B(G218gat), .ZN(new_n521));
  INV_X1    g320(.A(G85gat), .ZN(new_n522));
  INV_X1    g321(.A(G92gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT90), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n524), .B(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(KEYINPUT90), .B2(new_n525), .ZN(new_n528));
  AND3_X1   g327(.A1(KEYINPUT91), .A2(G99gat), .A3(G106gat), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT91), .B1(G99gat), .B2(G106gat), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT8), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G99gat), .B(G106gat), .Z(new_n532));
  AOI22_X1  g331(.A1(new_n532), .A2(KEYINPUT92), .B1(new_n522), .B2(new_n523), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(KEYINPUT92), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n534), .A2(new_n535), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n535), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT93), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545));
  INV_X1    g344(.A(G50gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(G43gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n547), .B2(KEYINPUT87), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n549));
  INV_X1    g348(.A(G29gat), .ZN(new_n550));
  INV_X1    g349(.A(G36gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G29gat), .A2(G36gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G43gat), .B(G50gat), .Z(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT15), .B1(new_n554), .B2(new_n555), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(KEYINPUT17), .A3(new_n561), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n540), .A2(new_n544), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n562), .ZN(new_n567));
  AND2_X1   g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n543), .A2(new_n567), .B1(KEYINPUT41), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n521), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT95), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT95), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n573), .B(new_n521), .C1(new_n566), .C2(new_n570), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OR3_X1    g374(.A1(new_n566), .A2(new_n570), .A3(new_n521), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n568), .A2(KEYINPUT41), .ZN(new_n577));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n575), .B(new_n576), .C1(KEYINPUT94), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n572), .A2(new_n576), .A3(new_n574), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n572), .A2(KEYINPUT94), .A3(new_n574), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n579), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(G57gat), .A2(G64gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(G57gat), .A2(G64gat), .ZN(new_n587));
  INV_X1    g386(.A(G71gat), .ZN(new_n588));
  INV_X1    g387(.A(G78gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n586), .B(new_n587), .C1(new_n590), .C2(KEYINPUT9), .ZN(new_n591));
  XOR2_X1   g390(.A(G71gat), .B(G78gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G127gat), .B(G155gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT89), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT16), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(G1gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G15gat), .B(G22gat), .ZN(new_n607));
  MUX2_X1   g406(.A(G1gat), .B(new_n606), .S(new_n607), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G8gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n593), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(KEYINPUT21), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n602), .A2(new_n614), .A3(new_n603), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n613), .B2(new_n615), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n609), .A2(new_n562), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n564), .A2(new_n565), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n609), .ZN(new_n622));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(KEYINPUT18), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(KEYINPUT13), .Z(new_n625));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n567), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(new_n626), .B2(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT18), .B1(new_n622), .B2(new_n623), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(new_n227), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n382), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n628), .A2(new_n629), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n634), .B1(new_n628), .B2(new_n629), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT88), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(KEYINPUT88), .B(new_n634), .C1(new_n628), .C2(new_n629), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT96), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n611), .B1(new_n536), .B2(new_n537), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n541), .A2(new_n593), .A3(new_n542), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT97), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n543), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n643), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n647), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n642), .B1(new_n649), .B2(new_n650), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n655), .B1(new_n658), .B2(new_n646), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n640), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n585), .A2(new_n619), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n520), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT98), .ZN(new_n664));
  INV_X1    g463(.A(new_n376), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(new_n664), .ZN(new_n668));
  OAI21_X1  g467(.A(G8gat), .B1(new_n668), .B2(new_n413), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  INV_X1    g469(.A(new_n413), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n664), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n673), .A2(KEYINPUT99), .A3(new_n670), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT99), .B1(new_n673), .B2(new_n670), .ZN(new_n675));
  OAI221_X1 g474(.A(new_n669), .B1(new_n670), .B2(new_n673), .C1(new_n674), .C2(new_n675), .ZN(G1325gat));
  INV_X1    g475(.A(new_n316), .ZN(new_n677));
  OAI21_X1  g476(.A(G15gat), .B1(new_n668), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n679), .A3(new_n505), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n456), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  AOI21_X1  g483(.A(new_n585), .B1(new_n504), .B2(new_n519), .ZN(new_n685));
  INV_X1    g484(.A(new_n619), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n661), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n550), .A3(new_n665), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n455), .A2(new_n505), .A3(new_n517), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n692), .B1(new_n488), .B2(new_n487), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT35), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n671), .B1(new_n373), .B2(new_n375), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n516), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT102), .B1(new_n507), .B2(new_n518), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n504), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n457), .B(KEYINPUT101), .C1(new_n486), .C2(new_n503), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n581), .A2(new_n584), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT100), .B1(new_n685), .B2(new_n705), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n709), .B(KEYINPUT44), .C1(new_n520), .C2(new_n585), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n711), .A2(new_n665), .A3(new_n688), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n691), .B1(new_n712), .B2(new_n550), .ZN(G1328gat));
  INV_X1    g512(.A(new_n689), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G36gat), .A3(new_n413), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT103), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n711), .A2(new_n671), .A3(new_n688), .ZN(new_n719));
  OAI221_X1 g518(.A(new_n718), .B1(new_n716), .B2(new_n715), .C1(new_n551), .C2(new_n719), .ZN(G1329gat));
  NAND3_X1  g519(.A1(new_n711), .A2(new_n316), .A3(new_n688), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G43gat), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n714), .A2(G43gat), .A3(new_n315), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n721), .B2(G43gat), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n729), .A2(new_n731), .A3(new_n723), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n728), .B1(KEYINPUT47), .B2(new_n732), .ZN(G1330gat));
  NAND4_X1  g532(.A1(new_n711), .A2(G50gat), .A3(new_n456), .A4(new_n688), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n546), .B1(new_n714), .B2(new_n455), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g536(.A(new_n640), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n686), .A2(new_n706), .A3(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n660), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n704), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n665), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT106), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n747), .A2(new_n413), .A3(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n749), .A2(KEYINPUT49), .A3(G64gat), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT49), .B(G64gat), .Z(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(G1333gat));
  NAND3_X1  g551(.A1(new_n743), .A2(new_n588), .A3(new_n505), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n747), .A2(new_n677), .A3(new_n748), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n588), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1334gat));
  NOR3_X1   g556(.A1(new_n747), .A2(new_n455), .A3(new_n748), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(new_n589), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n619), .A2(new_n738), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n704), .A2(new_n706), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n706), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(new_n522), .A3(new_n665), .A4(new_n660), .ZN(new_n766));
  INV_X1    g565(.A(new_n660), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n619), .A2(new_n738), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n711), .A2(KEYINPUT108), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT108), .B1(new_n711), .B2(new_n768), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n769), .A2(new_n770), .A3(new_n376), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n766), .B1(new_n771), .B2(new_n522), .ZN(G1336gat));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n763), .A2(new_n773), .A3(new_n764), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n767), .A2(G92gat), .A3(new_n413), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n761), .A2(KEYINPUT109), .A3(new_n762), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n769), .A2(new_n770), .A3(new_n413), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(G92gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n711), .A2(new_n768), .ZN(new_n781));
  OAI21_X1  g580(.A(G92gat), .B1(new_n781), .B2(new_n413), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n765), .B2(new_n775), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n782), .B2(new_n785), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n779), .A2(new_n780), .B1(new_n786), .B2(new_n787), .ZN(G1337gat));
  XNOR2_X1  g587(.A(KEYINPUT112), .B(G99gat), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n765), .A2(new_n505), .A3(new_n660), .A4(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n769), .A2(new_n770), .A3(new_n677), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(new_n789), .ZN(G1338gat));
  NOR3_X1   g591(.A1(new_n767), .A2(G106gat), .A3(new_n455), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n774), .A2(KEYINPUT113), .A3(new_n776), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n774), .A2(new_n776), .A3(new_n793), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n769), .A2(new_n770), .A3(new_n455), .ZN(new_n798));
  INV_X1    g597(.A(G106gat), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n794), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT53), .ZN(new_n801));
  OAI21_X1  g600(.A(G106gat), .B1(new_n781), .B2(new_n455), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT53), .B1(new_n765), .B2(new_n793), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n656), .B1(new_n658), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n652), .A2(KEYINPUT54), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n651), .A2(new_n643), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT55), .B(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n657), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n810), .A2(new_n657), .A3(KEYINPUT114), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n738), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n635), .ZN(new_n818));
  INV_X1    g617(.A(new_n633), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n622), .A2(new_n623), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n626), .A2(new_n620), .A3(new_n625), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n660), .A3(KEYINPUT115), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n818), .A2(new_n822), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n767), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n706), .B1(new_n817), .B2(new_n828), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n706), .A2(new_n816), .A3(new_n815), .A4(new_n823), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n686), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n686), .A2(new_n706), .A3(new_n738), .A4(new_n660), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n376), .A2(new_n671), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n506), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n738), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n660), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n619), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G127gat), .ZN(G1342gat));
  AOI21_X1  g642(.A(new_n585), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n834), .A2(new_n516), .A3(new_n835), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n845), .B(new_n846), .Z(G1343gat));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n316), .A2(new_n455), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n640), .A2(G141gat), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n836), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n677), .A2(new_n835), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n814), .A2(new_n813), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n657), .A3(new_n810), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n857), .A2(new_n640), .B1(new_n767), .B2(new_n826), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n585), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n706), .A2(new_n815), .A3(new_n816), .A4(new_n823), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n619), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n456), .B1(new_n861), .B2(new_n832), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n855), .B1(new_n862), .B2(KEYINPUT57), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n834), .A2(new_n864), .A3(new_n456), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n865), .A3(new_n738), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n853), .B1(G141gat), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT117), .B1(new_n866), .B2(G141gat), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  AOI221_X4 g669(.A(new_n853), .B1(KEYINPUT117), .B2(new_n870), .C1(G141gat), .C2(new_n866), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n848), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n873));
  INV_X1    g672(.A(new_n867), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n867), .B1(new_n868), .B2(KEYINPUT58), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(KEYINPUT118), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n872), .A2(new_n877), .ZN(G1344gat));
  OR2_X1    g677(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n455), .B1(new_n831), .B2(new_n833), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n879), .B(new_n660), .C1(new_n864), .C2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT59), .B(G148gat), .C1(new_n881), .C2(new_n855), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n836), .A2(new_n850), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n660), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n863), .A2(new_n865), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n660), .A2(new_n883), .ZN(new_n887));
  OAI221_X1 g686(.A(new_n882), .B1(G148gat), .B2(new_n885), .C1(new_n886), .C2(new_n887), .ZN(G1345gat));
  OAI21_X1  g687(.A(G155gat), .B1(new_n886), .B2(new_n686), .ZN(new_n889));
  INV_X1    g688(.A(G155gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n890), .A3(new_n619), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n886), .B2(new_n585), .ZN(new_n893));
  INV_X1    g692(.A(G162gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n884), .A2(new_n894), .A3(new_n706), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n665), .A2(new_n413), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n834), .A2(new_n516), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT119), .Z(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n227), .A3(new_n738), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n901));
  INV_X1    g700(.A(new_n897), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n831), .B2(new_n833), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n903), .A2(KEYINPUT121), .A3(new_n516), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT121), .B1(new_n903), .B2(new_n516), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n640), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n901), .A2(new_n907), .A3(new_n908), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n899), .B2(new_n660), .ZN(new_n910));
  OAI211_X1 g709(.A(G176gat), .B(new_n660), .C1(new_n904), .C2(new_n905), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT122), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n906), .B2(new_n686), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n903), .A2(new_n266), .A3(new_n516), .A4(new_n619), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g716(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(G1350gat));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n898), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n903), .A2(KEYINPUT121), .A3(new_n516), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n585), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT61), .B1(new_n923), .B2(new_n241), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n706), .B1(new_n904), .B2(new_n905), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(G190gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n931), .B(KEYINPUT61), .C1(new_n923), .C2(new_n241), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n926), .A2(KEYINPUT125), .A3(new_n927), .A4(G190gat), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n925), .A2(new_n930), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n899), .A2(new_n241), .A3(new_n706), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1351gat));
  AND2_X1   g735(.A1(new_n903), .A2(new_n849), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n382), .B1(new_n938), .B2(new_n640), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n902), .A2(new_n316), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n879), .B(new_n940), .C1(new_n880), .C2(new_n864), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n738), .A2(G197gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(G1352gat));
  NAND3_X1  g743(.A1(new_n937), .A2(new_n380), .A3(new_n660), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n940), .ZN(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n881), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(G1353gat));
  OAI21_X1  g751(.A(G211gat), .B1(new_n941), .B2(new_n686), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n686), .A2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n938), .B2(new_n956), .ZN(G1354gat));
  AOI21_X1  g756(.A(G218gat), .B1(new_n937), .B2(new_n706), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT127), .Z(new_n959));
  INV_X1    g758(.A(G218gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n941), .A2(new_n960), .A3(new_n585), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n959), .A2(new_n961), .ZN(G1355gat));
endmodule


