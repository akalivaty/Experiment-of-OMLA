//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G221), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n187), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(G125), .A2(G140), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT78), .B(G125), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G140), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n194), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  OR3_X1    g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  XOR2_X1   g015(.A(G125), .B(G140), .Z(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT70), .B(G128), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT24), .B(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n210), .A2(KEYINPUT23), .A3(G128), .ZN(new_n216));
  INV_X1    g030(.A(new_n211), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n215), .B1(G110), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n205), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n200), .B1(new_n197), .B2(new_n199), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n201), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n211), .A2(new_n212), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n218), .B2(G110), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT80), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n205), .A2(new_n219), .B1(new_n224), .B2(new_n222), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT80), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n192), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n191), .B1(new_n228), .B2(new_n229), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(KEYINPUT81), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT77), .B(G902), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n237), .B2(G234), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(G902), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT25), .B1(new_n233), .B2(new_n237), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n242));
  NOR4_X1   g056(.A1(new_n231), .A2(new_n242), .A3(new_n236), .A4(new_n232), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n238), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT66), .B(G137), .Z(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT11), .A3(G134), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT11), .B1(new_n248), .B2(G134), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(G134), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT67), .B(G131), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n246), .B2(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n200), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT69), .B(KEYINPUT1), .C1(new_n259), .C2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n206), .A2(KEYINPUT70), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G128), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT69), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n261), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(KEYINPUT71), .B(new_n261), .C1(new_n266), .C2(new_n267), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT65), .B1(new_n200), .B2(G143), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n259), .A3(G146), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n272), .A2(new_n274), .B1(G143), .B2(new_n200), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n206), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n270), .A2(new_n271), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT73), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n268), .A2(new_n269), .B1(new_n275), .B2(new_n276), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n271), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n257), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT66), .B(G137), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n285));
  INV_X1    g099(.A(G134), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n251), .ZN(new_n288));
  OAI21_X1  g102(.A(G131), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n289), .A2(new_n253), .ZN(new_n290));
  NAND2_X1  g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n275), .A2(new_n292), .B1(new_n294), .B2(new_n261), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT30), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n210), .A2(G116), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G119), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT2), .B(G113), .Z(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n304), .A2(new_n305), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n297), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n257), .B(KEYINPUT68), .ZN(new_n312));
  INV_X1    g126(.A(new_n278), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n299), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n310), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n298), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(G237), .A2(G953), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G210), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n317), .A2(new_n319), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT31), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n298), .A2(KEYINPUT28), .A3(new_n318), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n314), .A2(new_n310), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n325), .B(KEYINPUT74), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT31), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n317), .A2(new_n336), .A3(new_n319), .A4(new_n326), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n328), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(G472), .A2(G902), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n338), .A2(KEYINPUT32), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT32), .B1(new_n338), .B2(new_n339), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n317), .A2(new_n319), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT29), .B1(new_n343), .B2(new_n325), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n345));
  INV_X1    g159(.A(new_n334), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n330), .A2(new_n331), .A3(new_n332), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n310), .B1(new_n283), .B2(new_n297), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n329), .B1(new_n319), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT28), .B1(new_n298), .B2(new_n318), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT76), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n352), .A2(KEYINPUT29), .A3(new_n326), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n237), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n345), .B1(new_n344), .B2(new_n347), .ZN(new_n356));
  OAI21_X1  g170(.A(G472), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n245), .B1(new_n342), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G902), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT94), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G143), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n259), .A2(KEYINPUT94), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G214), .A4(new_n320), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n320), .A2(G214), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(new_n362), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n366), .A2(new_n252), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n252), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n366), .A2(new_n368), .A3(new_n252), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(new_n201), .A3(new_n221), .A4(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n203), .B1(G146), .B2(new_n195), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n366), .B(new_n376), .Z(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n374), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G113), .B(G122), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n372), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n372), .B2(new_n379), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n360), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G475), .ZN(new_n387));
  NOR2_X1   g201(.A1(G475), .A2(G902), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n202), .A2(KEYINPUT19), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(KEYINPUT19), .B2(new_n195), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n200), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n367), .A2(new_n369), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n201), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n379), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n382), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n389), .B1(new_n397), .B2(new_n383), .ZN(new_n398));
  XOR2_X1   g212(.A(KEYINPUT93), .B(KEYINPUT20), .Z(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI211_X1 g215(.A(KEYINPUT20), .B(new_n389), .C1(new_n397), .C2(new_n383), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n387), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G952), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G953), .ZN(new_n405));
  INV_X1    g219(.A(G237), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n189), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G953), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n409), .B(new_n237), .C1(G234), .C2(G237), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT21), .B(G898), .Z(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n403), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n259), .A2(G128), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n209), .A2(new_n259), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT13), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT97), .ZN(new_n419));
  OAI22_X1  g233(.A1(new_n418), .A2(new_n419), .B1(new_n417), .B2(new_n415), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  OAI21_X1  g235(.A(G134), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n416), .B1(G128), .B2(new_n259), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n286), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n301), .A2(G122), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT96), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n301), .A2(G122), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G107), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n422), .A2(new_n424), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n428), .B2(KEYINPUT14), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n429), .B(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n423), .B(new_n286), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT9), .B(G234), .Z(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(G217), .A3(new_n409), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n432), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n432), .B2(new_n436), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n237), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n432), .A2(new_n436), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n438), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n236), .B1(new_n448), .B2(new_n440), .ZN(new_n449));
  INV_X1    g263(.A(new_n445), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n446), .A2(new_n451), .A3(KEYINPUT98), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT98), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n443), .A2(new_n445), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n449), .A2(new_n450), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n414), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OR3_X1    g272(.A1(new_n381), .A2(KEYINPUT3), .A3(G107), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n381), .A2(G107), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n459), .B(new_n322), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT4), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n459), .B1(new_n461), .B2(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G101), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n463), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n310), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT5), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n210), .A3(G116), .ZN(new_n469));
  OAI211_X1 g283(.A(G113), .B(new_n469), .C1(new_n303), .C2(new_n468), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n306), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n470), .A2(new_n471), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n430), .A2(G104), .ZN(new_n476));
  OAI21_X1  g290(.A(G101), .B1(new_n460), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n462), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G122), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT88), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n467), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n462), .A2(new_n477), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n481), .B(KEYINPUT8), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n306), .A2(new_n470), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n484), .B(new_n485), .C1(new_n483), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G224), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(G953), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n493), .A2(KEYINPUT7), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n296), .A2(KEYINPUT89), .A3(new_n194), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n295), .B2(new_n198), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n313), .A2(new_n198), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n494), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n490), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(KEYINPUT90), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n504), .A3(new_n497), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n503), .A2(new_n505), .A3(new_n500), .A4(new_n494), .ZN(new_n506));
  AOI21_X1  g320(.A(G902), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n505), .A3(new_n500), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n492), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n503), .A2(new_n493), .A3(new_n500), .A4(new_n505), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n467), .A2(new_n479), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n513));
  INV_X1    g327(.A(new_n481), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n514), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n482), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G210), .B1(G237), .B2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n507), .A2(new_n520), .A3(new_n518), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(KEYINPUT92), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G214), .B1(G237), .B2(G902), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n523), .A2(KEYINPUT92), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n458), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n270), .A2(new_n271), .A3(new_n277), .A4(new_n483), .ZN(new_n529));
  INV_X1    g343(.A(new_n277), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n275), .A2(new_n276), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n478), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n290), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT84), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(KEYINPUT85), .A3(new_n536), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n290), .B1(new_n529), .B2(new_n532), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT84), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT12), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT85), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n539), .B2(KEYINPUT12), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n537), .A2(new_n538), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n478), .A2(KEYINPUT10), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AND4_X1   g360(.A1(new_n281), .A2(new_n270), .A3(new_n271), .A4(new_n277), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n281), .B1(new_n280), .B2(new_n271), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT83), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n553));
  AOI22_X1  g367(.A1(new_n466), .A2(new_n295), .B1(new_n532), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n551), .A2(new_n290), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G110), .B(G140), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n409), .A2(G227), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n556), .B(new_n557), .Z(new_n558));
  AND3_X1   g372(.A1(new_n544), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n545), .B1(new_n279), .B2(new_n282), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n554), .B1(new_n560), .B2(KEYINPUT83), .ZN(new_n561));
  INV_X1    g375(.A(new_n552), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n534), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n558), .B1(new_n563), .B2(new_n555), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G469), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n237), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT86), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n563), .A2(new_n555), .A3(new_n558), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n558), .B1(new_n544), .B2(new_n555), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n544), .A2(new_n555), .ZN(new_n572));
  INV_X1    g386(.A(new_n558), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n563), .A2(new_n555), .A3(new_n558), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(KEYINPUT86), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n571), .A2(G469), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n566), .A2(new_n360), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n567), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n188), .B1(new_n437), .B2(new_n360), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n528), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n359), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(new_n322), .ZN(G3));
  INV_X1    g400(.A(new_n245), .ZN(new_n587));
  INV_X1    g401(.A(G472), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n338), .B2(new_n237), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n338), .B2(new_n339), .ZN(new_n590));
  INV_X1    g404(.A(new_n525), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n522), .B2(new_n523), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n583), .A2(new_n587), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n443), .A2(G478), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n441), .B2(new_n442), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n448), .A2(KEYINPUT33), .A3(new_n440), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n237), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n598), .B2(G478), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n403), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n593), .A2(new_n413), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT34), .B(G104), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  INV_X1    g417(.A(new_n387), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n456), .B2(new_n452), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n413), .B(KEYINPUT99), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n398), .A2(new_n400), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n398), .A2(new_n400), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT100), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n605), .A2(KEYINPUT100), .A3(new_n609), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n593), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT35), .B(G107), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G9));
  NOR2_X1   g428(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n226), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n239), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n244), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n528), .A2(new_n583), .A3(new_n590), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G110), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n619), .B(new_n621), .ZN(G12));
  AND2_X1   g436(.A1(new_n244), .A2(new_n617), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n342), .B2(new_n357), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n580), .A2(new_n582), .A3(new_n592), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n607), .A2(new_n608), .ZN(new_n626));
  INV_X1    g440(.A(G900), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n408), .B1(new_n410), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n604), .B(new_n630), .C1(new_n452), .C2(new_n456), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n624), .A2(new_n625), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  AND2_X1   g447(.A1(new_n319), .A2(new_n349), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n327), .B1(new_n634), .B2(new_n346), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n360), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n342), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n524), .A2(new_n526), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT103), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n640), .B(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n403), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n456), .B2(new_n452), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n623), .A2(new_n525), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n639), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n628), .B(KEYINPUT39), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n583), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(KEYINPUT40), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(KEYINPUT40), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G143), .ZN(G45));
  NAND2_X1  g467(.A1(new_n598), .A2(G478), .ZN(new_n654));
  INV_X1    g468(.A(new_n594), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n654), .A2(new_n655), .A3(new_n403), .A4(new_n629), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n599), .A2(KEYINPUT104), .A3(new_n403), .A4(new_n629), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n624), .A2(new_n625), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G146), .ZN(G48));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n237), .B1(new_n559), .B2(new_n564), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G469), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n567), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(KEYINPUT105), .A3(G469), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n669), .A2(new_n582), .A3(new_n592), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n600), .A2(new_n413), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n358), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NOR2_X1   g488(.A1(new_n611), .A2(new_n610), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n670), .A2(new_n358), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  NAND3_X1  g491(.A1(new_n670), .A2(new_n624), .A3(new_n457), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G119), .ZN(G21));
  NAND2_X1  g493(.A1(new_n645), .A2(new_n592), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n645), .A2(KEYINPUT107), .A3(new_n592), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n606), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n339), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n352), .A2(new_n353), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT106), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n352), .A2(new_n688), .A3(new_n353), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n687), .A2(new_n334), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n328), .A2(new_n337), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n685), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n589), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n581), .B1(new_n667), .B2(new_n668), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n684), .A2(new_n693), .A3(new_n587), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT108), .B(G122), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G24));
  NAND3_X1  g511(.A1(new_n693), .A2(new_n618), .A3(new_n661), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n592), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT109), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n692), .A2(new_n623), .A3(new_n660), .A4(new_n589), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n702), .A3(new_n670), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n340), .B2(new_n341), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n338), .A2(new_n339), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT32), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n338), .A2(KEYINPUT32), .A3(new_n339), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(KEYINPUT110), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n712), .A3(new_n357), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n574), .A2(new_n575), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n567), .B(new_n579), .C1(new_n566), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n591), .B1(new_n524), .B2(new_n526), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n715), .A2(new_n716), .A3(new_n582), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n713), .A2(new_n587), .A3(new_n661), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n342), .A2(new_n357), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n717), .A2(new_n719), .A3(new_n587), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n660), .A2(KEYINPUT42), .ZN(new_n721));
  AOI22_X1  g535(.A1(KEYINPUT42), .A2(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  NAND3_X1  g537(.A1(new_n358), .A2(new_n631), .A3(new_n717), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n714), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n726), .A2(new_n566), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n566), .B1(new_n714), .B2(new_n568), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n729), .B1(new_n730), .B2(new_n576), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n728), .B1(new_n731), .B2(KEYINPUT111), .ZN(new_n732));
  INV_X1    g546(.A(new_n729), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n577), .A2(KEYINPUT111), .A3(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(KEYINPUT46), .B(new_n579), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT111), .B1(new_n577), .B2(new_n733), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n734), .A2(new_n739), .A3(new_n727), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n738), .B1(new_n740), .B2(new_n578), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n731), .A2(KEYINPUT111), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n577), .A2(new_n733), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n745), .A3(new_n728), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(KEYINPUT112), .A3(KEYINPUT46), .A4(new_n579), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n737), .A2(new_n567), .A3(new_n741), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n582), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT43), .B1(new_n644), .B2(KEYINPUT113), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n599), .A2(new_n644), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT114), .ZN(new_n754));
  INV_X1    g568(.A(new_n590), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n618), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n716), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n750), .A2(new_n758), .A3(new_n648), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  NAND2_X1  g576(.A1(new_n749), .A2(KEYINPUT47), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n748), .A2(new_n764), .A3(new_n582), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n719), .A2(new_n587), .A3(new_n660), .A4(new_n759), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NAND2_X1  g582(.A1(new_n404), .A2(new_n409), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n624), .B(new_n625), .C1(new_n631), .C2(new_n661), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n618), .B(new_n628), .C1(new_n682), .C2(new_n683), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n582), .A3(new_n638), .A4(new_n715), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n698), .A2(KEYINPUT109), .A3(new_n699), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n702), .B1(new_n701), .B2(new_n670), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n770), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n704), .A2(KEYINPUT52), .A3(new_n770), .A4(new_n772), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n692), .A2(new_n623), .A3(new_n589), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n661), .A3(new_n717), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n446), .A2(new_n451), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n630), .A2(new_n782), .A3(new_n604), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n716), .A2(new_n618), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n719), .A2(new_n784), .A3(new_n583), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n724), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n644), .A2(new_n782), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n600), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n527), .A3(new_n606), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n583), .A3(new_n587), .A4(new_n590), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n792), .B(new_n619), .C1(new_n359), .C2(new_n584), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n787), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n678), .A2(new_n676), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n672), .A2(new_n695), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n722), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n779), .A2(new_n796), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n795), .B(new_n799), .C1(new_n777), .C2(new_n778), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n803), .B(KEYINPUT54), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n799), .B1(new_n777), .B2(new_n778), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n787), .A2(new_n794), .A3(KEYINPUT116), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n786), .B2(new_n793), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n808), .A2(KEYINPUT53), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n812), .B(new_n813), .C1(new_n804), .C2(new_n801), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n806), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n245), .A2(new_n407), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n639), .A2(new_n694), .A3(new_n716), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n600), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n405), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n753), .A2(new_n408), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n821), .A2(new_n245), .A3(new_n589), .A4(new_n692), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n820), .B1(new_n670), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n713), .A2(new_n587), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n669), .A2(new_n582), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n821), .A2(new_n825), .A3(new_n759), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT48), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n823), .A2(KEYINPUT118), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT118), .B1(new_n823), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n643), .A2(new_n591), .A3(new_n694), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n822), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n822), .A2(KEYINPUT50), .A3(new_n832), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n669), .A2(new_n581), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n763), .B2(new_n765), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n822), .A2(new_n716), .ZN(new_n841));
  OAI211_X1 g655(.A(KEYINPUT117), .B(new_n837), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n599), .A2(new_n403), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n817), .A2(new_n843), .B1(new_n780), .B2(new_n826), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n837), .B(new_n844), .C1(new_n840), .C2(new_n841), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n845), .A3(KEYINPUT51), .ZN(new_n846));
  INV_X1    g660(.A(new_n837), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n748), .A2(new_n764), .A3(new_n582), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n764), .B1(new_n748), .B2(new_n582), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n838), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n841), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n852), .B(new_n844), .C1(KEYINPUT117), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n831), .B1(new_n846), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n815), .B1(new_n855), .B2(KEYINPUT119), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n857), .B(new_n831), .C1(new_n846), .C2(new_n854), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n769), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n669), .B(KEYINPUT49), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n245), .A2(new_n581), .A3(new_n591), .A4(new_n752), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n639), .A3(new_n643), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(G75));
  NAND2_X1  g677(.A1(new_n807), .A2(new_n796), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n802), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n237), .B1(new_n865), .B2(new_n812), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n521), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n517), .A2(new_n515), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n511), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n867), .B2(new_n868), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n409), .A2(G952), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G51));
  INV_X1    g689(.A(new_n812), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n801), .B1(new_n807), .B2(new_n796), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n878), .A2(KEYINPUT121), .A3(new_n237), .A4(new_n746), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n866), .B2(new_n740), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT54), .B1(new_n876), .B2(new_n877), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n814), .ZN(new_n884));
  XNOR2_X1  g698(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n578), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n565), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n874), .B1(new_n882), .B2(new_n888), .ZN(G54));
  AND2_X1   g703(.A1(KEYINPUT58), .A2(G475), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n236), .B(new_n890), .C1(new_n876), .C2(new_n877), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n397), .A3(new_n383), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n397), .A2(new_n383), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n866), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  INV_X1    g708(.A(new_n874), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT122), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(G60));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT59), .Z(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n806), .B2(new_n814), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n596), .A2(new_n597), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n895), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n906));
  INV_X1    g720(.A(new_n904), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n902), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n884), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n908), .ZN(new_n910));
  AOI211_X1 g724(.A(KEYINPUT123), .B(new_n910), .C1(new_n883), .C2(new_n814), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n905), .A2(new_n909), .A3(new_n911), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n616), .B(new_n915), .C1(new_n876), .C2(new_n877), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(new_n895), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  INV_X1    g733(.A(new_n234), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n878), .B2(new_n914), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n917), .A2(new_n918), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n918), .A2(new_n919), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n916), .A2(new_n895), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n865), .A2(new_n812), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n234), .B1(new_n926), .B2(new_n915), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n922), .A2(new_n928), .ZN(G66));
  OAI21_X1  g743(.A(G953), .B1(new_n412), .B2(new_n491), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n797), .A2(new_n798), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n793), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n932), .B2(G953), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n869), .B1(G898), .B2(new_n409), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  INV_X1    g749(.A(new_n770), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n700), .B2(new_n703), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n761), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n761), .A2(KEYINPUT126), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n682), .A2(new_n683), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n750), .A2(new_n648), .A3(new_n942), .A4(new_n824), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n722), .A2(new_n724), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n940), .A2(new_n767), .A3(new_n941), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n409), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n299), .A2(new_n316), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(new_n391), .Z(new_n949));
  OAI211_X1 g763(.A(new_n947), .B(new_n949), .C1(G227), .C2(new_n409), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n949), .A2(G227), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n409), .B1(new_n951), .B2(G900), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n789), .A2(KEYINPUT125), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n716), .B1(KEYINPUT125), .B2(new_n789), .ZN(new_n954));
  OR4_X1    g768(.A1(new_n359), .A2(new_n649), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n761), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n937), .A2(new_n652), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n937), .A2(KEYINPUT62), .A3(new_n652), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n956), .A2(new_n767), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n949), .A2(G953), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n952), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n950), .A2(new_n964), .ZN(G72));
  NAND4_X1  g779(.A1(new_n956), .A2(new_n961), .A3(new_n767), .A4(new_n932), .ZN(new_n966));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT63), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n326), .A3(new_n343), .ZN(new_n970));
  INV_X1    g784(.A(new_n968), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n343), .A2(new_n325), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n327), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n803), .B(new_n973), .C1(new_n804), .C2(new_n805), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n895), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n343), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n325), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n945), .A2(new_n767), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n979), .A2(new_n932), .A3(new_n940), .A4(new_n941), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n980), .B2(new_n968), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT127), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n932), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n968), .B1(new_n946), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n325), .A3(new_n977), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n986), .A3(new_n970), .A4(new_n975), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n982), .A2(new_n987), .ZN(G57));
endmodule


