//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT65), .ZN(G160));
  INV_X1    g048(.A(new_n469), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n462), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(G162));
  AND2_X1   g055(.A1(G126), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n462), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT66), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n462), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n464), .A2(G138), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n462), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n464), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n488), .A2(KEYINPUT67), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT67), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n462), .A2(KEYINPUT68), .A3(new_n487), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n462), .A2(KEYINPUT68), .A3(new_n487), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(new_n493), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n486), .A2(new_n492), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  OR2_X1    g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n507), .A2(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n505), .A2(new_n515), .ZN(G166));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n500), .A2(new_n501), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT69), .B(G89), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n525), .B1(new_n517), .B2(new_n518), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n521), .A2(new_n523), .A3(new_n524), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND2_X1  g104(.A1(new_n526), .A2(G52), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n519), .A2(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n502), .A2(G64), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n504), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n530), .B(new_n531), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(KEYINPUT70), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  OAI211_X1 g115(.A(G43), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n513), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n502), .A2(new_n506), .A3(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n546), .A2(KEYINPUT71), .A3(new_n541), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n510), .A2(new_n509), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n545), .A2(new_n547), .B1(G651), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n500), .A2(new_n559), .A3(new_n501), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT73), .B1(new_n510), .B2(new_n509), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT9), .B1(new_n507), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n526), .A2(new_n568), .A3(G53), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n519), .A2(KEYINPUT72), .A3(G91), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n513), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n565), .A2(new_n570), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G166), .ZN(G303));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n507), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n526), .A2(KEYINPUT74), .A3(G49), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n504), .B1(new_n549), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(G87), .B2(new_n519), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(G288));
  AOI22_X1  g162(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n504), .ZN(new_n589));
  INV_X1    g164(.A(G48), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n507), .A2(new_n590), .B1(new_n513), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AND2_X1   g169(.A1(G72), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n502), .B2(G60), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n504), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n519), .A2(G85), .B1(new_n526), .B2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n506), .A2(G54), .A3(G543), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n513), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT10), .A4(G92), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n560), .B2(new_n561), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT75), .Z(new_n611));
  OAI21_X1  g186(.A(G651), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g187(.A1(new_n607), .A2(KEYINPUT76), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(KEYINPUT76), .B1(new_n607), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n600), .B1(new_n615), .B2(G868), .ZN(G284));
  XOR2_X1   g191(.A(G284), .B(KEYINPUT77), .Z(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT78), .Z(new_n619));
  AOI21_X1  g194(.A(G868), .B1(G299), .B2(KEYINPUT79), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(KEYINPUT79), .B2(G299), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(G280));
  XOR2_X1   g197(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n615), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n607), .A2(new_n612), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n607), .A2(KEYINPUT76), .A3(new_n612), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  OR3_X1    g207(.A1(new_n631), .A2(KEYINPUT81), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT81), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G868), .C2(new_n552), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n462), .A2(new_n467), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT82), .B(G2100), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(G111), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(G2105), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n476), .B2(G123), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n474), .A2(new_n646), .A3(G135), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n646), .B1(new_n474), .B2(G135), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n639), .A2(new_n640), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(G2096), .ZN(new_n652));
  NAND4_X1  g227(.A1(new_n641), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(new_n668), .A3(G14), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(KEYINPUT17), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n675), .B2(new_n672), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT85), .Z(new_n677));
  NOR3_X1   g252(.A1(new_n675), .A2(new_n672), .A3(new_n671), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT86), .Z(new_n679));
  NAND3_X1  g254(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT19), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n687), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT20), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(G229));
  NAND3_X1  g280(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT25), .Z(new_n707));
  INV_X1    g282(.A(G139), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n469), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(new_n464), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G29), .ZN(new_n713));
  NOR2_X1   g288(.A1(G29), .A2(G33), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2072), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n474), .A2(G140), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n476), .A2(G128), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n464), .A2(G116), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n718), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G29), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G2067), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n717), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G11), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(G28), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n724), .B1(new_n732), .B2(G28), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n731), .B1(new_n733), .B2(new_n734), .C1(new_n649), .C2(new_n724), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n724), .A2(G32), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT26), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n476), .B2(G129), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n736), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n735), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2078), .ZN(new_n745));
  NAND2_X1  g320(.A1(G164), .A2(G29), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G27), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NOR2_X1   g324(.A1(G171), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G5), .B2(new_n749), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n744), .B1(new_n745), .B2(new_n747), .C1(new_n748), .C2(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n730), .B(new_n752), .C1(new_n745), .C2(new_n747), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(G20), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT23), .Z(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G299), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1956), .ZN(new_n757));
  NAND2_X1  g332(.A1(G168), .A2(G16), .ZN(new_n758));
  NOR2_X1   g333(.A1(G16), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(KEYINPUT95), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(KEYINPUT95), .B2(new_n758), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1966), .ZN(new_n762));
  NOR2_X1   g337(.A1(G29), .A2(G35), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G162), .B2(G29), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G2090), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(G160), .A2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G34), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n770), .B2(KEYINPUT24), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT24), .B2(new_n770), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(G2084), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n766), .A2(new_n767), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n762), .A2(new_n768), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT92), .B(G1341), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n749), .A2(G19), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n552), .B2(new_n749), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT93), .Z(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n753), .A2(new_n757), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n742), .A2(new_n743), .ZN(new_n783));
  AOI21_X1  g358(.A(G2084), .B1(new_n769), .B2(new_n772), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n783), .B(new_n784), .C1(new_n748), .C2(new_n751), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n615), .A2(new_n749), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G4), .B2(new_n749), .ZN(new_n788));
  INV_X1    g363(.A(G1348), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n790), .B(new_n791), .C1(new_n776), .C2(new_n780), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n782), .A2(new_n786), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n724), .A2(G25), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n476), .A2(G119), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT88), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n799));
  INV_X1    g374(.A(G107), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G2105), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n474), .B2(G131), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT89), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G1991), .Z(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n749), .A2(G24), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n596), .A2(new_n504), .ZN(new_n811));
  INV_X1    g386(.A(G47), .ZN(new_n812));
  INV_X1    g387(.A(G85), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n507), .A2(new_n812), .B1(new_n513), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n810), .B1(new_n815), .B2(new_n749), .ZN(new_n816));
  INV_X1    g391(.A(G1986), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n808), .A2(new_n809), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G6), .A2(G16), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n593), .B2(G16), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT32), .B(G1981), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT90), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n749), .A2(G22), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G166), .B2(new_n749), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1971), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n583), .A2(new_n586), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n749), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n749), .B2(G23), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT33), .B(G1976), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n824), .B(new_n832), .C1(new_n830), .C2(new_n831), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT91), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT34), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n819), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n833), .A2(KEYINPUT91), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(KEYINPUT91), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n837), .A2(KEYINPUT34), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n795), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n795), .A3(new_n839), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n794), .B1(new_n841), .B2(new_n842), .ZN(G311));
  INV_X1    g418(.A(new_n842), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n793), .B1(new_n844), .B2(new_n840), .ZN(G150));
  AOI22_X1  g420(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n504), .ZN(new_n847));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n507), .A2(new_n848), .B1(new_n513), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n615), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n551), .A2(G651), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n546), .A2(KEYINPUT71), .A3(new_n541), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT71), .B1(new_n546), .B2(new_n541), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g438(.A(KEYINPUT99), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n851), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n851), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n862), .A3(new_n861), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n857), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT100), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n852), .B1(new_n869), .B2(KEYINPUT39), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n854), .B1(new_n871), .B2(new_n872), .ZN(G145));
  NAND2_X1  g448(.A1(new_n474), .A2(G142), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n476), .A2(G130), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n464), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT102), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n638), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n803), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n712), .B(new_n741), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n722), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n492), .A2(new_n495), .ZN(new_n884));
  INV_X1    g459(.A(new_n485), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n484), .B1(new_n462), .B2(new_n481), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n497), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT101), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n488), .A2(KEYINPUT67), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n489), .A2(new_n491), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n889), .A2(new_n495), .A3(new_n890), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n483), .A2(new_n485), .B1(new_n496), .B2(new_n493), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n883), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n883), .A2(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n881), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n881), .A2(new_n900), .A3(new_n896), .A4(new_n897), .ZN(new_n901));
  INV_X1    g476(.A(new_n881), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n896), .A2(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(G160), .B(new_n649), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(G162), .Z(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT104), .B(G37), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n908), .B1(new_n902), .B2(new_n903), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(new_n898), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  INV_X1    g491(.A(new_n626), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(G299), .ZN(new_n918));
  NAND3_X1  g493(.A1(G299), .A2(new_n612), .A3(new_n607), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n567), .A2(new_n569), .B1(new_n571), .B2(new_n574), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n626), .A2(new_n920), .A3(KEYINPUT105), .A4(new_n565), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n864), .A2(new_n851), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n545), .A2(new_n547), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT99), .B1(new_n924), .B2(new_n858), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n552), .A2(KEYINPUT99), .A3(new_n851), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n926), .A2(new_n630), .A3(new_n927), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n867), .A2(new_n865), .B1(new_n615), .B2(new_n624), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n919), .ZN(new_n931));
  INV_X1    g506(.A(G299), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT105), .B1(new_n932), .B2(new_n626), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT41), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n630), .B1(new_n926), .B2(new_n927), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n865), .A2(new_n615), .A3(new_n624), .A4(new_n867), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n918), .A2(new_n937), .A3(new_n919), .A4(new_n921), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n930), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n934), .A2(new_n938), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n928), .A2(new_n929), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT106), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT109), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n949));
  NOR2_X1   g524(.A1(G288), .A2(G290), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n583), .A2(new_n586), .B1(new_n597), .B2(new_n598), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(G166), .A2(new_n593), .ZN(new_n953));
  OAI22_X1  g528(.A1(new_n505), .A2(new_n515), .B1(new_n589), .B2(new_n592), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G288), .A2(G290), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n815), .A2(new_n583), .A3(new_n586), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT107), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n952), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n955), .A2(KEYINPUT107), .A3(new_n957), .A4(new_n958), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT42), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT108), .B1(new_n960), .B2(new_n961), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(KEYINPUT108), .A3(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n947), .A2(new_n948), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT109), .B1(new_n941), .B2(new_n944), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n960), .A2(KEYINPUT108), .A3(new_n961), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(new_n964), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n962), .B1(new_n973), .B2(KEYINPUT42), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n632), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT110), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n866), .A2(new_n632), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n970), .A2(new_n979), .A3(new_n975), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(G295));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n978), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n979), .B1(new_n970), .B2(new_n975), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n977), .A2(KEYINPUT111), .A3(new_n978), .A4(new_n980), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(G331));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  OAI21_X1  g563(.A(G286), .B1(new_n536), .B2(new_n539), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n538), .A2(KEYINPUT70), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n534), .A2(new_n535), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n531), .A2(new_n530), .ZN(new_n992));
  NAND4_X1  g567(.A1(G168), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n868), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n989), .A2(new_n993), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(new_n867), .A3(new_n865), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n997), .A3(new_n922), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n996), .B1(new_n867), .B2(new_n865), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n868), .A2(new_n994), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n934), .A2(new_n938), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT112), .B1(new_n1003), .B2(new_n967), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n942), .B1(new_n1000), .B2(new_n999), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n973), .A3(new_n1006), .A4(new_n998), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n911), .B1(new_n1003), .B2(new_n967), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n1012));
  AOI21_X1  g587(.A(G37), .B1(new_n1003), .B2(new_n967), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n988), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1008), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1018));
  AND4_X1   g593(.A1(new_n1016), .A2(new_n1017), .A3(KEYINPUT44), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n988), .B1(new_n1010), .B2(KEYINPUT43), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1016), .B1(new_n1020), .B2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1015), .B1(new_n1019), .B2(new_n1021), .ZN(G397));
  XOR2_X1   g597(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n888), .A2(new_n1025), .A3(new_n894), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1024), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G40), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n465), .A2(new_n471), .A3(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n722), .B(new_n728), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n741), .B(G1996), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1030), .B(new_n1032), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT117), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n803), .B(new_n806), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT116), .B1(G290), .B2(G1986), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G290), .A2(G1986), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1384), .B1(new_n891), .B2(new_n892), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1032), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G305), .A2(G1981), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n589), .A2(new_n592), .A3(G1981), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  INV_X1    g627(.A(G1981), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n593), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1054), .B2(new_n1049), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1051), .A2(new_n1055), .A3(G8), .A4(new_n1047), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n828), .ZN(new_n1058));
  OAI211_X1 g633(.A(G8), .B(new_n1047), .C1(new_n1058), .C2(new_n1049), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n828), .A2(G1976), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1047), .A2(G8), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT52), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1047), .A2(new_n1060), .A3(new_n1063), .A4(G8), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1056), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1032), .B1(new_n1046), .B2(new_n1024), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1025), .A2(KEYINPUT45), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n888), .A2(new_n894), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT118), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n888), .A2(new_n894), .A3(new_n1072), .A4(new_n1069), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1068), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n472), .A2(G40), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1025), .B1(new_n884), .B2(new_n887), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(KEYINPUT50), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1046), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1074), .A2(G1971), .B1(G2090), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G303), .A2(G8), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT55), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(G8), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1059), .B1(new_n1067), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT120), .B(new_n1059), .C1(new_n1067), .C2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1078), .B1(new_n498), .B2(new_n1025), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT121), .B1(new_n1091), .B2(new_n1075), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(new_n1032), .C1(new_n1046), .C2(new_n1078), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1079), .A3(new_n1094), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1074), .A2(G1971), .B1(new_n1095), .B2(G2090), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G8), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1083), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1065), .A2(KEYINPUT122), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1056), .A2(new_n1062), .A3(new_n1100), .A4(new_n1064), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1098), .A2(new_n1085), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n498), .A2(new_n1025), .A3(new_n1024), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1104), .B(new_n1032), .C1(new_n1046), .C2(KEYINPUT45), .ZN(new_n1105));
  INV_X1    g680(.A(G1966), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G2084), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1077), .A2(new_n1108), .A3(new_n1079), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(G168), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G8), .ZN(new_n1111));
  AOI21_X1  g686(.A(G168), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT51), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1110), .A2(new_n1115), .A3(G8), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT62), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1074), .A2(new_n745), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1120), .A2(new_n1121), .B1(new_n748), .B2(new_n1080), .ZN(new_n1122));
  OR3_X1    g697(.A1(new_n1105), .A2(KEYINPUT127), .A3(G2078), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT127), .B1(new_n1105), .B2(G2078), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(KEYINPUT53), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1103), .A2(new_n1117), .A3(new_n1119), .A4(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1074), .A2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(G299), .B(KEYINPUT57), .Z(new_n1130));
  INV_X1    g705(.A(G1956), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1095), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1047), .A2(G2067), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1348), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1133), .B(new_n917), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1130), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1128), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1138), .B(new_n1068), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1076), .A2(KEYINPUT50), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1077), .B2(new_n1093), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1956), .B1(new_n1141), .B2(new_n1092), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1137), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1136), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(KEYINPUT61), .A3(new_n1133), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1047), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT58), .B(G1341), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(G1996), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1074), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1146), .B1(new_n1151), .B2(new_n861), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1074), .A2(new_n1150), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT59), .B(new_n552), .C1(new_n1153), .C2(new_n1149), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1145), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1143), .A2(new_n1133), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n626), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1134), .B1(new_n1080), .B2(new_n789), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT126), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n1164));
  NOR4_X1   g739(.A1(new_n1135), .A2(new_n1134), .A3(new_n1164), .A4(new_n1161), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1159), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1134), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1140), .A2(new_n1075), .A3(new_n1091), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1167), .B(new_n1162), .C1(new_n1168), .C2(G1348), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1164), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1159), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1160), .A2(KEYINPUT126), .A3(new_n1162), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1156), .A2(new_n1157), .B1(new_n1166), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1144), .B1(new_n1155), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(G171), .B(KEYINPUT54), .ZN(new_n1176));
  AOI211_X1 g751(.A(G2078), .B(new_n1068), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1177), .A2(KEYINPUT53), .B1(G1961), .B2(new_n1168), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1179), .A2(KEYINPUT53), .A3(new_n745), .A4(new_n1032), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1030), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1176), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1182), .B1(new_n1183), .B2(new_n1176), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1103), .A2(new_n1184), .A3(new_n1118), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1090), .B(new_n1127), .C1(new_n1175), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(G168), .A2(G8), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1098), .A2(new_n1085), .A3(new_n1102), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n1190));
  XNOR2_X1  g765(.A(KEYINPUT123), .B(KEYINPUT63), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1190), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1065), .B(KEYINPUT119), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1194), .A2(KEYINPUT63), .A3(new_n1188), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1081), .A2(G8), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1084), .A2(KEYINPUT125), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1195), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1192), .A2(new_n1193), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1045), .B1(new_n1186), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1038), .A2(new_n1150), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT46), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT46), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1038), .A2(new_n1205), .A3(new_n1150), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT47), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1038), .B1(new_n741), .B2(new_n1034), .ZN(new_n1209));
  AND3_X1   g784(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1208), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1038), .A2(new_n817), .A3(new_n815), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT48), .Z(new_n1213));
  OAI22_X1  g788(.A1(new_n1210), .A2(new_n1211), .B1(new_n1213), .B2(new_n1041), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1037), .A2(new_n806), .A3(new_n798), .A4(new_n802), .ZN(new_n1215));
  OR2_X1    g790(.A1(new_n722), .A2(G2067), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1039), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1202), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g794(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n914), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g796(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1223));
  NOR2_X1   g797(.A1(new_n1222), .A2(new_n1223), .ZN(G308));
  OR2_X1    g798(.A1(new_n1222), .A2(new_n1223), .ZN(G225));
endmodule


