//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT74), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n191), .A2(KEYINPUT74), .A3(G140), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n188), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n187), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n196), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n191), .A2(KEYINPUT74), .A3(G140), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(KEYINPUT74), .ZN(new_n201));
  OAI211_X1 g015(.A(G146), .B(new_n198), .C1(new_n201), .C2(new_n188), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n202), .A3(KEYINPUT75), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n195), .A2(new_n196), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G237), .ZN(new_n208));
  INV_X1    g022(.A(G953), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G214), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n212), .A2(KEYINPUT17), .A3(G131), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT90), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(G131), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n210), .B(G143), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n207), .A2(new_n224), .A3(new_n214), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n216), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G113), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n217), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT18), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n200), .A2(new_n187), .ZN(new_n232));
  INV_X1    g046(.A(new_n201), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n187), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n218), .B1(new_n235), .B2(new_n219), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(new_n229), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n221), .B(KEYINPUT89), .ZN(new_n239));
  XOR2_X1   g053(.A(new_n202), .B(KEYINPUT77), .Z(new_n240));
  MUX2_X1   g054(.A(new_n200), .B(new_n201), .S(KEYINPUT19), .Z(new_n241));
  OR2_X1    g055(.A1(new_n241), .A2(G146), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n237), .ZN(new_n244));
  INV_X1    g058(.A(new_n229), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(G475), .A2(G902), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT20), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT20), .ZN(new_n250));
  INV_X1    g064(.A(new_n248), .ZN(new_n251));
  AOI211_X1 g065(.A(new_n250), .B(new_n251), .C1(new_n238), .C2(new_n246), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n224), .B1(new_n207), .B2(new_n214), .ZN(new_n255));
  AOI211_X1 g069(.A(KEYINPUT90), .B(new_n213), .C1(new_n203), .C2(new_n206), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n255), .A2(new_n256), .A3(new_n222), .ZN(new_n257));
  INV_X1    g071(.A(new_n237), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n257), .A2(new_n245), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n229), .B1(new_n226), .B2(new_n237), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G475), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT92), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT13), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(KEYINPUT92), .A3(KEYINPUT13), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(G143), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n266), .A2(KEYINPUT13), .ZN(new_n273));
  OAI21_X1  g087(.A(G134), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n267), .A2(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G116), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(G122), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT91), .ZN(new_n280));
  INV_X1    g094(.A(G107), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(G122), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n274), .B(new_n277), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n275), .B(new_n276), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n280), .B(new_n282), .C1(KEYINPUT14), .C2(new_n281), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT9), .B(G234), .Z(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G217), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(new_n294), .A3(G953), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n285), .A2(new_n290), .A3(new_n295), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT93), .ZN(new_n299));
  OR3_X1    g113(.A1(new_n291), .A2(KEYINPUT93), .A3(new_n296), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(new_n254), .ZN(new_n301));
  INV_X1    g115(.A(G478), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(KEYINPUT15), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n301), .B(new_n303), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n263), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G952), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G953), .ZN(new_n308));
  NAND2_X1  g122(.A1(G234), .A2(G237), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT21), .B(G898), .Z(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(G902), .A3(G953), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n306), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G210), .B1(G237), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G143), .B(G146), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G128), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n187), .A2(G143), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n211), .A2(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n265), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n323), .B(new_n327), .C1(new_n322), .C2(new_n325), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n191), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT0), .A2(G128), .ZN(new_n330));
  OR2_X1    g144(.A1(KEYINPUT0), .A2(G128), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT64), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n321), .A2(KEYINPUT0), .A3(G128), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n326), .A2(KEYINPUT64), .A3(new_n330), .A4(new_n331), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n329), .B1(new_n337), .B2(new_n191), .ZN(new_n338));
  INV_X1    g152(.A(G224), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G953), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G122), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT85), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT3), .B1(new_n228), .B2(G107), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n281), .A3(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n228), .A2(G107), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G101), .ZN(new_n350));
  INV_X1    g164(.A(G101), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n345), .A2(new_n347), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n354));
  XNOR2_X1  g168(.A(G116), .B(G119), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT2), .B(G113), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n350), .A2(new_n360), .A3(KEYINPUT4), .A4(new_n352), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n354), .A2(new_n358), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n355), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(new_n356), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n278), .A2(KEYINPUT5), .A3(G119), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n355), .B2(KEYINPUT5), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(G113), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n228), .B2(G107), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n281), .A2(KEYINPUT80), .A3(G104), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n348), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G101), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n352), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT81), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n374), .B2(new_n352), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n369), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n344), .B1(new_n364), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n354), .A2(new_n361), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n381), .A2(new_n363), .A3(new_n358), .A4(new_n359), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n362), .A2(KEYINPUT84), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n342), .A3(new_n379), .A4(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT6), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n379), .A3(new_n383), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT6), .B1(new_n387), .B2(new_n343), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n341), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT7), .B1(new_n339), .B2(G953), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n338), .B(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n342), .B(KEYINPUT8), .Z(new_n393));
  INV_X1    g207(.A(new_n375), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT86), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n369), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n384), .B(new_n392), .C1(new_n393), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n254), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n320), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT87), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(new_n320), .C1(new_n390), .C2(new_n398), .ZN(new_n402));
  INV_X1    g216(.A(new_n398), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n387), .A2(new_n343), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n384), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n388), .B1(new_n405), .B2(KEYINPUT6), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n403), .B(new_n319), .C1(new_n406), .C2(new_n341), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT88), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n386), .A2(new_n389), .ZN(new_n409));
  INV_X1    g223(.A(new_n341), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT88), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n403), .A4(new_n319), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n400), .A2(new_n402), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G214), .B1(G237), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n318), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n418));
  INV_X1    g232(.A(G137), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G134), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(G134), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n423), .A2(new_n219), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n276), .A2(G137), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT67), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n421), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n429), .B(G131), .C1(new_n428), .C2(new_n421), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n328), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n422), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(new_n424), .A3(new_n425), .A4(new_n427), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G131), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(new_n426), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n431), .B(new_n357), .C1(new_n435), .C2(new_n337), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT28), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n208), .A2(new_n209), .A3(G210), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT26), .B(G101), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT66), .B1(new_n435), .B2(new_n337), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n434), .A2(new_n426), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n448), .A3(new_n431), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n358), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n437), .A2(new_n443), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n436), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n431), .B(KEYINPUT30), .C1(new_n435), .C2(new_n337), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(new_n449), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n452), .B1(new_n456), .B2(new_n358), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n418), .B(new_n451), .C1(new_n457), .C2(new_n443), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT70), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n457), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n442), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n462), .A2(KEYINPUT70), .A3(new_n418), .A4(new_n451), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n431), .B1(new_n435), .B2(new_n337), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n358), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n437), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT29), .A3(new_n443), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n460), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G472), .ZN(new_n470));
  NOR2_X1   g284(.A1(G472), .A2(G902), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n449), .A2(new_n455), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n358), .A3(new_n453), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT31), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n436), .A4(new_n443), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n437), .A2(new_n450), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n442), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n457), .B2(new_n443), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n471), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT69), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT32), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(KEYINPUT69), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n473), .A2(new_n436), .A3(new_n443), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT31), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n475), .A3(new_n477), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT32), .A3(new_n471), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n470), .A2(new_n482), .A3(new_n484), .A4(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n294), .B1(G234), .B2(new_n254), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n265), .A2(G119), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT72), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT73), .B(KEYINPUT23), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n265), .A2(G119), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n493), .B(new_n495), .C1(new_n499), .C2(new_n494), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n493), .A2(new_n498), .ZN(new_n501));
  XOR2_X1   g315(.A(KEYINPUT24), .B(G110), .Z(new_n502));
  OAI22_X1  g316(.A1(new_n500), .A2(G110), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n240), .A2(new_n503), .A3(new_n232), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(G110), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n203), .A2(new_n505), .A3(new_n206), .A4(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n507), .A2(KEYINPUT76), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(KEYINPUT76), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n209), .A2(G221), .A3(G234), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT22), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(G137), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n504), .B(new_n513), .C1(new_n508), .C2(new_n509), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n254), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT25), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n492), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n515), .A2(new_n516), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n492), .A2(G902), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n491), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G469), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n394), .A2(new_n328), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n394), .A2(new_n328), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n435), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n447), .B(KEYINPUT82), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT10), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n445), .A2(new_n354), .A3(new_n359), .A4(new_n361), .ZN(new_n538));
  OAI211_X1 g352(.A(KEYINPUT10), .B(new_n328), .C1(new_n376), .C2(new_n378), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n535), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n209), .A2(G227), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT78), .ZN(new_n543));
  INV_X1    g357(.A(G110), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n189), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n534), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n538), .A2(new_n539), .A3(new_n537), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT83), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT83), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n538), .A2(new_n539), .A3(new_n551), .A4(new_n537), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n447), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n546), .B1(new_n553), .B2(new_n540), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n529), .B(new_n254), .C1(new_n548), .C2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n529), .A2(new_n254), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n547), .B1(new_n534), .B2(new_n541), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n540), .A3(new_n546), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(G469), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n555), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n417), .A2(new_n528), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(G101), .ZN(G3));
  INV_X1    g380(.A(G472), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n487), .B2(new_n254), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT94), .B1(new_n487), .B2(new_n471), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n572), .A2(new_n525), .A3(new_n563), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n416), .B1(new_n399), .B2(new_n407), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n317), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n299), .A2(new_n300), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT33), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n302), .A2(G902), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n301), .A2(new_n302), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n263), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n573), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT34), .B(G104), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G6));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n229), .B1(new_n243), .B2(new_n237), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n255), .A2(new_n256), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n258), .B1(new_n590), .B2(new_n223), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n591), .B2(new_n229), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n250), .B1(new_n592), .B2(new_n251), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n247), .A2(KEYINPUT20), .A3(new_n248), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G475), .ZN(new_n596));
  INV_X1    g410(.A(new_n260), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n238), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n598), .B2(new_n254), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n305), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n588), .B1(new_n575), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n263), .A2(new_n304), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n603), .A2(KEYINPUT95), .A3(new_n317), .A4(new_n574), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n573), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  INV_X1    g422(.A(new_n572), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n514), .A2(KEYINPUT36), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n510), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n523), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n521), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT96), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n521), .A2(new_n615), .A3(new_n612), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n417), .A2(new_n564), .A3(new_n609), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT97), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT37), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(new_n544), .ZN(G12));
  AND3_X1   g435(.A1(new_n491), .A2(new_n614), .A3(new_n616), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT98), .B(G900), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n311), .B1(new_n315), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n601), .A2(new_n563), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n574), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G128), .ZN(G30));
  NOR2_X1   g441(.A1(new_n414), .A2(KEYINPUT38), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n414), .A2(KEYINPUT38), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n457), .A2(new_n442), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n465), .A2(new_n436), .A3(new_n442), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n254), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n482), .A2(new_n484), .A3(new_n490), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n629), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n624), .B(KEYINPUT39), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT40), .B1(new_n563), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n563), .A2(new_n637), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n600), .A2(new_n304), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NOR4_X1   g457(.A1(new_n636), .A2(new_n643), .A3(new_n416), .A4(new_n617), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n211), .ZN(G45));
  INV_X1    g459(.A(new_n624), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n263), .A2(new_n582), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n622), .A2(new_n564), .A3(new_n574), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  OR2_X1    g464(.A1(new_n548), .A2(new_n554), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n254), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G469), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n562), .A3(new_n555), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n527), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n584), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT41), .B(G113), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT99), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(G15));
  NAND2_X1  g473(.A1(new_n655), .A2(new_n605), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G116), .ZN(G18));
  NOR2_X1   g475(.A1(new_n318), .A2(new_n654), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n622), .A2(new_n574), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  OAI211_X1 g478(.A(new_n486), .B(new_n475), .C1(new_n467), .C2(new_n443), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n568), .B1(new_n471), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n526), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n654), .A2(new_n316), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n642), .A2(KEYINPUT100), .A3(new_n574), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT100), .B1(new_n642), .B2(new_n574), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n667), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  XNOR2_X1  g486(.A(new_n647), .B(KEYINPUT101), .ZN(new_n673));
  INV_X1    g487(.A(new_n654), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(new_n574), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n614), .A2(new_n616), .A3(new_n666), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G125), .ZN(G27));
  NAND2_X1  g492(.A1(new_n400), .A2(new_n402), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n408), .A2(new_n413), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n564), .A3(new_n415), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT102), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n414), .A2(new_n683), .A3(new_n564), .A4(new_n415), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n528), .A3(new_n673), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n480), .A2(new_n483), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n470), .A2(new_n488), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n690), .A2(new_n526), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n685), .A2(KEYINPUT42), .A3(new_n673), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G131), .ZN(G33));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n601), .B2(new_n624), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n603), .A2(KEYINPUT103), .A3(new_n646), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n685), .A2(new_n528), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n685), .A2(new_n701), .A3(new_n528), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G134), .ZN(G36));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n705));
  INV_X1    g519(.A(new_n582), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n595), .B2(new_n599), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n253), .A2(KEYINPUT106), .A3(new_n262), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n262), .A2(new_n593), .A3(new_n594), .A4(new_n582), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n715), .A3(new_n712), .ZN(new_n716));
  AOI22_X1  g530(.A1(KEYINPUT43), .A2(new_n710), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n614), .A2(new_n572), .A3(new_n616), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n705), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n716), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n595), .A2(new_n599), .A3(new_n707), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n253), .B2(new_n262), .ZN(new_n722));
  OAI211_X1 g536(.A(KEYINPUT43), .B(new_n582), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n614), .A2(new_n572), .A3(new_n616), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(KEYINPUT44), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n414), .A2(new_n415), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT45), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n558), .B2(new_n559), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n728), .B(G469), .C1(new_n732), .C2(G902), .ZN(new_n733));
  INV_X1    g547(.A(new_n731), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(G469), .A3(new_n729), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(KEYINPUT46), .A3(new_n557), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n555), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n562), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n637), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n719), .A2(new_n726), .A3(new_n727), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G137), .ZN(G39));
  NAND2_X1  g555(.A1(new_n738), .A2(KEYINPUT47), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n491), .A2(new_n526), .A3(new_n647), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n737), .A2(new_n744), .A3(new_n562), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n743), .A3(new_n727), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G140), .ZN(G42));
  NAND4_X1  g561(.A1(new_n656), .A2(new_n660), .A3(new_n663), .A4(new_n671), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT112), .Z(new_n749));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n688), .A2(new_n692), .B1(new_n700), .B2(new_n702), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n564), .B(new_n635), .C1(new_n669), .C2(new_n670), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n753), .A2(new_n613), .A3(new_n624), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n649), .A2(new_n626), .A3(new_n677), .ZN(new_n755));
  OR3_X1    g569(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT52), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n685), .A2(new_n676), .A3(new_n673), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT109), .B1(new_n306), .B2(new_n646), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n681), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n306), .A2(KEYINPUT109), .A3(new_n646), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n622), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n603), .A2(KEYINPUT108), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n601), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n767), .A3(new_n583), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n414), .A2(new_n416), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n317), .A4(new_n573), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n618), .A2(new_n565), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n764), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n751), .A2(new_n752), .A3(new_n758), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n748), .A2(new_n771), .ZN(new_n774));
  INV_X1    g588(.A(new_n764), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n752), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n756), .A2(new_n757), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n750), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(KEYINPUT54), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n742), .A2(new_n745), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n653), .A2(new_n555), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n562), .B2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n724), .A2(new_n311), .A3(new_n667), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n783), .A2(new_n727), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n727), .A2(new_n674), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT114), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(KEYINPUT114), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n787), .A2(new_n311), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT115), .A3(new_n676), .A4(new_n724), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n787), .A2(new_n311), .A3(new_n724), .A4(new_n788), .ZN(new_n792));
  INV_X1    g606(.A(new_n676), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n785), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n784), .A2(new_n674), .ZN(new_n796));
  INV_X1    g610(.A(new_n630), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n416), .B1(new_n797), .B2(new_n628), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  OAI22_X1  g614(.A1(new_n796), .A2(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n635), .A2(new_n525), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n789), .A2(KEYINPUT116), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n787), .A2(new_n311), .A3(new_n804), .A4(new_n788), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(new_n600), .A3(new_n706), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n795), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n795), .A2(new_n803), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n308), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT48), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n789), .A2(new_n816), .A3(new_n691), .A4(new_n724), .ZN(new_n817));
  INV_X1    g631(.A(new_n691), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT48), .B1(new_n792), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n784), .A2(new_n675), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n805), .A2(new_n263), .A3(new_n582), .A4(new_n808), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n820), .A2(new_n822), .A3(KEYINPUT117), .A4(new_n821), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n814), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n774), .A2(new_n775), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n703), .A2(new_n693), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n752), .A2(KEYINPUT110), .A3(new_n774), .A4(new_n775), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n758), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n750), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT111), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n776), .A2(new_n777), .A3(new_n750), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n834), .A2(new_n839), .A3(new_n750), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n780), .B(new_n828), .C1(KEYINPUT54), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(G952), .A2(G953), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT118), .ZN(new_n844));
  INV_X1    g658(.A(new_n710), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT107), .Z(new_n847));
  AOI211_X1 g661(.A(new_n845), .B(new_n847), .C1(KEYINPUT49), .C2(new_n782), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n628), .B2(new_n797), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n804), .A2(new_n562), .A3(new_n415), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n842), .A2(new_n844), .B1(new_n849), .B2(new_n850), .ZN(G75));
  AOI21_X1  g665(.A(new_n254), .B1(new_n773), .B2(new_n778), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(G210), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n406), .A2(new_n341), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n411), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT55), .Z(new_n856));
  XOR2_X1   g670(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n857));
  AND3_X1   g671(.A1(new_n853), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n856), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n209), .A2(G952), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(G51));
  XNOR2_X1  g676(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n557), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n773), .B2(new_n778), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n780), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n557), .A2(new_n863), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n651), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n852), .A2(G469), .A3(new_n732), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n861), .B1(new_n869), .B2(new_n870), .ZN(G54));
  NAND3_X1  g685(.A1(new_n852), .A2(KEYINPUT58), .A3(G475), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(new_n592), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n592), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(new_n861), .ZN(G60));
  NAND2_X1  g689(.A1(G478), .A2(G902), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT59), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n577), .A2(new_n578), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT121), .Z(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n877), .B(new_n880), .C1(new_n780), .C2(new_n866), .ZN(new_n881));
  INV_X1    g695(.A(new_n861), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n841), .A2(KEYINPUT54), .ZN(new_n884));
  INV_X1    g698(.A(new_n780), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n877), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n887), .B2(new_n879), .ZN(G63));
  NAND2_X1  g702(.A1(G217), .A2(G902), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT60), .Z(new_n890));
  NAND3_X1  g704(.A1(new_n779), .A2(new_n611), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n779), .A2(new_n890), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n882), .B(new_n891), .C1(new_n892), .C2(new_n522), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT61), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n893), .B(new_n895), .ZN(G66));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n209), .B1(new_n748), .B2(new_n771), .ZN(new_n898));
  OAI21_X1  g712(.A(G953), .B1(new_n313), .B2(new_n339), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n406), .B1(G898), .B2(new_n209), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n901), .B(new_n902), .Z(G69));
  AOI21_X1  g717(.A(new_n209), .B1(G227), .B2(G900), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n456), .B(new_n241), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n746), .A2(new_n649), .A3(new_n626), .A4(new_n677), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n719), .A2(new_n727), .A3(new_n726), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n691), .B1(new_n669), .B2(new_n670), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n911), .B2(new_n739), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n752), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n752), .A3(KEYINPUT124), .ZN(new_n916));
  AOI21_X1  g730(.A(G953), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n209), .A2(G900), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n907), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n912), .A2(new_n752), .A3(KEYINPUT124), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT124), .B1(new_n912), .B2(new_n752), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n209), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n918), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(KEYINPUT125), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n906), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n644), .A2(new_n755), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT62), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n746), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n528), .A2(new_n768), .A3(new_n639), .A4(new_n727), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n740), .A2(new_n929), .ZN(new_n930));
  AOI211_X1 g744(.A(G953), .B(new_n905), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n925), .A2(KEYINPUT126), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n922), .A2(KEYINPUT125), .A3(new_n923), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT125), .B1(new_n922), .B2(new_n923), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n905), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n928), .A2(new_n930), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n209), .A3(new_n906), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n933), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n904), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT126), .B1(new_n925), .B2(new_n931), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n936), .A2(new_n938), .A3(new_n933), .ZN(new_n942));
  INV_X1    g756(.A(new_n904), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n944), .ZN(G72));
  INV_X1    g759(.A(new_n631), .ZN(new_n946));
  NAND2_X1  g760(.A1(G472), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT63), .Z(new_n948));
  NAND2_X1  g762(.A1(new_n457), .A2(new_n442), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n841), .A2(new_n946), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n927), .A2(new_n746), .A3(new_n774), .A4(new_n930), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n946), .B1(new_n951), .B2(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n915), .A2(new_n774), .A3(new_n916), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n949), .B1(new_n953), .B2(new_n948), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n952), .A2(new_n954), .A3(new_n861), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT127), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n950), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(G57));
endmodule


