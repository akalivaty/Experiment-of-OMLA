//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  AOI21_X1  g004(.A(KEYINPUT67), .B1(new_n190), .B2(G119), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(G119), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT69), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n194), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n187), .B1(new_n188), .B2(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n188), .A2(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n200), .A4(new_n189), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n195), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n193), .A2(KEYINPUT68), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n204), .A3(new_n189), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n196), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT70), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n205), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n194), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT70), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n195), .A2(new_n201), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(G137), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n215), .A2(new_n218), .A3(new_n221), .A4(new_n216), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G143), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT65), .A3(G146), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n226), .A2(new_n228), .B1(G143), .B2(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(KEYINPUT64), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n225), .A2(G143), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(G146), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n229), .A2(new_n231), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  INV_X1    g053(.A(new_n228), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT65), .B1(new_n227), .B2(G146), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n234), .B(new_n239), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n234), .A2(new_n235), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G128), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(G143), .B2(new_n225), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n243), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n217), .A2(G134), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n214), .A2(G137), .ZN(new_n253));
  OAI21_X1  g067(.A(G131), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n222), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n223), .A2(new_n237), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n207), .A2(new_n212), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n207), .A2(new_n212), .A3(new_n259), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n256), .B(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n207), .A2(new_n212), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n267));
  NOR2_X1   g081(.A1(G237), .A2(G953), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT29), .B1(new_n266), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n257), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n256), .B1(new_n207), .B2(new_n212), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n258), .B2(new_n260), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n278), .B2(new_n275), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n274), .B1(new_n279), .B2(new_n273), .ZN(new_n280));
  INV_X1    g094(.A(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT28), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n282), .A2(KEYINPUT29), .A3(new_n276), .A4(new_n272), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT73), .B(G902), .Z(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n280), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G472), .ZN(new_n287));
  INV_X1    g101(.A(G472), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n261), .A2(new_n272), .A3(new_n265), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n261), .A2(KEYINPUT31), .A3(new_n272), .A4(new_n265), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n279), .A2(new_n273), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n290), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT32), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT32), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n293), .A2(new_n294), .B1(new_n279), .B2(new_n273), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n290), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n287), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G469), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT79), .B(G107), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(G104), .ZN(new_n305));
  INV_X1    g119(.A(G104), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G107), .ZN(new_n307));
  OAI21_X1  g121(.A(G101), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n309));
  AND2_X1   g123(.A1(KEYINPUT79), .A2(G107), .ZN(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT79), .A2(G107), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n309), .B(G104), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G101), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n306), .A2(G107), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n306), .B2(G107), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n251), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n238), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n249), .A2(KEYINPUT80), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n229), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n242), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n316), .B(new_n308), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n223), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT12), .ZN(new_n329));
  INV_X1    g143(.A(new_n317), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT10), .A3(new_n251), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT10), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n223), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G101), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT4), .A3(new_n316), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n338), .A3(G101), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n237), .A3(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n331), .A2(new_n333), .A3(new_n334), .A4(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT12), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n327), .A2(new_n342), .A3(new_n223), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n329), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G110), .B(G140), .ZN(new_n345));
  INV_X1    g159(.A(G227), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n345), .B(new_n347), .Z(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n331), .A2(new_n333), .A3(new_n340), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n223), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n352), .B2(new_n341), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n303), .B(new_n285), .C1(new_n350), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(G469), .A2(G902), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n344), .A2(new_n349), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n341), .A3(new_n348), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n354), .B(new_n355), .C1(new_n358), .C2(new_n303), .ZN(new_n359));
  INV_X1    g173(.A(G221), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT9), .B(G234), .Z(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(new_n289), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n268), .A2(G143), .A3(G214), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(G143), .B1(new_n268), .B2(G214), .ZN(new_n367));
  OAI21_X1  g181(.A(G131), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n221), .A3(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT88), .B1(new_n371), .B2(KEYINPUT17), .ZN(new_n372));
  INV_X1    g186(.A(G125), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n373), .A2(KEYINPUT16), .A3(G140), .ZN(new_n374));
  INV_X1    g188(.A(G140), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n373), .B2(KEYINPUT76), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(G125), .A3(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n374), .B1(new_n379), .B2(KEYINPUT16), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(G146), .ZN(new_n381));
  AOI211_X1 g195(.A(new_n225), .B(new_n374), .C1(new_n379), .C2(KEYINPUT16), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n369), .A2(new_n365), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT17), .A3(G131), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT88), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT17), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n368), .A2(new_n370), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n372), .A2(new_n383), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT18), .A2(G131), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n384), .B(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G125), .B(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n225), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n376), .A2(G146), .A3(new_n378), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n391), .B(new_n396), .C1(new_n394), .C2(new_n395), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G113), .B(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n306), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n398), .B(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G475), .B1(new_n401), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n382), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n392), .A2(KEYINPUT19), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(KEYINPUT19), .B2(new_n379), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n403), .B(new_n404), .C1(G146), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n405), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n379), .A2(KEYINPUT19), .ZN(new_n409));
  AOI21_X1  g223(.A(G146), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT87), .B1(new_n410), .B2(new_n382), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n411), .A3(new_n371), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n397), .ZN(new_n413));
  INV_X1    g227(.A(new_n400), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n414), .B2(new_n398), .ZN(new_n416));
  INV_X1    g230(.A(G475), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(KEYINPUT20), .A3(new_n417), .A4(new_n289), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n398), .A2(new_n414), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n400), .B1(new_n412), .B2(new_n397), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n417), .B(new_n289), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n402), .A2(new_n418), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT15), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G478), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n238), .A2(G143), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n227), .B1(new_n244), .B2(new_n246), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT13), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n427), .B(new_n429), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n247), .A2(G143), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n428), .B1(new_n433), .B2(KEYINPUT13), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT89), .B1(new_n429), .B2(new_n431), .ZN(new_n435));
  OAI211_X1 g249(.A(G134), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n304), .B(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n433), .A2(new_n214), .A3(new_n429), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G122), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G116), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(G116), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT14), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT90), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n444), .ZN(new_n448));
  OAI211_X1 g262(.A(KEYINPUT90), .B(new_n442), .C1(new_n443), .C2(new_n444), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G107), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n304), .A2(new_n437), .ZN(new_n452));
  OAI21_X1  g266(.A(G134), .B1(new_n430), .B2(new_n428), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n439), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n440), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G953), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n361), .A2(G217), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT91), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT92), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n460), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n440), .A2(new_n455), .A3(new_n463), .A4(new_n459), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n285), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n465), .B2(new_n285), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n426), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n425), .A3(G478), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n424), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n364), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT23), .B1(new_n238), .B2(G119), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n238), .A2(G119), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AND4_X1   g291(.A1(KEYINPUT75), .A2(new_n247), .A3(KEYINPUT23), .A4(G119), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n188), .B1(new_n244), .B2(new_n246), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT75), .B1(new_n479), .B2(KEYINPUT23), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT78), .B(G110), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n479), .A2(new_n476), .ZN(new_n483));
  OR2_X1    g297(.A1(KEYINPUT24), .A2(G110), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT24), .A2(G110), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT74), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(KEYINPUT74), .A3(new_n485), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI22_X1  g304(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n403), .A3(new_n393), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n481), .A2(G110), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n380), .B(G146), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n483), .A2(new_n488), .A3(new_n489), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AND4_X1   g310(.A1(KEYINPUT77), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n481), .B2(G110), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT77), .B1(new_n498), .B2(new_n494), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n492), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n457), .A2(G221), .A3(G234), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT22), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(G137), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n492), .B(new_n503), .C1(new_n497), .C2(new_n499), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G234), .ZN(new_n508));
  OAI21_X1  g322(.A(G217), .B1(new_n284), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n507), .A2(G902), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n285), .A3(new_n506), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT25), .A4(new_n285), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n511), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  OAI21_X1  g331(.A(G214), .B1(G237), .B2(G902), .ZN(new_n518));
  INV_X1    g332(.A(G952), .ZN(new_n519));
  AOI211_X1 g333(.A(G953), .B(new_n519), .C1(G234), .C2(G237), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G237), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n284), .B(G953), .C1(new_n508), .C2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT21), .B(G898), .Z(new_n524));
  OAI21_X1  g338(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G113), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT5), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n192), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n208), .B2(new_n527), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n330), .A2(new_n529), .A3(new_n211), .ZN(new_n530));
  XOR2_X1   g344(.A(G110), .B(G122), .Z(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n207), .A2(new_n212), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n337), .A2(new_n339), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n530), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n207), .B2(new_n212), .ZN(new_n536));
  INV_X1    g350(.A(new_n530), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n538), .A3(KEYINPUT6), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n540), .B(new_n531), .C1(new_n536), .C2(new_n537), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n232), .A2(new_n236), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n234), .B(new_n231), .C1(new_n240), .C2(new_n241), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n542), .A2(new_n543), .A3(G125), .ZN(new_n544));
  AOI21_X1  g358(.A(G125), .B1(new_n242), .B2(new_n250), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT81), .B(G224), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n457), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n548), .B(KEYINPUT82), .Z(new_n549));
  XNOR2_X1  g363(.A(new_n546), .B(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n539), .A2(new_n541), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT7), .B(new_n548), .C1(new_n544), .C2(new_n545), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT85), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n536), .A2(new_n537), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(new_n532), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n528), .B1(new_n193), .B2(new_n527), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n330), .A2(new_n211), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT83), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n529), .A2(new_n211), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n317), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT83), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n330), .A2(new_n561), .A3(new_n211), .A4(new_n556), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n531), .B(KEYINPUT8), .Z(new_n564));
  OR2_X1    g378(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n548), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n563), .A2(new_n564), .B1(new_n546), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n555), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G210), .B1(G237), .B2(G902), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n551), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n551), .B2(new_n569), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n518), .B(new_n525), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n302), .A2(new_n473), .A3(new_n517), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G101), .ZN(G3));
  NAND2_X1  g390(.A1(new_n465), .A2(new_n285), .ZN(new_n577));
  INV_X1    g391(.A(G478), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT96), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n581), .A3(new_n578), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n456), .A2(new_n583), .A3(new_n460), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT95), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n459), .A2(KEYINPUT94), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT33), .B1(new_n456), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n465), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n588), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT95), .B1(new_n592), .B2(new_n584), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n589), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n285), .A2(G478), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n580), .B(new_n582), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n402), .A2(new_n418), .A3(new_n423), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n573), .ZN(new_n599));
  INV_X1    g413(.A(new_n297), .ZN(new_n600));
  OAI21_X1  g414(.A(G472), .B1(new_n300), .B2(new_n284), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n517), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n364), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT34), .B(G104), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G6));
  INV_X1    g420(.A(new_n469), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n607), .A2(new_n467), .B1(new_n425), .B2(G478), .ZN(new_n608));
  INV_X1    g422(.A(new_n471), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n424), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n573), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n602), .A2(new_n611), .A3(new_n603), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT35), .B(G107), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G9));
  AOI21_X1  g428(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n615));
  OAI22_X1  g429(.A1(new_n615), .A2(new_n288), .B1(new_n290), .B2(new_n300), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n504), .A2(KEYINPUT36), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n500), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n500), .A2(new_n619), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n289), .A2(new_n620), .A3(new_n509), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n574), .A3(new_n473), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  OAI21_X1  g441(.A(new_n518), .B1(new_n571), .B2(new_n572), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n597), .B1(new_n470), .B2(new_n471), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n521), .B1(new_n523), .B2(G900), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n302), .A2(new_n629), .A3(new_n635), .A4(new_n603), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  XNOR2_X1  g451(.A(new_n634), .B(KEYINPUT39), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n359), .A2(new_n363), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n289), .B1(new_n281), .B2(new_n272), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n273), .B1(new_n261), .B2(new_n265), .ZN(new_n643));
  OAI21_X1  g457(.A(G472), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n298), .A2(new_n301), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n424), .B1(new_n470), .B2(new_n471), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n551), .A2(new_n569), .ZN(new_n648));
  INV_X1    g462(.A(new_n570), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n551), .A2(new_n569), .A3(new_n570), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT38), .ZN(new_n653));
  INV_X1    g467(.A(new_n518), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n617), .A2(new_n654), .A3(new_n622), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n641), .A2(new_n647), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT98), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  AND2_X1   g472(.A1(new_n302), .A2(new_n629), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n580), .A2(new_n582), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n591), .A2(new_n593), .ZN(new_n661));
  INV_X1    g475(.A(new_n589), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n595), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n597), .B(new_n634), .C1(new_n660), .C2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n596), .A2(KEYINPUT99), .A3(new_n597), .A4(new_n634), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n659), .A2(new_n668), .A3(new_n603), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G146), .ZN(G48));
  OAI21_X1  g484(.A(new_n285), .B1(new_n350), .B2(new_n353), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G469), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n363), .A3(new_n354), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n599), .A2(new_n302), .A3(new_n517), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND4_X1  g491(.A1(new_n611), .A2(new_n302), .A3(new_n517), .A4(new_n674), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  INV_X1    g493(.A(new_n472), .ZN(new_n680));
  INV_X1    g494(.A(new_n525), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n302), .A2(new_n629), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G119), .ZN(G21));
  AOI21_X1  g498(.A(new_n654), .B1(new_n650), .B2(new_n651), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n682), .A2(new_n685), .A3(new_n646), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n295), .A2(new_n296), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n285), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n297), .B1(new_n689), .B2(G472), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n687), .B1(new_n690), .B2(new_n517), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n687), .A2(new_n517), .A3(new_n600), .A4(new_n601), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n686), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  NOR2_X1   g508(.A1(new_n628), .A2(new_n673), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n624), .A2(new_n666), .A3(new_n667), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G125), .ZN(G27));
  NAND3_X1  g511(.A1(new_n650), .A2(new_n518), .A3(new_n651), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n356), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n344), .A2(KEYINPUT101), .A3(new_n349), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(G469), .A3(new_n357), .A4(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n354), .A3(new_n355), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n698), .A2(new_n703), .A3(new_n362), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n298), .A2(KEYINPUT102), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n297), .A2(new_n706), .A3(KEYINPUT32), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n705), .A2(new_n301), .A3(new_n287), .A4(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n668), .A2(new_n517), .A3(new_n704), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n704), .A2(new_n302), .A3(new_n517), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n666), .A2(new_n667), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(KEYINPUT42), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n709), .A2(KEYINPUT42), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G131), .ZN(G33));
  NAND4_X1  g529(.A1(new_n704), .A2(new_n302), .A3(new_n635), .A4(new_n517), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G134), .ZN(G36));
  NOR2_X1   g531(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n596), .A2(new_n424), .ZN(new_n720));
  NAND2_X1  g534(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n596), .A2(new_n424), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n718), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n690), .B(new_n623), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n698), .B1(new_n726), .B2(KEYINPUT44), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n357), .A4(new_n701), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n358), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(G469), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT46), .B1(new_n731), .B2(new_n355), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n732), .A2(KEYINPUT104), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n355), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n734), .A2(KEYINPUT103), .ZN(new_n735));
  INV_X1    g549(.A(new_n354), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n732), .B2(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(KEYINPUT103), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n733), .A2(new_n735), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n363), .A3(new_n638), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n727), .B(new_n740), .C1(KEYINPUT44), .C2(new_n726), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G137), .ZN(G39));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n739), .B2(new_n363), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n517), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n739), .A2(new_n743), .A3(new_n363), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n712), .A2(new_n302), .A3(new_n698), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G140), .ZN(G42));
  AOI21_X1  g564(.A(new_n521), .B1(new_n723), .B2(new_n725), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n698), .A2(new_n673), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n753), .A2(new_n616), .A3(new_n623), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n298), .A2(new_n301), .A3(new_n644), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n520), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n752), .A2(new_n517), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n756), .A2(new_n757), .A3(new_n597), .A4(new_n596), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n691), .A2(new_n692), .ZN(new_n759));
  INV_X1    g573(.A(new_n653), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n673), .A2(new_n518), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT114), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n759), .A2(new_n751), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n754), .B(new_n758), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  OR2_X1    g581(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n769));
  INV_X1    g583(.A(new_n747), .ZN(new_n770));
  INV_X1    g584(.A(new_n672), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n736), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT112), .ZN(new_n773));
  OAI22_X1  g587(.A1(new_n770), .A2(new_n744), .B1(new_n363), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n698), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n759), .A2(new_n751), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n708), .A2(new_n517), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n753), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT48), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n776), .A2(new_n695), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n781), .A2(new_n519), .A3(G953), .A4(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n777), .A2(KEYINPUT113), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n774), .A2(new_n786), .A3(new_n775), .A4(new_n776), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n785), .B(new_n787), .C1(new_n767), .C2(KEYINPUT115), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n769), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n675), .A2(new_n693), .A3(new_n678), .A4(new_n683), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT106), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n685), .A2(new_n791), .A3(new_n630), .A4(new_n525), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT106), .B1(new_n573), .B2(new_n610), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n602), .A4(new_n603), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(new_n575), .A3(new_n604), .A4(new_n625), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n704), .A2(new_n624), .A3(new_n666), .A4(new_n667), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n623), .A2(new_n698), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n302), .A2(new_n798), .A3(new_n473), .A4(new_n634), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n716), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n714), .A2(new_n790), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n302), .A2(new_n629), .A3(new_n603), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n696), .B(new_n636), .C1(new_n803), .C2(new_n712), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n703), .A2(new_n362), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n634), .B(KEYINPUT107), .Z(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT108), .B1(new_n623), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n617), .A2(new_n622), .A3(new_n809), .A4(new_n806), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n805), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n645), .A2(new_n685), .A3(new_n646), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT52), .B1(new_n804), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n659), .B(new_n603), .C1(new_n668), .C2(new_n635), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n646), .A2(new_n685), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n755), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n817), .B(new_n805), .C1(new_n808), .C2(new_n810), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n815), .A2(new_n818), .A3(new_n819), .A4(new_n696), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n802), .A2(KEYINPUT53), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n693), .A2(new_n675), .A3(new_n678), .A4(new_n683), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n795), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n714), .A3(new_n801), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n814), .A2(new_n820), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n822), .A2(KEYINPUT109), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT109), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n802), .A2(new_n830), .A3(new_n821), .A4(KEYINPUT53), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(KEYINPUT54), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n824), .A2(new_n795), .A3(new_n800), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n714), .A3(new_n814), .A4(new_n820), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n833), .B1(new_n835), .B2(new_n823), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n802), .A2(KEYINPUT110), .A3(new_n821), .A4(KEYINPUT53), .ZN(new_n837));
  XNOR2_X1  g651(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n836), .A2(new_n837), .A3(new_n828), .A4(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n784), .A2(new_n789), .A3(new_n832), .A4(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n756), .A2(new_n757), .A3(new_n598), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n841), .A2(new_n842), .B1(G952), .B2(G953), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n746), .A2(new_n724), .A3(new_n654), .A4(new_n362), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n772), .B(KEYINPUT49), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n760), .A2(new_n844), .A3(new_n755), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(G75));
  NOR2_X1   g661(.A1(new_n457), .A2(G952), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT116), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n836), .A2(new_n828), .A3(new_n837), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n284), .A3(new_n649), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n539), .A2(new_n541), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(new_n550), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT55), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n856), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(G51));
  NAND2_X1  g673(.A1(new_n850), .A2(new_n838), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n840), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n355), .B(KEYINPUT57), .Z(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n350), .A2(new_n353), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT117), .Z(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n731), .B(KEYINPUT118), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n850), .A2(new_n284), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n848), .B1(new_n866), .B2(new_n868), .ZN(G54));
  AND2_X1   g683(.A1(KEYINPUT58), .A2(G475), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n850), .A2(new_n284), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n416), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n848), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n850), .A2(new_n284), .A3(new_n416), .A4(new_n870), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n873), .A2(new_n878), .A3(new_n874), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(G60));
  NAND2_X1  g694(.A1(G478), .A2(G902), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT59), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n594), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n861), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n849), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n832), .B2(new_n840), .ZN(new_n887));
  INV_X1    g701(.A(new_n594), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT120), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n832), .A2(new_n840), .ZN(new_n890));
  INV_X1    g704(.A(new_n882), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n594), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n886), .B1(new_n889), .B2(new_n894), .ZN(G63));
  NAND2_X1  g709(.A1(G217), .A2(G902), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT121), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT60), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n850), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n507), .B(KEYINPUT122), .Z(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n850), .A2(new_n620), .A3(new_n621), .A4(new_n898), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n885), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n901), .A2(KEYINPUT61), .A3(new_n885), .A4(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(G66));
  NAND2_X1  g721(.A1(new_n524), .A2(new_n547), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(G953), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n825), .B2(G953), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n854), .B1(G898), .B2(new_n457), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(G69));
  AND2_X1   g726(.A1(new_n741), .A2(new_n749), .ZN(new_n913));
  INV_X1    g727(.A(new_n804), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n714), .A2(new_n716), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n779), .A2(new_n816), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n740), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n263), .B(KEYINPUT123), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(new_n406), .Z(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(G953), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n639), .A2(new_n698), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n598), .A2(new_n610), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(new_n302), .A3(new_n517), .A4(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT124), .Z(new_n926));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n927));
  INV_X1    g741(.A(new_n656), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n804), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n815), .A2(KEYINPUT62), .A3(new_n656), .A4(new_n696), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n741), .A3(new_n749), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n457), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n920), .ZN(new_n934));
  INV_X1    g748(.A(G900), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(G953), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n922), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT125), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n346), .B2(new_n935), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n922), .A2(new_n934), .A3(new_n940), .A4(new_n936), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n938), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(G72));
  NAND2_X1  g758(.A1(G472), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT63), .Z(new_n946));
  INV_X1    g760(.A(new_n825), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n918), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n266), .A2(new_n272), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n848), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n946), .B1(new_n932), .B2(new_n947), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT126), .B(new_n946), .C1(new_n932), .C2(new_n947), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(new_n643), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n643), .ZN(new_n957));
  INV_X1    g771(.A(new_n949), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n829), .A2(new_n957), .A3(new_n831), .A4(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n946), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT127), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n964), .A3(new_n950), .A4(new_n955), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(G57));
endmodule


