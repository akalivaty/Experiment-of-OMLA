//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G353));
  NOR2_X1   g0007(.A1(G97), .A2(G107), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(new_n203), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(G20), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(new_n220), .B2(new_n219), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n216), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n223), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n253), .A2(G223), .B1(G77), .B2(new_n251), .ZN(new_n254));
  INV_X1    g0054(.A(G222), .ZN(new_n255));
  OR2_X1    g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  AOI21_X1  g0057(.A(G1698), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n214), .B2(new_n261), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OR2_X1    g0067(.A1(KEYINPUT68), .A2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT68), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n266), .B(new_n267), .C1(G45), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(G226), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G190), .ZN(new_n278));
  XOR2_X1   g0078(.A(KEYINPUT71), .B(G200), .Z(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT10), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n284), .A2(new_n213), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n267), .A2(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G50), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n287), .A2(new_n289), .B1(G50), .B2(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G150), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  INV_X1    g0095(.A(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G33), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n294), .B1(new_n295), .B2(new_n297), .C1(new_n204), .C2(new_n296), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n284), .A2(new_n213), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n282), .A2(new_n283), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n303), .A2(new_n278), .A3(new_n305), .A4(new_n281), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n274), .A2(G244), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n271), .A2(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n253), .A2(G238), .B1(G107), .B2(new_n251), .ZN(new_n312));
  INV_X1    g0112(.A(G232), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n259), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n314), .B2(new_n263), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n315), .A2(G190), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n279), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n287), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n286), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n299), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT70), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(G77), .A3(new_n288), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n205), .ZN(new_n325));
  INV_X1    g0125(.A(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n296), .A2(new_n326), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n295), .A2(new_n327), .B1(new_n296), .B2(new_n205), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n297), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n299), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n324), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n316), .A2(new_n317), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(G169), .B2(new_n315), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n315), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n333), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n277), .A2(G169), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n276), .A2(G179), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n342), .A2(new_n343), .A3(new_n302), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n258), .A2(G223), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G87), .ZN(new_n347));
  INV_X1    g0147(.A(G226), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n256), .A2(new_n257), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n263), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n274), .A2(G232), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n271), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(new_n336), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n352), .B2(new_n354), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n295), .B1(new_n267), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n321), .B1(new_n320), .B2(new_n295), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n256), .A2(new_n296), .A3(new_n257), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n296), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G58), .A2(G68), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n296), .B1(new_n203), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G159), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n327), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT76), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(G58), .A2(G68), .ZN(new_n373));
  NOR2_X1   g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n293), .A2(G159), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n367), .A2(G68), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n285), .B1(new_n379), .B2(KEYINPUT16), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n202), .B1(new_n365), .B2(new_n366), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n375), .A2(new_n377), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n362), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT18), .B1(new_n359), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n358), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n336), .B2(new_n355), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n372), .A2(new_n378), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n251), .B2(new_n296), .ZN(new_n391));
  NOR4_X1   g0191(.A1(new_n249), .A2(new_n250), .A3(new_n364), .A4(G20), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n390), .A2(new_n393), .A3(KEYINPUT16), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n384), .A2(new_n394), .A3(new_n299), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n361), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n355), .A2(G200), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n352), .A2(new_n354), .A3(G190), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(new_n395), .A3(new_n361), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n385), .A2(KEYINPUT17), .A3(new_n399), .A4(new_n398), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n386), .A2(new_n397), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n309), .A2(new_n341), .A3(new_n345), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n274), .A2(G238), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n271), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n313), .A2(G1698), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n409), .B1(G226), .B2(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n262), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT13), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n411), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n263), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(new_n271), .A4(new_n407), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n413), .A2(new_n417), .A3(G179), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT73), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n413), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(KEYINPUT73), .B(KEYINPUT13), .C1(new_n408), .C2(new_n412), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G169), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n420), .A2(KEYINPUT14), .A3(G169), .A4(new_n421), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n418), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n202), .A2(G20), .ZN(new_n427));
  INV_X1    g0227(.A(G50), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n427), .B1(new_n297), .B2(new_n205), .C1(new_n428), .C2(new_n327), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n299), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT11), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT11), .B1(new_n436), .B2(new_n431), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n323), .A2(G68), .A3(new_n288), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n320), .A2(new_n202), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT12), .ZN(new_n440));
  AND4_X1   g0240(.A1(new_n435), .A2(new_n437), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n426), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n420), .A2(G200), .A3(new_n421), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT74), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT74), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n420), .A2(new_n445), .A3(G200), .A4(new_n421), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n413), .A2(new_n417), .A3(G190), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n444), .A2(new_n441), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n406), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT77), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT77), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(G33), .A3(G283), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n349), .A2(G250), .A3(G1698), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT4), .B1(new_n258), .B2(G244), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n263), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n267), .B(G45), .C1(new_n461), .C2(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n270), .B2(new_n461), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n263), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(G257), .B1(new_n266), .B2(new_n463), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G200), .ZN(new_n467));
  INV_X1    g0267(.A(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(KEYINPUT6), .A3(G97), .ZN(new_n469));
  XOR2_X1   g0269(.A(G97), .B(G107), .Z(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(KEYINPUT6), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(G20), .B1(G77), .B2(new_n293), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n367), .A2(G107), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n299), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n286), .A2(G97), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n287), .B1(new_n267), .B2(G33), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(G97), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n460), .A2(new_n465), .A3(G190), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n467), .A2(new_n475), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(new_n478), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n466), .A2(new_n357), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n460), .A2(new_n465), .A3(new_n336), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G20), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n296), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n468), .A2(KEYINPUT23), .A3(G20), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n296), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT24), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n491), .C1(new_n493), .C2(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n299), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n463), .A2(new_n266), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n464), .A2(G264), .ZN(new_n502));
  OAI211_X1 g0302(.A(G257), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G294), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n349), .A2(G250), .A3(new_n252), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT80), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n258), .A2(KEYINPUT80), .A3(G250), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n501), .B(new_n502), .C1(new_n510), .C2(new_n262), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  INV_X1    g0312(.A(new_n505), .ZN(new_n513));
  INV_X1    g0313(.A(G250), .ZN(new_n514));
  NOR4_X1   g0314(.A1(new_n251), .A2(new_n507), .A3(new_n514), .A4(G1698), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT80), .B1(new_n258), .B2(G250), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n263), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(G190), .A3(new_n501), .A4(new_n502), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT25), .B1(new_n320), .B2(new_n468), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n320), .A2(KEYINPUT25), .A3(new_n468), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n477), .A2(G107), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n500), .A2(new_n512), .A3(new_n519), .A4(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT79), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n349), .A2(G244), .A3(G1698), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n349), .A2(G238), .A3(new_n252), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n486), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n263), .ZN(new_n530));
  INV_X1    g0330(.A(G45), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n514), .B1(new_n531), .B2(G1), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n267), .A2(new_n265), .A3(G45), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n262), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G190), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n349), .A2(new_n296), .A3(G68), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n296), .B1(new_n411), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(G87), .B2(new_n209), .ZN(new_n541));
  INV_X1    g0341(.A(G97), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n539), .B1(new_n297), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n538), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n299), .B1(new_n320), .B2(new_n329), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n477), .A2(G87), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n534), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n529), .B2(new_n263), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(KEYINPUT79), .A3(G190), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n535), .A2(new_n280), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n537), .A2(new_n547), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n549), .A2(G169), .ZN(new_n553));
  AOI211_X1 g0353(.A(G179), .B(new_n548), .C1(new_n529), .C2(new_n263), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n477), .ZN(new_n556));
  XOR2_X1   g0356(.A(new_n329), .B(KEYINPUT78), .Z(new_n557));
  OAI21_X1  g0357(.A(new_n545), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n485), .A2(new_n525), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n511), .A2(new_n357), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n518), .A2(new_n336), .A3(new_n501), .A4(new_n502), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n285), .B1(new_n496), .B2(new_n498), .ZN(new_n564));
  INV_X1    g0364(.A(new_n523), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G116), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n284), .A2(new_n213), .B1(G20), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n456), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n296), .B1(new_n542), .B2(G33), .ZN(new_n571));
  OAI211_X1 g0371(.A(KEYINPUT20), .B(new_n569), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT20), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n571), .B1(new_n453), .B2(new_n455), .ZN(new_n574));
  INV_X1    g0374(.A(new_n569), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n568), .B1(new_n267), .B2(G33), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n319), .A2(new_n322), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n320), .A2(new_n568), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G264), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n582));
  OAI211_X1 g0382(.A(G257), .B(new_n252), .C1(new_n249), .C2(new_n250), .ZN(new_n583));
  INV_X1    g0383(.A(G303), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n349), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n263), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT5), .B1(new_n268), .B2(new_n269), .ZN(new_n587));
  OAI211_X1 g0387(.A(G270), .B(new_n262), .C1(new_n587), .C2(new_n462), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n501), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n581), .A2(G169), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n589), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n581), .A3(G179), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n581), .A2(KEYINPUT21), .A3(G169), .A4(new_n589), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n567), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n589), .A2(new_n536), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n581), .B(new_n598), .C1(G200), .C2(new_n589), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n450), .A2(new_n561), .A3(new_n600), .ZN(G372));
  NAND2_X1  g0401(.A1(new_n386), .A2(new_n397), .ZN(new_n602));
  INV_X1    g0402(.A(new_n448), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n340), .A2(new_n337), .A3(new_n335), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n442), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n402), .A2(new_n403), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n309), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n345), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT81), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n595), .A2(new_n594), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n501), .A2(new_n588), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n357), .B1(new_n613), .B2(new_n586), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT21), .B1(new_n614), .B2(new_n581), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n592), .A2(KEYINPUT81), .A3(new_n594), .A4(new_n595), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n566), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n561), .A3(KEYINPUT82), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT82), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n567), .B1(new_n616), .B2(new_n617), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n545), .B(new_n546), .C1(new_n549), .C2(new_n279), .ZN(new_n623));
  AND4_X1   g0423(.A1(KEYINPUT79), .A2(new_n530), .A3(G190), .A4(new_n534), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n625), .A2(new_n537), .B1(new_n558), .B2(new_n555), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(new_n524), .A3(new_n484), .A4(new_n480), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n621), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n560), .B2(new_n484), .ZN(new_n630));
  INV_X1    g0430(.A(new_n484), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(KEYINPUT26), .A3(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n630), .A2(new_n632), .B1(new_n558), .B2(new_n555), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n620), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n450), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n610), .A2(new_n635), .ZN(G369));
  NAND3_X1  g0436(.A1(new_n267), .A2(new_n296), .A3(G13), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(G213), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(G343), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n581), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n616), .B2(new_n617), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n599), .B(new_n644), .C1(new_n596), .C2(new_n643), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G330), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n564), .B2(new_n565), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n567), .B1(new_n524), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n566), .A2(new_n642), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n649), .ZN(new_n654));
  INV_X1    g0454(.A(new_n642), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n650), .A2(new_n596), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(G399));
  NOR3_X1   g0457(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT83), .Z(new_n659));
  INV_X1    g0459(.A(new_n217), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n270), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G1), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n659), .A2(new_n663), .B1(new_n211), .B2(new_n662), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT28), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n634), .A2(new_n655), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT29), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n561), .A2(new_n597), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n633), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n655), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n668), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G330), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n593), .A2(G179), .A3(new_n518), .A4(new_n502), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT30), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n460), .A2(new_n465), .A3(new_n549), .ZN(new_n676));
  OR3_X1    g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n674), .B2(new_n676), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n593), .A2(G179), .A3(new_n549), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n511), .A3(new_n466), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n642), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT31), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT31), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n684), .A3(new_n642), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n600), .A2(new_n561), .A3(new_n655), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n673), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n672), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n665), .B1(new_n691), .B2(G1), .ZN(G364));
  AND2_X1   g0492(.A1(new_n296), .A2(G13), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n267), .B1(new_n693), .B2(G45), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n662), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n645), .B2(G330), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(G330), .B2(new_n645), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n213), .B1(G20), .B2(new_n357), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G179), .A2(G200), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n296), .B1(new_n701), .B2(G190), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n542), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n336), .A2(G200), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n296), .A2(G190), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n536), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI221_X1 g0509(.A(new_n349), .B1(new_n706), .B2(new_n205), .C1(new_n709), .C2(new_n428), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n707), .A2(G190), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n703), .B(new_n710), .C1(G68), .C2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n280), .A2(new_n336), .A3(new_n705), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G107), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n296), .A2(new_n536), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n704), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT87), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(KEYINPUT87), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n280), .A2(new_n336), .A3(new_n716), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n722), .A2(G58), .B1(new_n724), .B2(G87), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n705), .A2(new_n701), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n370), .ZN(new_n727));
  XOR2_X1   g0527(.A(KEYINPUT88), .B(KEYINPUT32), .Z(new_n728));
  XNOR2_X1  g0528(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n712), .A2(new_n715), .A3(new_n725), .A4(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(G283), .A2(new_n714), .B1(new_n724), .B2(G303), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(G322), .ZN(new_n732));
  XNOR2_X1  g0532(.A(KEYINPUT89), .B(G326), .ZN(new_n733));
  INV_X1    g0533(.A(G294), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n709), .A2(new_n733), .B1(new_n734), .B2(new_n702), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT33), .B(G317), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n711), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G311), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n251), .B1(new_n706), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n726), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(G329), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n731), .A2(new_n732), .A3(new_n737), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n700), .B1(new_n730), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n699), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n244), .A2(G45), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n660), .A2(new_n349), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n748), .B(new_n749), .C1(G45), .C2(new_n211), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n349), .A2(new_n217), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT84), .ZN(new_n752));
  XOR2_X1   g0552(.A(G355), .B(KEYINPUT85), .Z(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G116), .B2(new_n217), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT86), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT86), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n750), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n695), .B(new_n743), .C1(new_n747), .C2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n746), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n645), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n698), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(G396));
  NAND2_X1  g0563(.A1(new_n335), .A2(new_n337), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n332), .A2(new_n642), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n764), .A2(new_n339), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n341), .B2(new_n765), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n666), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n333), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n604), .A2(new_n769), .A3(new_n765), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n604), .B2(new_n765), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n634), .A2(new_n771), .A3(new_n655), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n696), .B1(new_n773), .B2(new_n689), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n689), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n699), .A2(new_n744), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT90), .Z(new_n777));
  OAI21_X1  g0577(.A(new_n696), .B1(new_n777), .B2(G77), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n251), .B1(new_n726), .B2(new_n738), .C1(new_n568), .C2(new_n706), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n722), .B2(G294), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n709), .A2(new_n584), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n703), .B(new_n781), .C1(G283), .C2(new_n711), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G87), .A2(new_n714), .B1(new_n724), .B2(G107), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n706), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G159), .B1(G137), .B2(new_n708), .ZN(new_n786));
  INV_X1    g0586(.A(G150), .ZN(new_n787));
  INV_X1    g0587(.A(new_n711), .ZN(new_n788));
  INV_X1    g0588(.A(G143), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n786), .B1(new_n787), .B2(new_n788), .C1(new_n721), .C2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT91), .Z(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT34), .ZN(new_n792));
  INV_X1    g0592(.A(G132), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n349), .B1(new_n702), .B2(new_n201), .C1(new_n793), .C2(new_n726), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n714), .B2(G68), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n792), .B(new_n795), .C1(new_n428), .C2(new_n723), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n791), .A2(KEYINPUT34), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n784), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n778), .B1(new_n798), .B2(new_n699), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n745), .B2(new_n771), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n775), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G384));
  NAND2_X1  g0602(.A1(new_n426), .A2(new_n448), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT93), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n441), .A2(new_n655), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n805), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n807), .B(new_n448), .C1(new_n426), .C2(new_n441), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n804), .B1(new_n803), .B2(new_n805), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n338), .A2(new_n340), .A3(new_n655), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(new_n772), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n394), .A2(new_n299), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT16), .B1(new_n390), .B2(new_n393), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n361), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT94), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n640), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n376), .B1(new_n375), .B2(new_n377), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n381), .B1(new_n823), .B2(new_n382), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n824), .A2(new_n299), .A3(new_n394), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n825), .A2(KEYINPUT94), .A3(new_n361), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n819), .A2(new_n820), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT95), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n819), .A2(KEYINPUT95), .A3(new_n820), .A4(new_n826), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n819), .A2(new_n388), .A3(new_n826), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n829), .A2(new_n400), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT37), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n388), .A2(new_n396), .ZN(new_n834));
  XOR2_X1   g0634(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n835));
  XNOR2_X1  g0635(.A(new_n640), .B(KEYINPUT96), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n396), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n834), .A2(new_n400), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n829), .A2(new_n830), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n404), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n839), .A2(KEYINPUT98), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT98), .ZN(new_n844));
  INV_X1    g0644(.A(new_n838), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n832), .B2(KEYINPUT37), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n818), .B(new_n362), .C1(new_n380), .C2(new_n824), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT94), .B1(new_n825), .B2(new_n361), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT95), .B1(new_n849), .B2(new_n820), .ZN(new_n850));
  INV_X1    g0650(.A(new_n830), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n404), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT38), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n844), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n843), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n839), .A2(new_n852), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n840), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT99), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n843), .A2(new_n854), .B1(new_n856), .B2(new_n840), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT99), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n814), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n602), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n836), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT100), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n855), .A2(KEYINPUT99), .A3(new_n857), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT99), .B1(new_n855), .B2(new_n857), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n813), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT100), .ZN(new_n870));
  INV_X1    g0670(.A(new_n865), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n839), .A2(new_n842), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n405), .A2(new_n837), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n834), .A2(new_n400), .A3(new_n837), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(new_n835), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n840), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n873), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n858), .B2(KEYINPUT39), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n442), .A2(new_n642), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n866), .A2(new_n872), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n671), .A2(new_n667), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n667), .B2(new_n666), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n450), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n610), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n886), .B(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n767), .B1(new_n687), .B2(new_n686), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT101), .ZN(new_n893));
  INV_X1    g0693(.A(new_n810), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n808), .A3(new_n806), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n867), .B2(new_n868), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n873), .A2(new_n878), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n895), .A4(new_n892), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n450), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n687), .B2(new_n686), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n673), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n891), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n909), .A2(KEYINPUT102), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(KEYINPUT102), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n891), .A2(new_n908), .B1(new_n267), .B2(new_n693), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n213), .A2(new_n296), .A3(new_n568), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n471), .B(KEYINPUT92), .Z(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT35), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n917), .B2(new_n916), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n212), .A2(G77), .A3(new_n368), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n428), .A2(G68), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n267), .B(G13), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n913), .A2(new_n920), .A3(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n239), .A2(new_n749), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n925), .B(new_n747), .C1(new_n217), .C2(new_n329), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n695), .B1(new_n926), .B2(KEYINPUT109), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(KEYINPUT109), .B2(new_n926), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n721), .A2(new_n787), .B1(new_n205), .B2(new_n713), .ZN(new_n929));
  INV_X1    g0729(.A(new_n702), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n930), .A2(G68), .B1(G143), .B2(new_n708), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n370), .B2(new_n788), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n723), .A2(new_n201), .ZN(new_n933));
  INV_X1    g0733(.A(G137), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n349), .B1(new_n726), .B2(new_n934), .C1(new_n428), .C2(new_n706), .ZN(new_n935));
  NOR4_X1   g0735(.A1(new_n929), .A2(new_n932), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT110), .Z(new_n937));
  INV_X1    g0737(.A(G317), .ZN(new_n938));
  INV_X1    g0738(.A(G283), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n251), .B1(new_n726), .B2(new_n938), .C1(new_n939), .C2(new_n706), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n713), .A2(new_n542), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(new_n722), .C2(G303), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n930), .A2(G107), .B1(G311), .B2(new_n708), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n734), .B2(new_n788), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n723), .A2(new_n568), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(KEYINPUT46), .B2(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n942), .B(new_n946), .C1(KEYINPUT46), .C2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n937), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n928), .B1(new_n949), .B2(new_n699), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n547), .A2(new_n655), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n559), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n626), .B2(new_n951), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT103), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n950), .B1(new_n760), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n631), .A2(new_n642), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n481), .A2(new_n642), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n480), .A2(new_n484), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n650), .A2(new_n596), .A3(new_n655), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n484), .B1(new_n959), .B2(new_n566), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n961), .A2(KEYINPUT42), .B1(new_n655), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT105), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT42), .B2(new_n961), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(KEYINPUT105), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n955), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n652), .A2(KEYINPUT106), .A3(new_n960), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n967), .B1(new_n968), .B2(new_n955), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n652), .A2(new_n960), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT106), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n971), .A2(new_n976), .A3(new_n975), .A4(new_n973), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n694), .B(KEYINPUT108), .Z(new_n981));
  AOI21_X1  g0781(.A(new_n960), .B1(new_n656), .B2(new_n654), .ZN(new_n982));
  XOR2_X1   g0782(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n656), .A2(new_n654), .A3(new_n960), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT45), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n653), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n652), .B1(new_n984), .B2(new_n987), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n596), .A2(new_n655), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n651), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n656), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(new_n646), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n691), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n661), .B(KEYINPUT41), .Z(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n981), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n956), .B1(new_n980), .B2(new_n999), .ZN(G387));
  INV_X1    g0800(.A(new_n995), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n651), .A2(new_n746), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n785), .A2(G303), .B1(G311), .B2(new_n711), .ZN(new_n1003));
  INV_X1    g0803(.A(G322), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n709), .C1(new_n721), .C2(new_n938), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT48), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n724), .A2(G294), .B1(G283), .B2(new_n930), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT49), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n251), .B1(new_n733), .B2(new_n726), .C1(new_n713), .C2(new_n568), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT112), .B(G150), .Z(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n251), .B1(new_n1017), .B2(new_n740), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n202), .B2(new_n706), .C1(new_n295), .C2(new_n788), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n941), .B(new_n1019), .C1(G77), .C2(new_n724), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n722), .A2(G50), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n557), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n930), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n708), .A2(G159), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT113), .Z(new_n1025));
  NAND4_X1  g0825(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n700), .B1(new_n1015), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n747), .ZN(new_n1028));
  AOI211_X1 g0828(.A(G45), .B(new_n659), .C1(G68), .C2(G77), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n295), .A2(G50), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n749), .C1(new_n531), .C2(new_n236), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n659), .A2(new_n752), .B1(new_n468), .B2(new_n660), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT111), .Z(new_n1035));
  AOI21_X1  g0835(.A(new_n1028), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1027), .A2(new_n695), .A3(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1001), .A2(new_n981), .B1(new_n1002), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n690), .A2(new_n995), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n691), .A2(new_n1001), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n661), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1039), .A2(KEYINPUT114), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1038), .B1(new_n1042), .B2(new_n1043), .ZN(G393));
  INV_X1    g0844(.A(new_n981), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT115), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n989), .A2(new_n1046), .A3(new_n990), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n985), .A2(new_n988), .A3(KEYINPUT115), .A4(new_n653), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n721), .A2(new_n738), .B1(new_n938), .B2(new_n709), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT117), .Z(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT116), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n715), .B1(new_n939), .B2(new_n723), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n251), .B1(new_n726), .B2(new_n1004), .C1(new_n734), .C2(new_n706), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n788), .A2(new_n584), .B1(new_n702), .B2(new_n568), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1053), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n721), .A2(new_n370), .B1(new_n787), .B2(new_n709), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT51), .Z(new_n1061));
  AOI22_X1  g0861(.A1(G87), .A2(new_n714), .B1(new_n724), .B2(G68), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n349), .B1(new_n726), .B2(new_n789), .C1(new_n295), .C2(new_n706), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n702), .A2(new_n205), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n711), .B2(G50), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1059), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n699), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n957), .A2(new_n959), .A3(new_n746), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1028), .B1(G97), .B2(new_n660), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n247), .A2(new_n749), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n695), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1069), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OR3_X1    g0875(.A1(new_n1049), .A2(KEYINPUT118), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT118), .B1(new_n1049), .B2(new_n1075), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1047), .A2(new_n1041), .A3(new_n1048), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n661), .B1(new_n991), .B2(new_n1041), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1078), .A2(new_n1082), .ZN(G390));
  INV_X1    g0883(.A(new_n685), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n684), .B1(new_n681), .B2(new_n642), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NOR4_X1   g0886(.A1(new_n597), .A2(new_n627), .A3(new_n599), .A4(new_n642), .ZN(new_n1087));
  OAI211_X1 g0887(.A(G330), .B(new_n771), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1088), .A2(new_n811), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n879), .B1(new_n861), .B2(new_n874), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n813), .A2(new_n882), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n812), .B1(new_n671), .B2(new_n767), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n895), .A2(KEYINPUT119), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT119), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n811), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1097), .A2(new_n883), .A3(new_n902), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1089), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n883), .A3(new_n902), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n688), .A2(new_n895), .A3(new_n771), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1103), .A2(new_n1045), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n295), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n723), .A2(new_n1016), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n349), .B1(new_n726), .B2(new_n1108), .C1(new_n706), .C2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n722), .B2(G132), .ZN(new_n1111));
  INV_X1    g0911(.A(G128), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n709), .A2(new_n1112), .B1(new_n702), .B2(new_n370), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G137), .B2(new_n711), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n714), .A2(G50), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1107), .A2(new_n1111), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n722), .A2(G116), .B1(G68), .B2(new_n714), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n708), .A2(G283), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1065), .B1(new_n711), .B2(G107), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n251), .B1(new_n726), .B2(new_n734), .C1(new_n542), .C2(new_n706), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n724), .B2(G87), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n696), .B1(new_n1105), .B2(new_n777), .C1(new_n1123), .C2(new_n700), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n881), .B2(new_n744), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1104), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT120), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n688), .A2(new_n450), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n889), .A2(new_n610), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1094), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n895), .A2(KEYINPUT119), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n1088), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1088), .A2(new_n811), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1101), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n772), .A2(new_n812), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1130), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n662), .B1(new_n1103), .B2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1131), .A2(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(new_n1129), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1099), .A2(new_n1144), .A3(new_n1102), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1127), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1102), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n879), .B1(new_n813), .B2(new_n882), .C1(new_n874), .C2(new_n861), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1101), .B1(new_n1148), .B2(new_n1100), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1141), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  AND4_X1   g0950(.A1(new_n1127), .A2(new_n1150), .A3(new_n661), .A4(new_n1145), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1126), .B1(new_n1146), .B2(new_n1151), .ZN(G378));
  NAND2_X1  g0952(.A1(new_n301), .A2(new_n820), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT122), .Z(new_n1154));
  AOI211_X1 g0954(.A(new_n344), .B(new_n1154), .C1(new_n308), .C2(new_n306), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1154), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n309), .B2(new_n345), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1159));
  OR2_X1    g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n903), .A2(G330), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n901), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1162), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1166), .B(new_n1163), .C1(new_n899), .C2(new_n900), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n886), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n860), .A2(new_n862), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT40), .B1(new_n1169), .B2(new_n898), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1166), .B1(new_n1170), .B2(new_n1163), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n869), .A2(new_n871), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n884), .B1(new_n1172), .B2(KEYINPUT100), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n901), .A2(new_n1164), .A3(new_n1162), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1173), .A3(new_n872), .A4(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1168), .A2(new_n1175), .A3(new_n981), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n695), .B1(new_n428), .B2(new_n776), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT121), .Z(new_n1178));
  NOR2_X1   g0978(.A1(new_n349), .A2(new_n270), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n428), .B1(G33), .B2(G41), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G107), .A2(new_n722), .B1(new_n1022), .B2(new_n785), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n788), .A2(new_n542), .B1(new_n709), .B2(new_n568), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1179), .B1(new_n939), .B2(new_n726), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G68), .C2(new_n930), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n724), .A2(G77), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n714), .A2(G58), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1182), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1181), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n721), .A2(new_n1112), .B1(new_n723), .B2(new_n1109), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n706), .A2(new_n934), .B1(new_n702), .B2(new_n787), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n788), .A2(new_n793), .B1(new_n709), .B2(new_n1108), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n714), .A2(G159), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n740), .C2(G124), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1190), .B1(new_n1189), .B2(new_n1188), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1178), .B1(new_n1201), .B2(new_n699), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n1166), .B2(new_n745), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1176), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1145), .A2(new_n1130), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1168), .A2(new_n1175), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1168), .A2(new_n1175), .A3(KEYINPUT57), .A4(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n661), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1204), .B1(new_n1208), .B2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n1143), .A2(new_n1129), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1141), .A2(new_n998), .A3(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1132), .A2(new_n744), .A3(new_n1133), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n696), .B1(new_n777), .B2(G68), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n722), .A2(G283), .B1(new_n724), .B2(G97), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(new_n1023), .C1(new_n205), .C2(new_n713), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n349), .B1(new_n740), .B2(G303), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G116), .A2(new_n711), .B1(new_n708), .B2(G294), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n468), .C2(new_n706), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n722), .A2(G137), .B1(new_n724), .B2(G159), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n349), .B1(new_n726), .B2(new_n1112), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G150), .B2(new_n785), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1187), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n708), .A2(G132), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n702), .B2(new_n428), .C1(new_n788), .C2(new_n1109), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1217), .A2(new_n1220), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1215), .B1(new_n1227), .B2(new_n699), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1140), .A2(new_n981), .B1(new_n1214), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1213), .A2(new_n1229), .ZN(G381));
  NAND2_X1  g1030(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1126), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1081), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1235));
  INV_X1    g1035(.A(G387), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(G375), .A2(new_n1237), .ZN(G407));
  INV_X1    g1038(.A(G213), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(G343), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(G375), .A2(new_n1232), .A3(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT123), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1044(.A(KEYINPUT63), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1204), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1206), .A2(new_n997), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1176), .A2(new_n1203), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1233), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1240), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1141), .A2(new_n661), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT60), .B1(new_n1212), .B2(KEYINPUT124), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1212), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1252), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1229), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n801), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1255), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(new_n1253), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G384), .B(new_n1229), .C1(new_n1260), .C2(new_n1252), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1245), .B1(new_n1251), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1240), .A2(KEYINPUT125), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1258), .A2(new_n1261), .A3(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(G2897), .A3(new_n1240), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1240), .A2(G2897), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1258), .A2(new_n1261), .A3(new_n1267), .A4(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(KEYINPUT126), .A3(new_n1268), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1251), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1262), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G393), .B(new_n762), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(G390), .B2(G387), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1236), .A2(new_n1235), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT127), .B1(new_n1236), .B2(new_n1235), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1276), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1281), .B(new_n1282), .C1(new_n1236), .C2(new_n1235), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(KEYINPUT61), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1263), .A2(new_n1273), .A3(new_n1275), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1250), .A2(new_n1287), .A3(new_n1274), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n1250), .B2(new_n1269), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1250), .B2(new_n1274), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1286), .B1(new_n1292), .B2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(G375), .A2(new_n1233), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1246), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1284), .A2(new_n1246), .A3(new_n1295), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1262), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1297), .A2(new_n1274), .A3(new_n1298), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(G402));
endmodule


