//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1034, new_n1035, new_n1036, new_n1037;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT27), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n211));
  AOI21_X1  g010(.A(G190gat), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT68), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n214));
  NOR3_X1   g013(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT28), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT28), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  AND2_X1   g016(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n216), .B1(new_n220), .B2(KEYINPUT67), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n213), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT28), .B1(new_n212), .B2(new_n214), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(KEYINPUT67), .A3(new_n216), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(KEYINPUT68), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT26), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229));
  INV_X1    g028(.A(G169gat), .ZN(new_n230));
  INV_X1    g029(.A(G176gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n226), .B(new_n228), .C1(new_n232), .C2(new_n227), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n222), .A2(new_n225), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT23), .B1(new_n230), .B2(new_n231), .ZN(new_n236));
  INV_X1    g035(.A(new_n227), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT25), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n226), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n209), .A2(new_n217), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT64), .B(G169gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n230), .A2(KEYINPUT64), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G169gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n247), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT65), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n243), .A2(KEYINPUT66), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n257), .A2(G169gat), .A3(G176gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n237), .B2(new_n236), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n242), .A3(new_n260), .A4(new_n241), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n244), .A2(new_n255), .B1(new_n262), .B2(KEYINPUT25), .ZN(new_n263));
  INV_X1    g062(.A(G134gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G127gat), .ZN(new_n265));
  AND2_X1   g064(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n267));
  OAI21_X1  g066(.A(G120gat), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G120gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G113gat), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n265), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT1), .B1(new_n264), .B2(G127gat), .ZN(new_n272));
  AND2_X1   g071(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n274));
  OAI21_X1  g073(.A(G127gat), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n265), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278));
  INV_X1    g077(.A(new_n270), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n269), .A2(G113gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n271), .A2(new_n272), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n235), .A2(new_n263), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n235), .B2(new_n263), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n207), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT33), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n205), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n284), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n235), .A2(new_n263), .A3(new_n282), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n206), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT34), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(new_n206), .B2(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n294), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n290), .A2(new_n206), .A3(new_n291), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n285), .B(KEYINPUT32), .C1(new_n286), .C2(new_n205), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n289), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n298), .B1(new_n289), .B2(new_n299), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G141gat), .B(G148gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(G155gat), .B2(G162gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G141gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G148gat), .ZN(new_n312));
  INV_X1    g111(.A(G148gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G141gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G155gat), .B(G162gat), .ZN(new_n316));
  INV_X1    g115(.A(G155gat), .ZN(new_n317));
  INV_X1    g116(.A(G162gat), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT2), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n310), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G211gat), .A2(G218gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(G211gat), .A2(G218gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(G197gat), .A2(G204gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G211gat), .B(G218gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G197gat), .B(G204gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n332), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n310), .A2(new_n320), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT29), .B1(new_n333), .B2(new_n337), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(KEYINPUT3), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n340), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n342), .B1(new_n340), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(G22gat), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n343), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n338), .A2(new_n323), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n321), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n338), .B1(new_n322), .B2(new_n323), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n341), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G22gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n340), .A2(new_n345), .A3(new_n342), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n348), .A2(KEYINPUT78), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G78gat), .B(G106gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT31), .B(G50gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n353), .A2(new_n355), .A3(new_n362), .A4(new_n354), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n357), .A2(KEYINPUT79), .A3(new_n361), .A4(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n356), .A2(new_n360), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n369), .A2(new_n348), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n368), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n303), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT35), .ZN(new_n377));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n235), .A2(new_n263), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(new_n323), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n235), .B2(new_n263), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n339), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n379), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n235), .B2(new_n263), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n384), .B(new_n338), .C1(new_n379), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT73), .B(G64gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G92gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT74), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT74), .ZN(new_n394));
  AOI211_X1 g193(.A(new_n394), .B(new_n391), .C1(new_n383), .C2(new_n386), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n383), .A2(KEYINPUT30), .A3(new_n386), .A4(new_n391), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n393), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n391), .A3(new_n386), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT76), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  INV_X1    g205(.A(G85gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n271), .A2(new_n272), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n277), .A2(new_n281), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(new_n343), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n282), .A2(new_n349), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n282), .A2(new_n349), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n282), .B2(new_n349), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(KEYINPUT77), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT77), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n424), .A3(new_n420), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n412), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n415), .A2(new_n322), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n419), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n422), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n432), .A2(new_n433), .A3(new_n411), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n410), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436));
  INV_X1    g235(.A(new_n410), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n433), .A3(new_n411), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n412), .B(new_n428), .C1(new_n423), .C2(new_n425), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n419), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT6), .B(new_n410), .C1(new_n430), .C2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n398), .A2(new_n405), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n398), .A2(new_n405), .A3(new_n443), .A4(KEYINPUT83), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n376), .A2(new_n377), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n298), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n300), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n374), .B1(new_n368), .B2(new_n371), .ZN(new_n453));
  AOI211_X1 g252(.A(KEYINPUT80), .B(new_n370), .C1(new_n366), .C2(new_n367), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n387), .A2(new_n392), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n394), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n387), .A2(KEYINPUT74), .A3(new_n392), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n396), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT75), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n457), .A2(KEYINPUT75), .A3(new_n396), .A4(new_n458), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n443), .A3(new_n462), .A4(new_n405), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT35), .B1(new_n455), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n373), .A2(KEYINPUT81), .A3(new_n375), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n453), .B2(new_n454), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n468), .A3(new_n463), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n387), .A2(KEYINPUT37), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n383), .B2(new_n386), .ZN(new_n472));
  OR3_X1    g271(.A1(new_n470), .A2(new_n391), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n443), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n470), .A2(new_n472), .ZN(new_n477));
  INV_X1    g276(.A(new_n474), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n392), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n475), .A2(new_n476), .A3(new_n399), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n373), .A2(new_n375), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n398), .A2(new_n405), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n432), .A2(KEYINPUT39), .A3(new_n411), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n410), .ZN(new_n484));
  OR3_X1    g283(.A1(new_n416), .A2(new_n417), .A3(new_n412), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(KEYINPUT39), .C1(new_n432), .C2(new_n411), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n484), .A2(KEYINPUT40), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT40), .B1(new_n484), .B2(new_n486), .ZN(new_n488));
  INV_X1    g287(.A(new_n435), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n480), .A2(new_n481), .A3(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT36), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n452), .B2(KEYINPUT36), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n469), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n465), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT84), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n465), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(G8gat), .ZN(new_n503));
  INV_X1    g302(.A(G15gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n354), .ZN(new_n505));
  NAND2_X1  g304(.A1(G15gat), .A2(G22gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT90), .ZN(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n505), .A2(new_n510), .A3(new_n506), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n508), .A2(new_n511), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n509), .A2(KEYINPUT16), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n503), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n514), .B1(new_n508), .B2(new_n511), .ZN(new_n517));
  OAI21_X1  g316(.A(G8gat), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  OR2_X1    g320(.A1(G43gat), .A2(G50gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(G43gat), .A2(G50gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  OR3_X1    g331(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n526), .A3(new_n530), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT87), .B(G36gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G29gat), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n525), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT89), .B(G50gat), .Z(new_n539));
  XOR2_X1   g338(.A(KEYINPUT88), .B(G43gat), .Z(new_n540));
  OAI22_X1  g339(.A1(G43gat), .A2(new_n539), .B1(new_n540), .B2(G50gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n521), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n529), .A2(new_n530), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n543), .A2(new_n533), .B1(G29gat), .B2(new_n536), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n542), .A2(new_n544), .A3(new_n525), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n520), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n519), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n534), .A2(new_n533), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n537), .B1(new_n549), .B2(new_n531), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n524), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n524), .B1(new_n541), .B2(new_n521), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n519), .A2(new_n547), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n520), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(KEYINPUT18), .B(new_n502), .C1(new_n548), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(KEYINPUT93), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n550), .A2(new_n524), .B1(new_n552), .B2(new_n544), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n561), .A3(new_n519), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n502), .B(KEYINPUT13), .Z(new_n563));
  INV_X1    g362(.A(new_n519), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(new_n564), .A3(KEYINPUT93), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n557), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n547), .B1(new_n559), .B2(KEYINPUT17), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n555), .A2(new_n520), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n564), .A2(new_n569), .B1(new_n570), .B2(new_n559), .ZN(new_n571));
  INV_X1    g370(.A(new_n502), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  INV_X1    g374(.A(G197gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT11), .B(G169gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT12), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n567), .B(new_n573), .C1(new_n574), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n557), .A2(new_n574), .A3(new_n566), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n557), .A2(new_n566), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n564), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n559), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT18), .B1(new_n587), .B2(new_n502), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n581), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT94), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n501), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT9), .ZN(new_n598));
  INV_X1    g397(.A(G64gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G57gat), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n599), .A2(G57gat), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G71gat), .B(G78gat), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  OR2_X1    g404(.A1(KEYINPUT95), .A2(G57gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(KEYINPUT95), .A2(G57gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G64gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT96), .A3(new_n600), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n599), .B1(new_n606), .B2(new_n607), .ZN(new_n612));
  INV_X1    g411(.A(new_n600), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G71gat), .A2(G78gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n598), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n619), .A3(new_n598), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n603), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n605), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  AOI211_X1 g422(.A(KEYINPUT98), .B(new_n621), .C1(new_n610), .C2(new_n614), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n604), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n519), .B1(new_n626), .B2(KEYINPUT21), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n629), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n626), .A2(KEYINPUT21), .ZN(new_n636));
  XOR2_X1   g435(.A(G183gat), .B(G211gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n630), .A2(new_n632), .ZN(new_n641));
  INV_X1    g440(.A(new_n631), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n640), .B1(new_n643), .B2(new_n633), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n597), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n638), .B1(new_n634), .B2(new_n635), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n640), .A3(new_n633), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n596), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(G85gat), .A3(G92gat), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT7), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G99gat), .A2(G106gat), .ZN(new_n656));
  INV_X1    g455(.A(G92gat), .ZN(new_n657));
  AOI22_X1  g456(.A1(KEYINPUT8), .A2(new_n656), .B1(new_n407), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n652), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G99gat), .B(G106gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n520), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n538), .B2(new_n545), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n551), .A2(new_n520), .A3(new_n553), .A4(new_n662), .ZN(new_n665));
  NAND2_X1  g464(.A1(G232gat), .A2(G233gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT101), .Z(new_n667));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G190gat), .B(G218gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n664), .A2(new_n665), .A3(new_n669), .A4(new_n671), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n651), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n667), .A2(new_n668), .ZN(new_n676));
  XOR2_X1   g475(.A(G134gat), .B(G162gat), .Z(new_n677));
  XOR2_X1   g476(.A(new_n676), .B(new_n677), .Z(new_n678));
  AND2_X1   g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n673), .A2(new_n651), .A3(new_n674), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n675), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(G230gat), .A2(G233gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n625), .A2(new_n662), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n660), .B(new_n661), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n604), .B(new_n687), .C1(new_n623), .C2(new_n624), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT10), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n686), .A2(new_n695), .A3(new_n688), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n688), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT104), .B1(new_n698), .B2(new_n685), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  INV_X1    g499(.A(new_n685), .ZN(new_n701));
  AOI211_X1 g500(.A(new_n700), .B(new_n701), .C1(new_n696), .C2(new_n697), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n690), .B(new_n694), .C1(new_n699), .C2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n696), .B2(new_n697), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n693), .B1(new_n704), .B2(new_n689), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n649), .A2(new_n650), .A3(new_n684), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n645), .A2(new_n648), .A3(new_n684), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT105), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n593), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n443), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n509), .ZN(G1324gat));
  XNOR2_X1  g513(.A(KEYINPUT16), .B(G8gat), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n715), .B(new_n712), .C1(new_n398), .C2(new_n405), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n717));
  INV_X1    g516(.A(new_n482), .ZN(new_n718));
  OAI21_X1  g517(.A(G8gat), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(G1325gat));
  NOR3_X1   g520(.A1(new_n712), .A2(new_n504), .A3(new_n495), .ZN(new_n722));
  INV_X1    g521(.A(new_n303), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n593), .A2(new_n723), .A3(new_n711), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n504), .B2(new_n724), .ZN(G1326gat));
  NAND2_X1  g524(.A1(new_n466), .A2(new_n468), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n712), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT43), .B(G22gat), .Z(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n465), .A2(new_n496), .A3(new_n499), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n499), .B1(new_n465), .B2(new_n496), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(new_n591), .A3(new_n683), .A4(new_n707), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(new_n443), .A3(new_n649), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  INV_X1    g535(.A(G29gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n730), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n740), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(KEYINPUT45), .A3(new_n738), .ZN(new_n743));
  INV_X1    g542(.A(new_n649), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n469), .A2(new_n745), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n373), .A2(new_n375), .B1(new_n482), .B2(new_n490), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n494), .B1(new_n747), .B2(new_n480), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n466), .A2(new_n468), .A3(new_n463), .A4(KEYINPUT107), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n684), .B1(new_n750), .B2(new_n465), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n744), .B1(new_n751), .B2(KEYINPUT44), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n684), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n731), .A2(new_n732), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(new_n590), .A3(new_n707), .ZN(new_n758));
  OAI21_X1  g557(.A(G29gat), .B1(new_n758), .B2(new_n443), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n743), .A3(new_n759), .ZN(G1328gat));
  OAI21_X1  g559(.A(new_n536), .B1(new_n758), .B2(new_n718), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n501), .A2(new_n592), .A3(new_n684), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(new_n482), .A3(new_n744), .A4(new_n707), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT46), .B1(new_n763), .B2(new_n536), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n734), .A2(new_n649), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n766));
  INV_X1    g565(.A(new_n536), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n482), .A4(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n761), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT108), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n761), .A2(new_n764), .A3(new_n771), .A4(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1329gat));
  INV_X1    g572(.A(new_n540), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n758), .B2(new_n495), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n765), .A2(new_n723), .A3(new_n540), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1330gat));
  INV_X1    g579(.A(new_n539), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n758), .B2(new_n481), .ZN(new_n782));
  INV_X1    g581(.A(new_n726), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n783), .A3(new_n539), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(KEYINPUT48), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n784), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n758), .A2(new_n726), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n781), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n788), .B2(KEYINPUT48), .ZN(G1331gat));
  OAI211_X1 g588(.A(new_n723), .B(new_n377), .C1(new_n453), .C2(new_n454), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n446), .A2(new_n447), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n462), .A2(new_n443), .A3(new_n405), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n481), .A2(new_n461), .A3(new_n793), .A4(new_n452), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n791), .A2(new_n792), .B1(new_n794), .B2(KEYINPUT35), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n749), .A2(new_n495), .A3(new_n492), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n746), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n707), .A2(new_n590), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n797), .A2(new_n709), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n476), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(new_n608), .Z(G1332gat));
  NAND2_X1  g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n482), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT109), .ZN(new_n805));
  NOR2_X1   g604(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n805), .B(new_n806), .Z(G1333gat));
  XOR2_X1   g606(.A(new_n303), .B(KEYINPUT110), .Z(new_n808));
  AOI21_X1  g607(.A(G71gat), .B1(new_n800), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n494), .A2(G71gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n800), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g611(.A1(new_n800), .A2(new_n783), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g613(.A(new_n753), .B1(new_n797), .B2(new_n684), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n498), .A2(new_n500), .A3(new_n754), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n815), .A2(new_n744), .A3(new_n816), .A4(new_n798), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n407), .A3(new_n443), .ZN(new_n818));
  INV_X1    g617(.A(new_n590), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n751), .A2(new_n819), .A3(new_n744), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT51), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n751), .A2(new_n822), .A3(new_n819), .A4(new_n744), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n706), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n476), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n818), .B1(new_n826), .B2(new_n407), .ZN(G1336gat));
  INV_X1    g626(.A(new_n817), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n657), .B1(new_n828), .B2(new_n482), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n718), .A2(G92gat), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n821), .A2(new_n706), .A3(new_n823), .A4(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT52), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n817), .B2(new_n718), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n757), .A2(KEYINPUT112), .A3(new_n482), .A4(new_n798), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(G92gat), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n838));
  AND2_X1   g637(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n837), .A2(KEYINPUT113), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT113), .B1(new_n837), .B2(new_n839), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n833), .B1(new_n840), .B2(new_n841), .ZN(G1337gat));
  INV_X1    g641(.A(G99gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n843), .A3(new_n723), .ZN(new_n844));
  OAI21_X1  g643(.A(G99gat), .B1(new_n817), .B2(new_n495), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1338gat));
  INV_X1    g645(.A(new_n481), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n821), .A2(new_n847), .A3(new_n706), .A4(new_n823), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(G106gat), .ZN(new_n850));
  INV_X1    g649(.A(G106gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n851), .B1(new_n828), .B2(new_n783), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT53), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n854));
  OAI22_X1  g653(.A1(new_n848), .A2(G106gat), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g654(.A(KEYINPUT53), .B(new_n851), .C1(new_n828), .C2(new_n847), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(G1339gat));
  NAND3_X1  g656(.A1(new_n696), .A2(new_n701), .A3(new_n697), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT54), .B(new_n858), .C1(new_n699), .C2(new_n702), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n694), .B1(new_n704), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(KEYINPUT55), .A3(new_n861), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n864), .A2(new_n590), .A3(new_n703), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n573), .A2(new_n557), .A3(new_n566), .A4(new_n580), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n587), .A2(new_n502), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n563), .B1(new_n562), .B2(new_n565), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n579), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n705), .B2(new_n703), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n866), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n684), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n865), .A2(new_n683), .A3(new_n703), .ZN(new_n879));
  INV_X1    g678(.A(new_n871), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n879), .A2(KEYINPUT115), .A3(new_n864), .A4(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n880), .A2(new_n865), .A3(new_n683), .A4(new_n703), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT55), .B1(new_n859), .B2(new_n861), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n649), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n709), .A2(new_n590), .A3(new_n706), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n443), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n455), .A2(new_n482), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n893), .B(new_n590), .C1(new_n267), .C2(new_n266), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n783), .A2(new_n303), .A3(new_n482), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n591), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT117), .B1(new_n898), .B2(G113gat), .ZN(new_n899));
  OAI211_X1 g698(.A(KEYINPUT117), .B(G113gat), .C1(new_n896), .C2(new_n592), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n894), .B1(new_n899), .B2(new_n901), .ZN(G1340gat));
  OAI21_X1  g701(.A(G120gat), .B1(new_n896), .B2(new_n707), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n706), .A2(new_n269), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n892), .B2(new_n904), .ZN(G1341gat));
  NAND3_X1  g704(.A1(new_n893), .A2(KEYINPUT118), .A3(new_n649), .ZN(new_n906));
  INV_X1    g705(.A(G127gat), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n892), .B2(new_n744), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n897), .A2(G127gat), .A3(new_n649), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1342gat));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n683), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n273), .A2(new_n274), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n892), .A2(new_n914), .A3(new_n684), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n916));
  AOI22_X1  g715(.A1(G134gat), .A2(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n893), .A2(new_n683), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n918), .B(KEYINPUT56), .C1(new_n919), .C2(new_n914), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT119), .B1(new_n915), .B2(new_n916), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(G1343gat));
  NOR2_X1   g721(.A1(new_n889), .A2(new_n481), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n494), .A2(new_n443), .A3(new_n482), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n923), .A2(new_n311), .A3(new_n591), .A4(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n924), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n884), .A2(KEYINPUT120), .ZN(new_n928));
  INV_X1    g727(.A(new_n703), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n863), .B1(new_n862), .B2(KEYINPUT120), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n872), .B1(new_n931), .B2(new_n591), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n886), .B1(new_n932), .B2(new_n683), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n744), .ZN(new_n934));
  INV_X1    g733(.A(new_n888), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(KEYINPUT57), .A3(new_n783), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT57), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n938), .B1(new_n889), .B2(new_n481), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n927), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n590), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n926), .B1(new_n941), .B2(G141gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT58), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n311), .B1(new_n940), .B2(new_n591), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n942), .A2(new_n943), .B1(new_n944), .B2(new_n945), .ZN(G1344gat));
  NAND3_X1  g745(.A1(new_n923), .A2(new_n313), .A3(new_n476), .ZN(new_n947));
  OR4_X1    g746(.A1(new_n494), .A2(new_n947), .A3(new_n482), .A4(new_n707), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n949));
  OAI211_X1 g748(.A(KEYINPUT57), .B(new_n847), .C1(new_n887), .C2(new_n888), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n881), .A2(new_n885), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n865), .A2(new_n703), .ZN(new_n954));
  AOI22_X1  g753(.A1(new_n862), .A2(new_n863), .B1(new_n581), .B2(new_n589), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT116), .B(new_n872), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n876), .B1(new_n866), .B2(new_n873), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n953), .B1(new_n958), .B2(new_n684), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n935), .B1(new_n959), .B2(new_n649), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n960), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n847), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n708), .A2(new_n592), .A3(new_n710), .ZN(new_n962));
  OAI22_X1  g761(.A1(new_n932), .A2(new_n683), .B1(new_n884), .B2(new_n883), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n744), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n938), .B1(new_n964), .B2(new_n726), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n952), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n706), .A3(new_n924), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n949), .B1(new_n967), .B2(G148gat), .ZN(new_n968));
  AOI211_X1 g767(.A(KEYINPUT59), .B(new_n313), .C1(new_n940), .C2(new_n706), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n948), .B1(new_n968), .B2(new_n969), .ZN(G1345gat));
  NOR2_X1   g769(.A1(new_n744), .A2(new_n317), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n923), .A2(new_n649), .A3(new_n924), .ZN(new_n972));
  AOI22_X1  g771(.A1(new_n940), .A2(new_n971), .B1(new_n317), .B2(new_n972), .ZN(G1346gat));
  NOR2_X1   g772(.A1(new_n684), .A2(new_n318), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n923), .A2(new_n683), .A3(new_n924), .ZN(new_n975));
  AOI22_X1  g774(.A1(new_n940), .A2(new_n974), .B1(new_n318), .B2(new_n975), .ZN(G1347gat));
  INV_X1    g775(.A(new_n455), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n718), .A2(new_n476), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n252), .A3(new_n590), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n960), .A2(new_n726), .A3(new_n808), .A4(new_n978), .ZN(new_n982));
  OAI21_X1  g781(.A(G169gat), .B1(new_n982), .B2(new_n592), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n983), .A2(KEYINPUT122), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(KEYINPUT122), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(G1348gat));
  AOI21_X1  g785(.A(G176gat), .B1(new_n980), .B2(new_n706), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n982), .A2(new_n231), .A3(new_n707), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(G1349gat));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n990), .B1(new_n982), .B2(new_n744), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n808), .B(new_n978), .C1(new_n887), .C2(new_n888), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n993), .A2(KEYINPUT123), .A3(new_n726), .A4(new_n649), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n991), .A2(new_n994), .A3(G183gat), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n744), .B1(new_n210), .B2(new_n211), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n980), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT60), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT60), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n995), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1350gat));
  NOR3_X1   g802(.A1(new_n979), .A2(G190gat), .A3(new_n684), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT125), .ZN(new_n1005));
  OAI21_X1  g804(.A(G190gat), .B1(new_n982), .B2(new_n684), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G1351gat));
  NAND2_X1  g808(.A1(new_n495), .A2(new_n978), .ZN(new_n1010));
  INV_X1    g809(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n966), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g811(.A(G197gat), .B1(new_n1012), .B2(new_n592), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n923), .A2(new_n576), .A3(new_n590), .A4(new_n1011), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(G1352gat));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n960), .A2(new_n847), .A3(new_n1011), .ZN(new_n1017));
  NOR3_X1   g816(.A1(new_n1017), .A2(G204gat), .A3(new_n707), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1016), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OR2_X1    g822(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1024), .A2(KEYINPUT62), .A3(new_n1020), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n966), .A2(new_n706), .A3(new_n1011), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1026), .A2(G204gat), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1023), .A2(new_n1025), .A3(new_n1027), .ZN(G1353gat));
  OR3_X1    g827(.A1(new_n1017), .A2(G211gat), .A3(new_n744), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n966), .A2(new_n649), .A3(new_n1011), .ZN(new_n1030));
  AND3_X1   g829(.A1(new_n1030), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1031));
  AOI21_X1  g830(.A(KEYINPUT63), .B1(new_n1030), .B2(G211gat), .ZN(new_n1032));
  OAI21_X1  g831(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(G1354gat));
  INV_X1    g832(.A(G218gat), .ZN(new_n1034));
  NOR3_X1   g833(.A1(new_n1012), .A2(new_n1034), .A3(new_n684), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1034), .B1(new_n1017), .B2(new_n684), .ZN(new_n1036));
  XNOR2_X1  g835(.A(new_n1036), .B(KEYINPUT127), .ZN(new_n1037));
  NOR2_X1   g836(.A1(new_n1035), .A2(new_n1037), .ZN(G1355gat));
endmodule


