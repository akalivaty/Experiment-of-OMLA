//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n215));
  AND3_X1   g0015(.A1(new_n214), .A2(G50), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT67), .B(G238), .Z(new_n220));
  AND2_X1   g0020(.A1(KEYINPUT66), .A2(G68), .ZN(new_n221));
  NOR2_X1   g0021(.A1(KEYINPUT66), .A2(G68), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT5), .B(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G274), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n253), .B1(new_n250), .B2(new_n248), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n254), .B1(G270), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G264), .A3(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(G257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G303), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n258), .B(new_n260), .C1(new_n261), .C2(new_n257), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n253), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n256), .A2(G179), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n207), .A2(G13), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n208), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n217), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT75), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT75), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(new_n267), .B2(new_n269), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n271), .A2(G116), .A3(new_n273), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G283), .ZN(new_n278));
  INV_X1    g0078(.A(G97), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n278), .B(new_n208), .C1(G33), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G116), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G20), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n269), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT20), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n277), .B(new_n285), .C1(new_n266), .C2(new_n282), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n265), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n256), .B2(new_n263), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT92), .B1(new_n289), .B2(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT21), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI211_X1 g0092(.A(KEYINPUT92), .B(KEYINPUT21), .C1(new_n289), .C2(new_n286), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n256), .A2(G190), .A3(new_n263), .ZN(new_n294));
  INV_X1    g0094(.A(G200), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n256), .B2(new_n263), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n294), .A2(new_n296), .A3(new_n286), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n292), .A2(new_n293), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n253), .A2(new_n252), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  AOI21_X1  g0102(.A(G1), .B1(new_n302), .B2(new_n249), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n253), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G226), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n257), .A2(G222), .A3(new_n259), .ZN(new_n306));
  INV_X1    g0106(.A(G77), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n257), .A2(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(G223), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n306), .B1(new_n307), .B2(new_n257), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT68), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n253), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n301), .B(new_n305), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT9), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT69), .ZN(new_n318));
  INV_X1    g0118(.A(G58), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT8), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n208), .A2(G33), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G20), .A2(G33), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n269), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n269), .B1(new_n207), .B2(G20), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G50), .ZN(new_n332));
  INV_X1    g0132(.A(G13), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G1), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G20), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n332), .B1(G50), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n317), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n330), .A2(new_n336), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT9), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n316), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n315), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g0143(.A(new_n343), .B(KEYINPUT10), .Z(new_n344));
  AOI21_X1  g0144(.A(new_n338), .B1(new_n315), .B2(new_n288), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G179), .B2(new_n315), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n322), .A2(new_n335), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n322), .B2(new_n331), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT3), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT7), .B1(new_n353), .B2(new_n208), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  AOI211_X1 g0155(.A(new_n355), .B(G20), .C1(new_n350), .C2(new_n352), .ZN(new_n356));
  OAI21_X1  g0156(.A(G68), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n355), .B1(new_n257), .B2(G20), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n351), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT7), .B(new_n208), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(KEYINPUT80), .A3(G68), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G58), .B1(new_n221), .B2(new_n222), .ZN(new_n367));
  INV_X1    g0167(.A(new_n201), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n208), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  INV_X1    g0170(.A(G159), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n371), .A2(G20), .A3(G33), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT81), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT80), .B1(new_n364), .B2(G68), .ZN(new_n375));
  INV_X1    g0175(.A(G68), .ZN(new_n376));
  AOI211_X1 g0176(.A(new_n358), .B(new_n376), .C1(new_n360), .C2(new_n363), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT81), .B(new_n373), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n269), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n369), .A2(new_n372), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n223), .B1(new_n360), .B2(new_n363), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT82), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI211_X1 g0184(.A(KEYINPUT82), .B(new_n223), .C1(new_n360), .C2(new_n363), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n370), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT83), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT83), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n370), .C1(new_n384), .C2(new_n385), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n349), .B1(new_n380), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT84), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n373), .B1(new_n375), .B2(new_n377), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT81), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n329), .B1(new_n395), .B2(new_n378), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n387), .A3(new_n389), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT84), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(new_n349), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  INV_X1    g0200(.A(G226), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n257), .A2(new_n259), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n400), .B1(new_n308), .B2(new_n401), .C1(new_n309), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n253), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n304), .A2(G232), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT85), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n304), .A2(KEYINPUT85), .A3(G232), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n300), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G179), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(G169), .B2(new_n410), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n392), .A2(new_n399), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n392), .A2(new_n399), .A3(new_n417), .A4(new_n414), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n410), .A2(new_n341), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n295), .B1(new_n404), .B2(new_n409), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n349), .B(new_n421), .C1(new_n380), .C2(new_n390), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n349), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n416), .A2(new_n418), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n223), .A2(G20), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n307), .B2(new_n323), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n326), .A2(G50), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n429), .B(new_n433), .C1(new_n307), .C2(new_n323), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n269), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT11), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(KEYINPUT11), .A3(new_n269), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT78), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT78), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n442), .A3(new_n439), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n207), .A2(G20), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n271), .A2(G68), .A3(new_n273), .A4(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n223), .A2(KEYINPUT12), .A3(G20), .A4(new_n334), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT12), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n335), .B2(G68), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  XOR2_X1   g0249(.A(new_n449), .B(KEYINPUT79), .Z(new_n450));
  NAND3_X1  g0250(.A1(new_n441), .A2(new_n443), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n257), .A2(G232), .A3(G1698), .ZN(new_n452));
  OAI221_X1 g0252(.A(new_n452), .B1(new_n274), .B2(new_n279), .C1(new_n402), .C2(new_n401), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n453), .A2(new_n253), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n300), .A2(KEYINPUT76), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n300), .A2(KEYINPUT76), .B1(new_n304), .B2(G238), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT13), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n253), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT13), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n455), .A4(new_n456), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT14), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(G169), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n458), .A2(G179), .A3(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n462), .B2(G169), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n451), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n449), .B(KEYINPUT79), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n440), .B2(KEYINPUT78), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n458), .A2(G190), .A3(new_n461), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n462), .A2(G200), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n443), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT72), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n321), .B(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(new_n326), .B1(G20), .B2(G77), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n477), .A2(KEYINPUT73), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT15), .B(G87), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n479), .A2(KEYINPUT74), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(KEYINPUT74), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n323), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n477), .B2(KEYINPUT73), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n329), .B1(new_n478), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n271), .A2(G77), .A3(new_n273), .A4(new_n444), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G77), .B2(new_n335), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n257), .A2(G232), .A3(new_n259), .ZN(new_n489));
  XOR2_X1   g0289(.A(KEYINPUT70), .B(G107), .Z(new_n490));
  OAI221_X1 g0290(.A(new_n489), .B1(new_n490), .B2(new_n257), .C1(new_n308), .C2(new_n220), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n253), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n300), .B1(G244), .B2(new_n304), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n288), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G179), .B2(new_n494), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT71), .ZN(new_n499));
  INV_X1    g0299(.A(new_n494), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n295), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(G190), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n485), .A2(new_n487), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n499), .A3(G190), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  NOR4_X1   g0307(.A1(new_n347), .A2(new_n428), .A3(new_n474), .A4(new_n507), .ZN(new_n508));
  OR2_X1    g0308(.A1(G238), .A2(G1698), .ZN(new_n509));
  INV_X1    g0309(.A(G244), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G1698), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n257), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT88), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n513), .B1(new_n512), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n253), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n253), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(G250), .C1(G1), .C2(new_n249), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n253), .A2(new_n252), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n250), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n295), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n257), .A2(new_n208), .A3(G68), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT19), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n323), .B2(new_n279), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G87), .A2(G97), .ZN(new_n529));
  NAND3_X1  g0329(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n490), .A2(new_n529), .B1(new_n208), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n269), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n482), .A2(new_n267), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n270), .A2(G87), .A3(new_n276), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT90), .B1(new_n524), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT90), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n512), .A2(new_n514), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT88), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n522), .B1(new_n542), .B2(new_n253), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n537), .B(new_n538), .C1(new_n543), .C2(new_n295), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(KEYINPUT91), .A3(G190), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT91), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n517), .A2(new_n523), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n341), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n536), .A2(new_n544), .A3(new_n545), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n270), .A2(new_n276), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n532), .B(new_n533), .C1(new_n482), .C2(new_n550), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n551), .A2(KEYINPUT89), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(KEYINPUT89), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n543), .A2(new_n288), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n547), .A2(new_n411), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n552), .B(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n402), .B2(new_n510), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n559), .A2(new_n278), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n253), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n520), .A2(new_n250), .A3(new_n248), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n251), .A2(new_n518), .A3(G257), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n288), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n562), .B2(new_n253), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n411), .ZN(new_n571));
  XNOR2_X1  g0371(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n572));
  INV_X1    g0372(.A(G107), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g0375(.A(G97), .B(G107), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(G20), .C1(new_n572), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n326), .A2(G77), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n490), .B1(new_n360), .B2(new_n363), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n579), .B1(KEYINPUT87), .B2(new_n580), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n580), .A2(KEYINPUT87), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n329), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n267), .A2(new_n279), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n550), .B2(new_n279), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n569), .B(new_n571), .C1(new_n583), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n257), .A2(G257), .A3(G1698), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n257), .A2(G250), .A3(new_n259), .ZN(new_n588));
  INV_X1    g0388(.A(G294), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n587), .B(new_n588), .C1(new_n274), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n253), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n255), .A2(G264), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n564), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n288), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n590), .A2(new_n253), .B1(new_n255), .B2(G264), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n411), .A3(new_n564), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n257), .A2(new_n208), .A3(G87), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT22), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT22), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n257), .A2(new_n600), .A3(new_n208), .A4(G87), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n573), .A2(G20), .ZN(new_n604));
  OAI22_X1  g0404(.A1(KEYINPUT23), .A2(new_n604), .B1(new_n323), .B2(new_n281), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n490), .A2(G20), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(KEYINPUT23), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n603), .B1(new_n602), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n269), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n334), .A2(G20), .A3(new_n573), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT25), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT93), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n612), .A2(KEYINPUT93), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n573), .B2(new_n550), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n611), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n597), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n580), .A2(KEYINPUT87), .ZN(new_n623));
  INV_X1    g0423(.A(new_n579), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n582), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n585), .B1(new_n625), .B2(new_n269), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n568), .A2(G190), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n570), .A2(G200), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n593), .A2(G190), .ZN(new_n630));
  AOI21_X1  g0430(.A(G200), .B1(new_n595), .B2(new_n564), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n611), .B(new_n620), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n586), .A2(new_n622), .A3(new_n629), .A4(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n298), .A2(new_n508), .A3(new_n557), .A4(new_n633), .ZN(G372));
  INV_X1    g0434(.A(new_n346), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n391), .A2(new_n414), .ZN(new_n636));
  XNOR2_X1  g0436(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n636), .B(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n468), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n504), .A2(new_n496), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n473), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(new_n426), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n635), .B1(new_n643), .B2(new_n344), .ZN(new_n644));
  INV_X1    g0444(.A(new_n508), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n571), .B1(G169), .B2(new_n570), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n626), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n549), .A2(new_n647), .A3(new_n556), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(KEYINPUT26), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n650));
  INV_X1    g0450(.A(new_n524), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n543), .A2(G190), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n538), .A2(KEYINPUT94), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT94), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n535), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n651), .B(new_n652), .C1(new_n653), .C2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n647), .A2(new_n656), .A3(new_n650), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n650), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT95), .B1(new_n649), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n656), .A2(new_n650), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(new_n647), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n648), .A2(KEYINPUT26), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT95), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n650), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n290), .A2(new_n291), .ZN(new_n666));
  INV_X1    g0466(.A(new_n293), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n622), .A4(new_n287), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n629), .A2(new_n586), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n660), .A4(new_n632), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n659), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n644), .B1(new_n645), .B2(new_n672), .ZN(G369));
  OR3_X1    g0473(.A1(new_n266), .A2(KEYINPUT27), .A3(G20), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT27), .B1(new_n266), .B2(G20), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n286), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n298), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n292), .A2(new_n293), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g0482(.A(KEYINPUT97), .B(G330), .Z(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n621), .A2(new_n678), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n622), .A2(new_n686), .A3(new_n632), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n597), .A2(new_n621), .A3(new_n678), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n678), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n292), .B2(new_n293), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n622), .A2(new_n632), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n622), .A2(new_n678), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n690), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n211), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n490), .A2(new_n281), .A3(new_n529), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n699), .A2(new_n207), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n216), .B2(new_n699), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  INV_X1    g0503(.A(new_n650), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n670), .B(new_n705), .C1(KEYINPUT26), .C2(new_n648), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n691), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n672), .A2(new_n678), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(KEYINPUT29), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n543), .A2(new_n570), .A3(new_n595), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT30), .B1(new_n712), .B2(new_n264), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n517), .A2(new_n595), .A3(new_n523), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n265), .A3(new_n715), .A4(new_n570), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(G179), .B1(new_n256), .B2(new_n263), .ZN(new_n718));
  AND4_X1   g0518(.A1(new_n547), .A2(new_n568), .A3(new_n718), .A4(new_n593), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT98), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n691), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n719), .B1(new_n713), .B2(new_n716), .ZN(new_n726));
  INV_X1    g0526(.A(new_n724), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT98), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n633), .A2(new_n557), .A3(new_n298), .A4(new_n691), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n723), .B1(new_n726), .B2(new_n691), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n683), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT99), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(KEYINPUT99), .A3(new_n683), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n711), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n703), .B1(new_n739), .B2(G1), .ZN(G364));
  NOR2_X1   g0540(.A1(new_n333), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n207), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n699), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n685), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n683), .B2(new_n682), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n698), .A2(new_n353), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G355), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G116), .B2(new_n211), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n698), .A2(new_n257), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n216), .B2(new_n249), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n243), .A2(new_n249), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT100), .Z(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n217), .B1(G20), .B2(new_n288), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n744), .B1(new_n754), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(G20), .A2(G179), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT101), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n341), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(G190), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G50), .A2(new_n767), .B1(new_n768), .B2(G68), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n208), .A2(G179), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n371), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(G87), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n341), .A2(G200), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n208), .B1(new_n778), .B2(new_n411), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n279), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n770), .A2(new_n341), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n573), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n777), .A2(new_n353), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n769), .A2(new_n774), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT102), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n765), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n765), .A2(new_n785), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n786), .A2(new_n778), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n786), .A2(new_n771), .A3(new_n787), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n319), .A2(new_n788), .B1(new_n789), .B2(new_n307), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n781), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n772), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n257), .B(new_n792), .C1(G329), .C2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n768), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n767), .A2(G326), .ZN(new_n797));
  INV_X1    g0597(.A(new_n779), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G294), .B1(new_n776), .B2(G303), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n794), .A2(new_n796), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n789), .B1(new_n788), .B2(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n784), .A2(new_n790), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT103), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n760), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n804), .B2(new_n805), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n763), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n682), .B2(new_n758), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n746), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  INV_X1    g0612(.A(new_n744), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n488), .A2(KEYINPUT105), .A3(new_n497), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT105), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n504), .B2(new_n496), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n506), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n671), .A2(new_n691), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n488), .A2(new_n678), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n814), .A2(new_n823), .A3(new_n817), .A4(new_n506), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n498), .B2(new_n691), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n710), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n813), .B1(new_n826), .B2(new_n738), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(KEYINPUT106), .B1(new_n738), .B2(new_n826), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(KEYINPUT106), .B2(new_n827), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n807), .A2(new_n756), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n744), .B1(G77), .B2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n257), .B(new_n780), .C1(G311), .C2(new_n793), .ZN(new_n832));
  INV_X1    g0632(.A(new_n781), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n776), .A2(G107), .B1(new_n833), .B2(G87), .ZN(new_n834));
  INV_X1    g0634(.A(new_n768), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n832), .B(new_n834), .C1(new_n791), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G303), .B2(new_n767), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n281), .B2(new_n789), .C1(new_n589), .C2(new_n788), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G137), .A2(new_n767), .B1(new_n768), .B2(G150), .ZN(new_n839));
  INV_X1    g0639(.A(G143), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n840), .B2(new_n788), .C1(new_n371), .C2(new_n789), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT34), .Z(new_n842));
  OAI22_X1  g0642(.A1(new_n202), .A2(new_n775), .B1(new_n781), .B2(new_n376), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT104), .Z(new_n844));
  AOI21_X1  g0644(.A(new_n353), .B1(new_n793), .B2(G132), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n844), .B(new_n845), .C1(new_n319), .C2(new_n779), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n838), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n831), .B1(new_n847), .B2(new_n760), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n825), .B2(new_n756), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n829), .A2(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n741), .A2(new_n207), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT16), .B1(new_n366), .B2(new_n381), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n349), .B1(new_n380), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n676), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n426), .B1(KEYINPUT18), .B2(new_n415), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n418), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n392), .A2(new_n399), .A3(new_n855), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n422), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n415), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n856), .A2(new_n422), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n854), .A2(new_n414), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n852), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n856), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n428), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n862), .A2(new_n865), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n451), .A2(new_n678), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n468), .A2(new_n473), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n451), .B(new_n678), .C1(new_n466), .C2(new_n467), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n825), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n726), .A2(new_n727), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n721), .A2(new_n678), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n880), .B2(new_n723), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT109), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n881), .A2(new_n882), .A3(new_n730), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n881), .B2(new_n730), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n872), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n859), .B1(new_n639), .B2(new_n427), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT108), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n859), .A2(new_n422), .A3(new_n636), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n890), .A2(new_n862), .B1(new_n891), .B2(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n415), .A2(new_n859), .A3(KEYINPUT108), .A4(new_n861), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n871), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n881), .A2(new_n882), .A3(new_n730), .ZN(new_n896));
  INV_X1    g0696(.A(new_n879), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n730), .A2(new_n897), .A3(new_n731), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT109), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n888), .B(new_n877), .C1(new_n896), .C2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n887), .A2(new_n888), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n883), .A2(new_n884), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n902), .B1(new_n645), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n899), .A2(new_n896), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n508), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n683), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n862), .A2(new_n890), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n392), .A2(new_n399), .A3(new_n855), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n636), .A2(new_n422), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(new_n893), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n639), .A2(new_n427), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n910), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AOI221_X4 g0716(.A(new_n852), .B1(new_n862), .B2(new_n865), .C1(new_n428), .C2(new_n868), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n908), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n640), .A2(new_n691), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n639), .A2(new_n855), .ZN(new_n923));
  INV_X1    g0723(.A(new_n876), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n819), .A2(new_n678), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n822), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n872), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n644), .B1(new_n711), .B2(new_n645), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n851), .B1(new_n907), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n907), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n575), .B1(new_n572), .B2(new_n576), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT35), .ZN(new_n935));
  OAI211_X1 g0735(.A(G116), .B(new_n218), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  XNOR2_X1  g0737(.A(KEYINPUT107), .B(KEYINPUT36), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n216), .A2(G77), .A3(new_n367), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(G50), .B2(new_n376), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n333), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n933), .A2(new_n939), .A3(new_n942), .ZN(G367));
  OAI21_X1  g0743(.A(new_n669), .B1(new_n626), .B2(new_n691), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n647), .A2(new_n678), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n694), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT42), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n944), .A2(new_n622), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n678), .B1(new_n952), .B2(new_n586), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n950), .B2(KEYINPUT42), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n653), .A2(new_n655), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n660), .B1(new_n955), .B2(new_n691), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n955), .A2(new_n650), .A3(new_n691), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n951), .A2(new_n954), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n959), .B(new_n960), .Z(new_n961));
  NOR2_X1   g0761(.A1(new_n690), .A2(new_n947), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n696), .A2(new_n946), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT45), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n696), .A2(new_n946), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT44), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n965), .A2(new_n690), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n690), .B1(new_n965), .B2(new_n967), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n684), .A2(KEYINPUT111), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n692), .A2(new_n687), .A3(new_n688), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT110), .Z(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n973), .A3(new_n948), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n684), .A2(KEYINPUT111), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n739), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n739), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n699), .B(KEYINPUT41), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n963), .B1(new_n980), .B2(new_n743), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n761), .B1(new_n482), .B2(new_n211), .C1(new_n239), .C2(new_n751), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n813), .B1(new_n982), .B2(KEYINPUT112), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(KEYINPUT112), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n779), .A2(new_n376), .ZN(new_n985));
  INV_X1    g0785(.A(G137), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n257), .B1(new_n772), .B2(new_n986), .C1(new_n307), .C2(new_n781), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(G58), .C2(new_n776), .ZN(new_n988));
  INV_X1    g0788(.A(new_n767), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n988), .B1(new_n840), .B2(new_n989), .C1(new_n371), .C2(new_n835), .ZN(new_n990));
  INV_X1    g0790(.A(G150), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n202), .A2(new_n789), .B1(new_n788), .B2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G294), .A2(new_n768), .B1(new_n767), .B2(G311), .ZN(new_n993));
  INV_X1    g0793(.A(G317), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n353), .B1(new_n772), .B2(new_n994), .C1(new_n779), .C2(new_n490), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G97), .B2(new_n833), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n776), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT46), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n775), .B2(new_n281), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n993), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n791), .A2(new_n789), .B1(new_n788), .B2(new_n261), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n990), .A2(new_n992), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT47), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n984), .B1(new_n1003), .B2(new_n760), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n758), .B2(new_n958), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n981), .A2(new_n1005), .ZN(G387));
  AOI22_X1  g0806(.A1(new_n747), .A2(new_n700), .B1(new_n573), .B2(new_n698), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n476), .A2(new_n202), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n249), .B1(new_n376), .B2(new_n307), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1009), .A2(new_n700), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n750), .B1(new_n236), .B2(new_n249), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1007), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n761), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n744), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n689), .A2(new_n758), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n257), .B1(new_n793), .B2(G326), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n779), .A2(new_n791), .B1(new_n775), .B2(new_n589), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G311), .A2(new_n768), .B1(new_n767), .B2(G322), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n261), .B2(new_n789), .C1(new_n994), .C2(new_n788), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT48), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n1021), .B2(new_n1020), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT49), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1017), .B1(new_n281), .B2(new_n781), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G159), .A2(new_n767), .B1(new_n768), .B2(new_n322), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n257), .B1(new_n772), .B2(new_n991), .C1(new_n279), .C2(new_n781), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G77), .B2(new_n776), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(new_n482), .C2(new_n779), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n202), .A2(new_n788), .B1(new_n789), .B2(new_n376), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1025), .A2(new_n1026), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1015), .B(new_n1016), .C1(new_n1032), .C2(new_n760), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n976), .B2(new_n743), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n739), .A2(new_n976), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n699), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n739), .A2(new_n976), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(G393));
  NAND2_X1  g0838(.A1(new_n977), .A2(new_n699), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n970), .B1(new_n739), .B2(new_n976), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n1039), .A2(KEYINPUT114), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT114), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n970), .A2(new_n743), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n761), .B1(new_n279), .B2(new_n211), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n751), .A2(new_n246), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n744), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n353), .B1(new_n833), .B2(G87), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n775), .A2(new_n223), .B1(new_n772), .B2(new_n840), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT113), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1048), .B1(new_n307), .B2(new_n779), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n835), .A2(new_n202), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n1050), .C2(new_n1049), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n476), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n789), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n371), .A2(new_n788), .B1(new_n989), .B2(new_n991), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT51), .Z(new_n1057));
  OAI22_X1  g0857(.A1(new_n801), .A2(new_n788), .B1(new_n989), .B2(new_n994), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT52), .Z(new_n1059));
  OAI22_X1  g0859(.A1(new_n779), .A2(new_n281), .B1(new_n775), .B2(new_n791), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n353), .B1(new_n772), .B2(new_n802), .C1(new_n573), .C2(new_n781), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(G303), .C2(new_n768), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n589), .B2(new_n789), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1055), .A2(new_n1057), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1047), .B1(new_n1064), .B2(new_n760), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n946), .B2(new_n758), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1043), .A2(new_n1044), .A3(new_n1066), .ZN(G390));
  OAI211_X1 g0867(.A(G330), .B(new_n825), .C1(new_n883), .C2(new_n884), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n924), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n732), .A2(KEYINPUT99), .A3(new_n683), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT99), .B1(new_n732), .B2(new_n683), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n878), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n926), .B1(new_n707), .B2(new_n820), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1069), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT115), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1073), .B1(new_n737), .B2(new_n878), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(KEYINPUT115), .A3(new_n1069), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n822), .A2(new_n926), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n905), .A2(G330), .A3(new_n878), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n825), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n735), .B2(new_n736), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n1083), .B2(new_n876), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1077), .A2(new_n1079), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n508), .A2(G330), .A3(new_n905), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n644), .B(new_n1086), .C1(new_n711), .C2(new_n645), .ZN(new_n1087));
  OAI21_X1  g0887(.A(KEYINPUT116), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n918), .A2(new_n921), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n920), .B1(new_n1080), .B2(new_n876), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n919), .B1(new_n1074), .B2(new_n924), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n916), .A2(new_n917), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1072), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1081), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1090), .B1(new_n918), .B2(new_n921), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1088), .A2(new_n1096), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1084), .A2(new_n1080), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT115), .B1(new_n1078), .B2(new_n1069), .ZN(new_n1103));
  AND4_X1   g0903(.A1(KEYINPUT115), .A2(new_n1069), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1087), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1081), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1072), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1098), .A2(new_n1099), .A3(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1107), .B(KEYINPUT116), .C1(new_n1108), .C2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1101), .A2(new_n1111), .A3(new_n699), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1096), .A2(new_n1100), .A3(new_n743), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1089), .A2(new_n755), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n744), .B1(new_n322), .B2(new_n830), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n353), .B1(new_n772), .B2(new_n589), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n779), .A2(new_n307), .B1(new_n781), .B2(new_n376), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(G87), .C2(new_n776), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n791), .B2(new_n989), .C1(new_n490), .C2(new_n835), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n279), .A2(new_n789), .B1(new_n788), .B2(new_n281), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n257), .B1(new_n781), .B2(new_n202), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT117), .Z(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  INV_X1    g0923(.A(G132), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1122), .B1(new_n789), .B2(new_n1123), .C1(new_n1124), .C2(new_n788), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n775), .A2(new_n991), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n768), .A2(G137), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n767), .A2(G128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n798), .A2(G159), .B1(new_n793), .B2(G125), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1119), .A2(new_n1120), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1115), .B1(new_n1132), .B2(new_n760), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1114), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1113), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1112), .A2(new_n1136), .ZN(G378));
  AND2_X1   g0937(.A1(new_n922), .A2(new_n928), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n900), .B1(new_n916), .B2(new_n917), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n885), .B1(new_n867), .B2(new_n871), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(G330), .C1(KEYINPUT40), .C2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n338), .A2(new_n676), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n347), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n347), .A2(new_n1142), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1141), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n887), .A2(new_n888), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1152), .A2(new_n1153), .A3(G330), .A4(new_n1139), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1138), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1151), .A2(new_n1154), .B1(new_n922), .B2(new_n928), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT57), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1096), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1158), .A2(new_n1106), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n699), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT120), .B1(new_n922), .B2(new_n928), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1161), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1154), .B2(new_n1151), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1158), .A2(new_n1106), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT57), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1150), .A2(new_n755), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n744), .B1(G50), .B2(new_n830), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n768), .A2(G132), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n798), .A2(G150), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n775), .A2(new_n1123), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(G128), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1174), .A2(new_n788), .B1(new_n789), .B2(new_n986), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G125), .C2(new_n767), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1179));
  OR2_X1    g0979(.A1(KEYINPUT118), .A2(G124), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(KEYINPUT118), .A2(G124), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n793), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n274), .A3(new_n302), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G159), .B2(new_n833), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1178), .A2(new_n1179), .A3(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n573), .A2(new_n788), .B1(new_n789), .B2(new_n482), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n353), .A2(new_n302), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1187), .B(new_n985), .C1(G283), .C2(new_n793), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n781), .A2(new_n319), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G77), .B2(new_n776), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(new_n279), .C2(new_n835), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1186), .B(new_n1191), .C1(G116), .C2(new_n767), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT58), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1192), .A2(KEYINPUT58), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1187), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1185), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1169), .B1(new_n1196), .B2(new_n760), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1168), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT119), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1164), .B2(new_n743), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1167), .A2(new_n1200), .ZN(G375));
  OAI211_X1 g1001(.A(new_n1102), .B(new_n1087), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1107), .A2(new_n979), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n924), .A2(new_n755), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n744), .B1(G68), .B2(new_n830), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n257), .B1(new_n772), .B2(new_n1174), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n779), .A2(new_n202), .B1(new_n775), .B2(new_n371), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G58), .C2(new_n833), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n1124), .B2(new_n989), .C1(new_n835), .C2(new_n1123), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n986), .A2(new_n788), .B1(new_n789), .B2(new_n991), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G116), .A2(new_n768), .B1(new_n767), .B2(G294), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n781), .A2(new_n307), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n353), .B1(new_n772), .B2(new_n261), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G97), .C2(new_n776), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1211), .B(new_n1214), .C1(new_n482), .C2(new_n779), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n791), .A2(new_n788), .B1(new_n789), .B2(new_n490), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1209), .A2(new_n1210), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1205), .B1(new_n1217), .B2(new_n760), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1105), .A2(new_n743), .B1(new_n1204), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1203), .A2(new_n1219), .ZN(G381));
  NOR3_X1   g1020(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT121), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1222), .A2(G390), .A3(G387), .A4(G381), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT122), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n699), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n1088), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1135), .B1(new_n1227), .B2(new_n1111), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1167), .A2(new_n1228), .A3(new_n1200), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1224), .A2(new_n1229), .ZN(G407));
  OAI211_X1 g1030(.A(G407), .B(G213), .C1(G343), .C2(new_n1229), .ZN(G409));
  NAND2_X1  g1031(.A1(new_n677), .A2(G213), .ZN(new_n1232));
  INV_X1    g1032(.A(G384), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1107), .A2(new_n699), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT60), .B1(new_n1202), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1202), .A2(new_n1235), .A3(KEYINPUT60), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1234), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1219), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1233), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1238), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(new_n1236), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G384), .B(new_n1219), .C1(new_n1243), .C2(new_n1234), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1200), .C1(new_n1160), .C2(new_n1166), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1198), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1153), .B1(new_n901), .B2(G330), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1141), .A2(new_n1150), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n929), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1138), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1247), .B1(new_n1252), .B2(new_n743), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1161), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1248), .A2(new_n1249), .B1(new_n1138), .B2(KEYINPUT120), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1165), .A2(new_n979), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(KEYINPUT123), .A3(new_n1228), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1246), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT123), .B1(new_n1257), .B2(new_n1228), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1232), .B(new_n1245), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1232), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n677), .A2(G213), .A3(G2897), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1241), .A2(new_n1244), .A3(new_n1264), .A4(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1241), .A2(new_n1244), .A3(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1265), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1264), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1263), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1257), .A2(new_n1228), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT123), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1246), .A3(new_n1258), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1232), .A4(new_n1245), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1262), .A2(new_n1272), .A3(new_n1273), .A4(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(KEYINPUT127), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1271), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1282), .A2(new_n1262), .A3(new_n1283), .A4(new_n1279), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(G393), .B(new_n811), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G390), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(G390), .A2(new_n1285), .ZN(new_n1288));
  OAI21_X1  g1088(.A(G387), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  OR2_X1    g1089(.A1(G390), .A2(new_n1285), .ZN(new_n1290));
  INV_X1    g1090(.A(G387), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1286), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1281), .A2(new_n1284), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1289), .A2(new_n1273), .A3(new_n1292), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(KEYINPUT126), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1261), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1261), .A2(new_n1297), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1296), .A2(new_n1272), .A3(new_n1298), .A4(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1294), .A2(new_n1300), .ZN(G405));
  NAND2_X1  g1101(.A1(G375), .A2(G378), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1229), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(new_n1245), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1293), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1304), .B(new_n1305), .ZN(G402));
endmodule


