//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT80), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT67), .B(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(KEYINPUT23), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OR3_X1    g015(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n207), .B(new_n210), .C1(new_n216), .C2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n223));
  OR2_X1    g022(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n225));
  AOI21_X1  g024(.A(G190gat), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n216), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n213), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n230), .A2(KEYINPUT69), .A3(new_n214), .A4(new_n215), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(KEYINPUT23), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n227), .A2(new_n231), .A3(new_n234), .A4(new_n210), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n222), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT27), .B(G183gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(KEYINPUT28), .A3(new_n213), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n224), .A2(KEYINPUT27), .A3(new_n225), .ZN(new_n241));
  NOR2_X1   g040(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n244), .B2(new_n213), .ZN(new_n245));
  AOI211_X1 g044(.A(KEYINPUT70), .B(G190gat), .C1(new_n241), .C2(new_n243), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n239), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n233), .A2(KEYINPUT26), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n206), .A2(new_n208), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n233), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n204), .B(new_n236), .C1(new_n249), .C2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n228), .A2(new_n229), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n242), .B1(new_n256), .B2(KEYINPUT27), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT70), .B1(new_n257), .B2(G190gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(new_n240), .A3(new_n213), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n248), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n254), .B1(new_n260), .B2(new_n238), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n222), .A2(new_n235), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT78), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n255), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n267), .B(new_n264), .C1(new_n261), .C2(new_n262), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G197gat), .B(G204gat), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT76), .B(G218gat), .ZN(new_n272));
  INV_X1    g071(.A(G211gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n271), .B1(new_n274), .B2(KEYINPUT22), .ZN(new_n275));
  XOR2_X1   g074(.A(G211gat), .B(G218gat), .Z(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n276), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(new_n271), .C1(new_n274), .C2(KEYINPUT22), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT77), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT77), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(new_n275), .B2(new_n276), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n203), .B1(new_n269), .B2(new_n284), .ZN(new_n285));
  AOI211_X1 g084(.A(KEYINPUT80), .B(new_n283), .C1(new_n266), .C2(new_n268), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n255), .A2(new_n263), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(new_n265), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n283), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n202), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n284), .B(new_n288), .C1(new_n289), .C2(new_n291), .ZN(new_n295));
  NOR4_X1   g094(.A1(new_n285), .A2(new_n286), .A3(new_n295), .A4(KEYINPUT81), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT37), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298));
  INV_X1    g097(.A(G64gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G92gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n269), .A2(new_n284), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT80), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT37), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n269), .A2(new_n203), .A3(new_n284), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n293), .A4(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n297), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT38), .ZN(new_n309));
  INV_X1    g108(.A(new_n302), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n310), .A2(KEYINPUT38), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n305), .B1(new_n292), .B2(new_n284), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n269), .A2(new_n283), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT1), .B1(new_n318), .B2(new_n319), .ZN(new_n321));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT72), .A4(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G113gat), .ZN(new_n326));
  INV_X1    g125(.A(G113gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G120gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n328), .A3(new_n319), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n322), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n318), .A2(new_n319), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n324), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n318), .A2(KEYINPUT1), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n335), .A2(new_n322), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G141gat), .B(G148gat), .Z(new_n342));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(KEYINPUT82), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n347), .A3(new_n340), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n342), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n340), .A2(KEYINPUT2), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT83), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n345), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n334), .A3(new_n336), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(KEYINPUT3), .ZN(new_n358));
  XOR2_X1   g157(.A(KEYINPUT84), .B(KEYINPUT3), .Z(new_n359));
  OAI211_X1 g158(.A(new_n337), .B(new_n358), .C1(new_n352), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(KEYINPUT5), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n354), .A2(new_n357), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n362), .ZN(new_n365));
  AND4_X1   g164(.A1(new_n357), .A2(new_n354), .A3(new_n360), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n355), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n353), .B1(new_n336), .B2(new_n334), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT5), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n364), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT0), .B(G57gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(G85gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n375), .B(new_n364), .C1(new_n366), .C2(new_n370), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n371), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n287), .A2(new_n293), .A3(new_n310), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n307), .A2(KEYINPUT90), .A3(new_n314), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n317), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT91), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n384), .A2(new_n383), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n388), .A2(KEYINPUT91), .A3(new_n382), .A4(new_n317), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n309), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n267), .B1(new_n280), .B2(new_n282), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n353), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n280), .ZN(new_n394));
  INV_X1    g193(.A(new_n282), .ZN(new_n395));
  INV_X1    g194(.A(new_n290), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n352), .B2(new_n359), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G228gat), .ZN(new_n399));
  INV_X1    g198(.A(G233gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n393), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n283), .A2(new_n397), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n290), .B1(new_n277), .B2(new_n279), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n352), .B1(new_n405), .B2(new_n359), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(G22gat), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  INV_X1    g210(.A(G50gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT86), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n413), .B(new_n415), .ZN(new_n416));
  OR3_X1    g215(.A1(new_n393), .A2(new_n398), .A3(new_n402), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n407), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n410), .A2(new_n416), .B1(new_n420), .B2(new_n408), .ZN(new_n421));
  AND4_X1   g220(.A1(KEYINPUT87), .A2(new_n420), .A3(new_n408), .A4(new_n416), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n302), .B1(new_n294), .B2(new_n296), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(KEYINPUT30), .A3(new_n383), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n383), .A2(KEYINPUT30), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n354), .A2(new_n357), .A3(new_n360), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n362), .ZN(new_n431));
  OR3_X1    g230(.A1(new_n367), .A2(new_n368), .A3(new_n362), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n431), .A2(KEYINPUT39), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n375), .B1(new_n431), .B2(KEYINPUT39), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n377), .B1(new_n435), .B2(KEYINPUT40), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n436), .B1(KEYINPUT40), .B2(new_n435), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n428), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n390), .A2(new_n424), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT36), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n440), .A2(KEYINPUT36), .ZN(new_n442));
  XNOR2_X1  g241(.A(G15gat), .B(G43gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G71gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(G99gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n446), .B(KEYINPUT64), .Z(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n260), .A2(new_n238), .ZN(new_n449));
  INV_X1    g248(.A(new_n254), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n338), .B1(new_n451), .B2(new_n236), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n261), .A2(new_n262), .A3(new_n337), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n445), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n451), .A2(new_n338), .A3(new_n236), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n337), .B1(new_n261), .B2(new_n262), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n447), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT32), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT73), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT73), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n454), .A2(new_n462), .A3(KEYINPUT32), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n456), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n454), .B(KEYINPUT32), .C1(new_n455), .C2(new_n445), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT74), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT74), .B1(new_n464), .B2(new_n465), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n453), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n447), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n468), .A2(new_n446), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(new_n469), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n466), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  AND4_X1   g272(.A1(KEYINPUT74), .A2(new_n472), .A3(new_n464), .A4(new_n465), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n441), .B(new_n442), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n467), .A2(new_n472), .ZN(new_n476));
  INV_X1    g275(.A(new_n466), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n474), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n440), .A3(KEYINPUT36), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n380), .A2(new_n381), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n304), .A2(new_n293), .A3(new_n306), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n287), .A2(new_n202), .A3(new_n293), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n310), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n487));
  INV_X1    g286(.A(new_n383), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n482), .B1(new_n489), .B2(new_n427), .ZN(new_n490));
  XOR2_X1   g289(.A(new_n423), .B(KEYINPUT88), .Z(new_n491));
  AOI21_X1  g290(.A(new_n481), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n423), .B1(new_n478), .B2(new_n479), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(new_n482), .C1(new_n489), .C2(new_n427), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n382), .B1(new_n426), .B2(new_n428), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n493), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n439), .A2(new_n492), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G71gat), .A2(G78gat), .ZN(new_n500));
  OR2_X1    g299(.A1(G71gat), .A2(G78gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT9), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n299), .A2(G57gat), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n504), .A2(KEYINPUT99), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(KEYINPUT99), .ZN(new_n506));
  INV_X1    g305(.A(G57gat), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n505), .B(new_n506), .C1(new_n507), .C2(G64gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n500), .A2(new_n502), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(G64gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(new_n504), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n511), .A2(new_n501), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n500), .B(KEYINPUT98), .Z(new_n513));
  AOI22_X1  g312(.A1(new_n503), .A2(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT21), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G1gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G1gat), .B2(new_n516), .ZN(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT100), .ZN(new_n523));
  AND2_X1   g322(.A1(G231gat), .A2(G233gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n514), .A2(KEYINPUT21), .ZN(new_n526));
  XNOR2_X1  g325(.A(G127gat), .B(G155gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n525), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n530));
  XNOR2_X1  g329(.A(G183gat), .B(G211gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G190gat), .B(G218gat), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT102), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n540));
  OR3_X1    g339(.A1(new_n540), .A2(G29gat), .A3(G36gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT93), .B(G29gat), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G43gat), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT15), .B1(new_n546), .B2(G50gat), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n546), .B2(G50gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT96), .B(G50gat), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n546), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n412), .A2(G43gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT15), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(new_n545), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n548), .B(KEYINPUT95), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT17), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(G99gat), .ZN(new_n563));
  INV_X1    g362(.A(G106gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT8), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(KEYINPUT101), .B(G92gat), .Z(new_n566));
  OAI211_X1 g365(.A(new_n562), .B(new_n565), .C1(G85gat), .C2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n560), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n559), .A2(new_n569), .ZN(new_n572));
  NAND3_X1  g371(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n539), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT41), .ZN(new_n576));
  INV_X1    g375(.A(G232gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n400), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n575), .B(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n538), .A2(KEYINPUT102), .ZN(new_n580));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n579), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n537), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT105), .Z(new_n586));
  NOR2_X1   g385(.A1(new_n569), .A2(new_n514), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT103), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT104), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n568), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n514), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n514), .A3(KEYINPUT10), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n586), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n597), .B1(new_n588), .B2(new_n593), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G148gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT106), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n325), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT107), .ZN(new_n605));
  OR3_X1    g404(.A1(new_n596), .A2(new_n598), .A3(new_n603), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(KEYINPUT107), .A3(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n521), .B1(new_n551), .B2(new_n558), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n560), .B2(new_n521), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(KEYINPUT18), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT18), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(KEYINPUT97), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n559), .B(new_n521), .Z(new_n618));
  XOR2_X1   g417(.A(new_n613), .B(KEYINPUT13), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n612), .A2(new_n614), .A3(KEYINPUT18), .A4(new_n613), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G169gat), .B(G197gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n617), .A2(new_n620), .A3(new_n621), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n610), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n499), .A2(new_n584), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n382), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  INV_X1    g437(.A(new_n636), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n489), .A2(new_n427), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n517), .A2(new_n520), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n647), .B(new_n648), .C1(new_n520), .C2(new_n642), .ZN(G1325gat));
  NAND2_X1  g448(.A1(new_n478), .A2(new_n479), .ZN(new_n650));
  AOI21_X1  g449(.A(G15gat), .B1(new_n636), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n481), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n639), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n653), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n491), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  NOR3_X1   g456(.A1(new_n499), .A2(new_n583), .A3(new_n635), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n536), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n382), .A2(new_n543), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n659), .A2(KEYINPUT45), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT45), .B1(new_n659), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n543), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n439), .A2(new_n492), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n495), .A2(new_n498), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n583), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(KEYINPUT44), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n499), .B2(new_n583), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n536), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT108), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n634), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n664), .B1(new_n680), .B2(new_n482), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT110), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n663), .A2(new_n681), .A3(KEYINPUT110), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1328gat));
  NOR3_X1   g485(.A1(new_n659), .A2(G36gat), .A3(new_n641), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT46), .ZN(new_n688));
  OAI21_X1  g487(.A(G36gat), .B1(new_n680), .B2(new_n641), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n669), .A2(new_n671), .A3(new_n481), .A4(new_n679), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G43gat), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n658), .A2(new_n546), .A3(new_n650), .A4(new_n536), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n691), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n693), .A2(new_n695), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT111), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(KEYINPUT47), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n698), .A2(new_n702), .ZN(G1330gat));
  OAI21_X1  g502(.A(new_n552), .B1(new_n680), .B2(new_n424), .ZN(new_n704));
  INV_X1    g503(.A(new_n491), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n659), .A2(new_n705), .A3(new_n552), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(KEYINPUT48), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n552), .B1(new_n680), .B2(new_n705), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(new_n706), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g509(.A1(new_n584), .A2(new_n632), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n499), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n610), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n482), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n507), .ZN(G1332gat));
  NOR2_X1   g515(.A1(new_n714), .A2(KEYINPUT112), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n713), .B2(new_n610), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n641), .ZN(new_n721));
  NOR2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  AND2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n721), .B2(new_n722), .ZN(G1333gat));
  NAND2_X1  g524(.A1(new_n610), .A2(new_n650), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n499), .A2(G71gat), .A3(new_n712), .A4(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n481), .B1(new_n717), .B2(new_n719), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(G71gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT50), .ZN(G1334gat));
  OAI21_X1  g529(.A(new_n491), .B1(new_n717), .B2(new_n719), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n537), .A2(new_n632), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n499), .A2(new_n583), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(KEYINPUT114), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n667), .A2(new_n668), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n733), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n734), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n737), .B2(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n735), .A2(KEYINPUT114), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(KEYINPUT51), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n740), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n742), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n743), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n609), .A2(G85gat), .A3(new_n482), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT116), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n741), .A2(new_n609), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n669), .A2(new_n671), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT113), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n669), .A2(new_n671), .A3(new_n754), .A4(new_n751), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n482), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(G85gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n750), .B1(new_n756), .B2(new_n757), .ZN(G1336gat));
  INV_X1    g557(.A(new_n566), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n755), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n640), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n641), .A2(new_n609), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n301), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n740), .B2(new_n744), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n763), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n746), .A2(new_n747), .A3(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n768));
  NAND3_X1  g567(.A1(new_n672), .A2(new_n640), .A3(new_n751), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n566), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n771), .ZN(G1337gat));
  AOI211_X1 g571(.A(new_n563), .B(new_n652), .C1(new_n753), .C2(new_n755), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n746), .A2(new_n650), .A3(new_n610), .A4(new_n747), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n563), .ZN(G1338gat));
  XOR2_X1   g574(.A(KEYINPUT118), .B(G106gat), .Z(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n760), .B2(new_n491), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n609), .A2(new_n424), .A3(G106gat), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n740), .B2(new_n744), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT53), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n746), .A2(new_n747), .A3(new_n779), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n672), .A2(new_n423), .A3(new_n751), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT53), .B1(new_n784), .B2(new_n776), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(G1339gat));
  NOR2_X1   g586(.A1(new_n640), .A2(new_n482), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n650), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n594), .A2(new_n595), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n597), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n594), .A2(new_n586), .A3(new_n595), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(KEYINPUT54), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n603), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n596), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n606), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n796), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n632), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n612), .A2(new_n613), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n618), .A2(new_n619), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n627), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n631), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n608), .A3(new_n607), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n668), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n801), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n797), .A2(new_n606), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n809), .A2(new_n583), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n676), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n711), .A2(new_n609), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n705), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(KEYINPUT119), .A3(new_n705), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n789), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820), .B2(new_n633), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n814), .A2(new_n493), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n788), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n327), .A3(new_n632), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(G1340gat));
  AOI21_X1  g624(.A(G120gat), .B1(new_n823), .B2(new_n610), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n820), .A2(new_n325), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(new_n610), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n823), .B2(new_n537), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n819), .A2(G127gat), .ZN(new_n830));
  INV_X1    g629(.A(new_n676), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n823), .A2(new_n833), .A3(new_n668), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n668), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n837), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT120), .B1(new_n837), .B2(G134gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(G1343gat));
  AOI21_X1  g639(.A(new_n424), .B1(new_n812), .B2(new_n813), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n788), .A2(new_n652), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(G141gat), .A3(new_n633), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(KEYINPUT58), .ZN(new_n846));
  INV_X1    g645(.A(G141gat), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n800), .B1(new_n799), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT121), .B1(new_n793), .B2(new_n796), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n798), .B(new_n632), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n668), .B1(new_n851), .B2(new_n807), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n536), .B1(new_n852), .B2(new_n811), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n705), .B1(new_n853), .B2(new_n813), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n843), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT57), .B(new_n424), .C1(new_n812), .C2(new_n813), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n856), .A2(new_n633), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n846), .B1(new_n847), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n853), .A2(new_n813), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n491), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n842), .B1(new_n862), .B2(KEYINPUT57), .ZN(new_n863));
  INV_X1    g662(.A(new_n857), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n856), .A2(KEYINPUT122), .A3(new_n857), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n632), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n845), .B1(new_n867), .B2(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n859), .B1(new_n868), .B2(new_n869), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n841), .A2(new_n855), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n855), .B2(new_n854), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(KEYINPUT59), .A3(new_n610), .A4(new_n843), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n863), .A2(new_n860), .A3(new_n864), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT122), .B1(new_n856), .B2(new_n857), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n609), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n876), .B2(KEYINPUT59), .ZN(new_n877));
  INV_X1    g676(.A(new_n844), .ZN(new_n878));
  AOI21_X1  g677(.A(G148gat), .B1(new_n878), .B2(new_n610), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n877), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n879), .ZN(G1345gat));
  AOI21_X1  g679(.A(G155gat), .B1(new_n878), .B2(new_n537), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n676), .B1(new_n874), .B2(new_n875), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(G155gat), .ZN(G1346gat));
  NOR3_X1   g682(.A1(new_n844), .A2(G162gat), .A3(new_n583), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT123), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n583), .B1(new_n874), .B2(new_n875), .ZN(new_n886));
  INV_X1    g685(.A(G162gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n641), .A2(new_n382), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n822), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT124), .Z(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n206), .A3(new_n632), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n817), .A2(new_n818), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(new_n650), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n633), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n892), .A2(new_n897), .ZN(G1348gat));
  NOR3_X1   g697(.A1(new_n896), .A2(new_n205), .A3(new_n609), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n891), .A2(new_n610), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n208), .ZN(G1349gat));
  OAI21_X1  g700(.A(new_n256), .B1(new_n896), .B2(new_n676), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n822), .A2(new_n237), .A3(new_n537), .A4(new_n889), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT60), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n668), .A3(new_n895), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G190gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT125), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(new_n912), .A3(G190gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(KEYINPUT61), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n891), .A2(new_n213), .A3(new_n668), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n910), .A2(KEYINPUT125), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n641), .A2(new_n382), .A3(new_n481), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n841), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(G197gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n632), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n872), .A2(new_n919), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(new_n632), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n924), .B2(new_n921), .ZN(G1352gat));
  INV_X1    g724(.A(G204gat), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n841), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n762), .A2(new_n652), .A3(new_n482), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT62), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT126), .Z(new_n930));
  OR2_X1    g729(.A1(new_n927), .A2(new_n928), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n872), .A2(new_n610), .A3(new_n919), .ZN(new_n932));
  OAI221_X1 g731(.A(new_n930), .B1(KEYINPUT62), .B2(new_n931), .C1(new_n926), .C2(new_n932), .ZN(G1353gat));
  NAND3_X1  g732(.A1(new_n920), .A2(new_n273), .A3(new_n537), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n872), .A2(new_n537), .A3(new_n919), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n920), .B2(new_n668), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n583), .A2(new_n272), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT127), .Z(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n923), .B2(new_n941), .ZN(G1355gat));
endmodule


