

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n551), .A2(G2104), .ZN(n883) );
  NOR2_X2 U552 ( .A1(G2104), .A2(n551), .ZN(n879) );
  INV_X1 U553 ( .A(G2105), .ZN(n551) );
  AND2_X1 U554 ( .A1(G2105), .A2(G2104), .ZN(n880) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n787) );
  NAND2_X2 U556 ( .A1(n534), .A2(n533), .ZN(n739) );
  AND2_X1 U557 ( .A1(n787), .A2(n535), .ZN(n534) );
  XNOR2_X1 U558 ( .A(n517), .B(KEYINPUT17), .ZN(n552) );
  XNOR2_X1 U559 ( .A(n739), .B(KEYINPUT95), .ZN(n723) );
  NOR2_X1 U560 ( .A1(n819), .A2(n529), .ZN(n528) );
  NAND2_X1 U561 ( .A1(n821), .A2(n828), .ZN(n529) );
  XNOR2_X1 U562 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U563 ( .A1(n524), .A2(n516), .ZN(n523) );
  NOR2_X1 U564 ( .A1(n967), .A2(KEYINPUT100), .ZN(n524) );
  NAND2_X1 U565 ( .A1(n520), .A2(n519), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n522), .A2(n521), .ZN(n519) );
  AND2_X1 U567 ( .A1(n525), .A2(n523), .ZN(n520) );
  INV_X1 U568 ( .A(KEYINPUT100), .ZN(n521) );
  NAND2_X1 U569 ( .A1(n531), .A2(n748), .ZN(n530) );
  INV_X1 U570 ( .A(n784), .ZN(n535) );
  INV_X1 U571 ( .A(KEYINPUT101), .ZN(n767) );
  NOR2_X1 U572 ( .A1(n542), .A2(n541), .ZN(n653) );
  INV_X1 U573 ( .A(KEYINPUT66), .ZN(n517) );
  NOR2_X1 U574 ( .A1(G651), .A2(n542), .ZN(n659) );
  NAND2_X1 U575 ( .A1(n527), .A2(n834), .ZN(n835) );
  NAND2_X1 U576 ( .A1(n800), .A2(n528), .ZN(n527) );
  OR2_X1 U577 ( .A1(n774), .A2(n759), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n518), .B(n760), .ZN(n762) );
  INV_X1 U579 ( .A(n770), .ZN(n522) );
  NAND2_X1 U580 ( .A1(n770), .A2(n526), .ZN(n525) );
  AND2_X1 U581 ( .A1(n967), .A2(KEYINPUT100), .ZN(n526) );
  XNOR2_X1 U582 ( .A(n530), .B(KEYINPUT32), .ZN(n757) );
  NAND2_X1 U583 ( .A1(n532), .A2(n751), .ZN(n531) );
  AND2_X1 U584 ( .A1(n750), .A2(n745), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n723), .A2(G2072), .ZN(n722) );
  INV_X1 U586 ( .A(n785), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n737), .A2(n736), .ZN(n751) );
  NOR2_X1 U588 ( .A1(n714), .A2(n955), .ZN(n719) );
  INV_X1 U589 ( .A(KEYINPUT28), .ZN(n729) );
  XNOR2_X1 U590 ( .A(n702), .B(n701), .ZN(n703) );
  INV_X1 U591 ( .A(KEYINPUT29), .ZN(n733) );
  XNOR2_X1 U592 ( .A(n734), .B(n733), .ZN(n737) );
  INV_X1 U593 ( .A(KEYINPUT64), .ZN(n760) );
  INV_X1 U594 ( .A(KEYINPUT102), .ZN(n777) );
  INV_X1 U595 ( .A(KEYINPUT13), .ZN(n591) );
  XNOR2_X1 U596 ( .A(n592), .B(n591), .ZN(n593) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n650) );
  INV_X1 U598 ( .A(G651), .ZN(n541) );
  NOR2_X1 U599 ( .A1(G543), .A2(n541), .ZN(n537) );
  XNOR2_X1 U600 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(n664) );
  NAND2_X1 U602 ( .A1(G64), .A2(n664), .ZN(n539) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n542) );
  NAND2_X1 U604 ( .A1(G52), .A2(n659), .ZN(n538) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U606 ( .A(KEYINPUT71), .B(n540), .Z(n547) );
  NAND2_X1 U607 ( .A1(G77), .A2(n653), .ZN(n544) );
  NAND2_X1 U608 ( .A1(G90), .A2(n650), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n545), .Z(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(G171) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  NAND2_X1 U615 ( .A1(G126), .A2(n879), .ZN(n549) );
  NAND2_X1 U616 ( .A1(G114), .A2(n880), .ZN(n548) );
  NAND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(KEYINPUT86), .B(n550), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n883), .A2(G102), .ZN(n555) );
  NOR2_X1 U620 ( .A1(G2105), .A2(G2104), .ZN(n553) );
  XNOR2_X2 U621 ( .A(n553), .B(n552), .ZN(n626) );
  NAND2_X1 U622 ( .A1(G138), .A2(n626), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(G164) );
  NAND2_X1 U625 ( .A1(n650), .A2(G88), .ZN(n560) );
  NAND2_X1 U626 ( .A1(G75), .A2(n653), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT83), .B(n558), .Z(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G62), .A2(n664), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G50), .A2(n659), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U632 ( .A1(n564), .A2(n563), .ZN(G166) );
  NAND2_X1 U633 ( .A1(G89), .A2(n650), .ZN(n565) );
  XOR2_X1 U634 ( .A(KEYINPUT4), .B(n565), .Z(n566) );
  XNOR2_X1 U635 ( .A(n566), .B(KEYINPUT77), .ZN(n568) );
  NAND2_X1 U636 ( .A1(G76), .A2(n653), .ZN(n567) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n569), .B(KEYINPUT5), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G63), .A2(n664), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G51), .A2(n659), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U642 ( .A(KEYINPUT6), .B(n572), .Z(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n575), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(G101), .A2(n883), .ZN(n576) );
  XNOR2_X1 U647 ( .A(n576), .B(KEYINPUT65), .ZN(n577) );
  XNOR2_X1 U648 ( .A(n577), .B(KEYINPUT23), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n626), .A2(G137), .ZN(n578) );
  XOR2_X1 U650 ( .A(KEYINPUT67), .B(n578), .Z(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n785) );
  NAND2_X1 U652 ( .A1(G125), .A2(n879), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G113), .A2(n880), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n694) );
  NOR2_X1 U655 ( .A1(n785), .A2(n694), .ZN(G160) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n583), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U658 ( .A(G223), .B(KEYINPUT74), .Z(n836) );
  NAND2_X1 U659 ( .A1(n836), .A2(G567), .ZN(n584) );
  XOR2_X1 U660 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U661 ( .A1(G56), .A2(n664), .ZN(n585) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(n585), .Z(n594) );
  NAND2_X1 U663 ( .A1(n653), .A2(G68), .ZN(n586) );
  XNOR2_X1 U664 ( .A(n586), .B(KEYINPUT76), .ZN(n590) );
  XOR2_X1 U665 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n588) );
  NAND2_X1 U666 ( .A1(G81), .A2(n650), .ZN(n587) );
  XNOR2_X1 U667 ( .A(n588), .B(n587), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n592) );
  NOR2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n659), .A2(G43), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n955) );
  INV_X1 U672 ( .A(G860), .ZN(n634) );
  OR2_X1 U673 ( .A1(n955), .A2(n634), .ZN(G153) );
  INV_X1 U674 ( .A(G171), .ZN(G301) );
  NAND2_X1 U675 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G79), .A2(n653), .ZN(n598) );
  NAND2_X1 U677 ( .A1(G66), .A2(n664), .ZN(n597) );
  NAND2_X1 U678 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U679 ( .A1(G92), .A2(n650), .ZN(n600) );
  NAND2_X1 U680 ( .A1(G54), .A2(n659), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U682 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U683 ( .A(KEYINPUT15), .B(n603), .Z(n956) );
  INV_X1 U684 ( .A(n956), .ZN(n617) );
  INV_X1 U685 ( .A(G868), .ZN(n677) );
  NAND2_X1 U686 ( .A1(n617), .A2(n677), .ZN(n604) );
  NAND2_X1 U687 ( .A1(n605), .A2(n604), .ZN(G284) );
  NAND2_X1 U688 ( .A1(G65), .A2(n664), .ZN(n607) );
  NAND2_X1 U689 ( .A1(G53), .A2(n659), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U691 ( .A(KEYINPUT72), .B(n608), .Z(n612) );
  NAND2_X1 U692 ( .A1(G78), .A2(n653), .ZN(n610) );
  NAND2_X1 U693 ( .A1(G91), .A2(n650), .ZN(n609) );
  AND2_X1 U694 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(G299) );
  NOR2_X1 U696 ( .A1(G286), .A2(n677), .ZN(n614) );
  NOR2_X1 U697 ( .A1(G868), .A2(G299), .ZN(n613) );
  NOR2_X1 U698 ( .A1(n614), .A2(n613), .ZN(G297) );
  NAND2_X1 U699 ( .A1(n634), .A2(G559), .ZN(n615) );
  NAND2_X1 U700 ( .A1(n615), .A2(n956), .ZN(n616) );
  XNOR2_X1 U701 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U702 ( .A1(n617), .A2(n677), .ZN(n618) );
  XOR2_X1 U703 ( .A(KEYINPUT78), .B(n618), .Z(n619) );
  NOR2_X1 U704 ( .A1(G559), .A2(n619), .ZN(n621) );
  NOR2_X1 U705 ( .A1(G868), .A2(n955), .ZN(n620) );
  NOR2_X1 U706 ( .A1(n621), .A2(n620), .ZN(G282) );
  XOR2_X1 U707 ( .A(G2100), .B(KEYINPUT80), .Z(n632) );
  NAND2_X1 U708 ( .A1(G123), .A2(n879), .ZN(n622) );
  XOR2_X1 U709 ( .A(KEYINPUT18), .B(n622), .Z(n623) );
  XNOR2_X1 U710 ( .A(n623), .B(KEYINPUT79), .ZN(n625) );
  NAND2_X1 U711 ( .A1(G111), .A2(n880), .ZN(n624) );
  NAND2_X1 U712 ( .A1(n625), .A2(n624), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n883), .A2(G99), .ZN(n628) );
  NAND2_X1 U714 ( .A1(G135), .A2(n626), .ZN(n627) );
  NAND2_X1 U715 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n935) );
  XNOR2_X1 U717 ( .A(n935), .B(G2096), .ZN(n631) );
  NAND2_X1 U718 ( .A1(n632), .A2(n631), .ZN(G156) );
  NAND2_X1 U719 ( .A1(G559), .A2(n956), .ZN(n633) );
  XOR2_X1 U720 ( .A(n955), .B(n633), .Z(n674) );
  NAND2_X1 U721 ( .A1(n634), .A2(n674), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G80), .A2(n653), .ZN(n636) );
  NAND2_X1 U723 ( .A1(G67), .A2(n664), .ZN(n635) );
  NAND2_X1 U724 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G93), .A2(n650), .ZN(n638) );
  NAND2_X1 U726 ( .A1(G55), .A2(n659), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U728 ( .A1(n640), .A2(n639), .ZN(n676) );
  XOR2_X1 U729 ( .A(n641), .B(n676), .Z(G145) );
  NAND2_X1 U730 ( .A1(G72), .A2(n653), .ZN(n643) );
  NAND2_X1 U731 ( .A1(G85), .A2(n650), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U733 ( .A(KEYINPUT68), .B(n644), .Z(n649) );
  NAND2_X1 U734 ( .A1(n659), .A2(G47), .ZN(n646) );
  NAND2_X1 U735 ( .A1(n664), .A2(G60), .ZN(n645) );
  NAND2_X1 U736 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U737 ( .A(KEYINPUT70), .B(n647), .Z(n648) );
  NAND2_X1 U738 ( .A1(n649), .A2(n648), .ZN(G290) );
  NAND2_X1 U739 ( .A1(G86), .A2(n650), .ZN(n652) );
  NAND2_X1 U740 ( .A1(G61), .A2(n664), .ZN(n651) );
  NAND2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U742 ( .A1(n653), .A2(G73), .ZN(n654) );
  XOR2_X1 U743 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U744 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U745 ( .A1(n659), .A2(G48), .ZN(n657) );
  NAND2_X1 U746 ( .A1(n658), .A2(n657), .ZN(G305) );
  NAND2_X1 U747 ( .A1(n659), .A2(G49), .ZN(n660) );
  XOR2_X1 U748 ( .A(KEYINPUT81), .B(n660), .Z(n662) );
  NAND2_X1 U749 ( .A1(G651), .A2(G74), .ZN(n661) );
  NAND2_X1 U750 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U751 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U752 ( .A(n665), .B(KEYINPUT82), .ZN(n667) );
  NAND2_X1 U753 ( .A1(G87), .A2(n542), .ZN(n666) );
  NAND2_X1 U754 ( .A1(n667), .A2(n666), .ZN(G288) );
  XNOR2_X1 U755 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n668) );
  XNOR2_X1 U756 ( .A(n668), .B(n676), .ZN(n669) );
  XNOR2_X1 U757 ( .A(n669), .B(G290), .ZN(n672) );
  INV_X1 U758 ( .A(G299), .ZN(n959) );
  XNOR2_X1 U759 ( .A(G166), .B(n959), .ZN(n670) );
  XNOR2_X1 U760 ( .A(n670), .B(G305), .ZN(n671) );
  XNOR2_X1 U761 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U762 ( .A(n673), .B(G288), .ZN(n906) );
  XOR2_X1 U763 ( .A(n906), .B(n674), .Z(n675) );
  NOR2_X1 U764 ( .A1(n677), .A2(n675), .ZN(n679) );
  AND2_X1 U765 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U766 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U767 ( .A1(G2078), .A2(G2084), .ZN(n680) );
  XOR2_X1 U768 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U769 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U770 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n683), .A2(G2072), .ZN(n684) );
  XOR2_X1 U772 ( .A(KEYINPUT85), .B(n684), .Z(G158) );
  XNOR2_X1 U773 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  XNOR2_X1 U774 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U775 ( .A1(G108), .A2(G120), .ZN(n685) );
  NOR2_X1 U776 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U777 ( .A1(G69), .A2(n686), .ZN(n925) );
  NAND2_X1 U778 ( .A1(n925), .A2(G567), .ZN(n691) );
  NOR2_X1 U779 ( .A1(G220), .A2(G219), .ZN(n687) );
  XOR2_X1 U780 ( .A(KEYINPUT22), .B(n687), .Z(n688) );
  NOR2_X1 U781 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U782 ( .A1(G96), .A2(n689), .ZN(n926) );
  NAND2_X1 U783 ( .A1(n926), .A2(G2106), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n840) );
  NAND2_X1 U785 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U786 ( .A1(n840), .A2(n692), .ZN(n839) );
  NAND2_X1 U787 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U788 ( .A(G166), .ZN(G303) );
  INV_X1 U789 ( .A(G40), .ZN(n693) );
  OR2_X1 U790 ( .A1(n694), .A2(n693), .ZN(n784) );
  NAND2_X1 U791 ( .A1(n739), .A2(G8), .ZN(n696) );
  XNOR2_X2 U792 ( .A(n696), .B(KEYINPUT94), .ZN(n774) );
  NOR2_X1 U793 ( .A1(n774), .A2(G1966), .ZN(n753) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n739), .ZN(n749) );
  INV_X1 U795 ( .A(n749), .ZN(n697) );
  NAND2_X1 U796 ( .A1(G8), .A2(n697), .ZN(n698) );
  NOR2_X1 U797 ( .A1(n753), .A2(n698), .ZN(n702) );
  XOR2_X1 U798 ( .A(KEYINPUT30), .B(KEYINPUT97), .Z(n700) );
  INV_X1 U799 ( .A(KEYINPUT98), .ZN(n699) );
  NOR2_X1 U800 ( .A1(G168), .A2(n703), .ZN(n707) );
  INV_X1 U801 ( .A(G1961), .ZN(n981) );
  NAND2_X1 U802 ( .A1(n981), .A2(n739), .ZN(n705) );
  XNOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .ZN(n1008) );
  NAND2_X1 U804 ( .A1(n723), .A2(n1008), .ZN(n704) );
  NAND2_X1 U805 ( .A1(n705), .A2(n704), .ZN(n735) );
  NOR2_X1 U806 ( .A1(G171), .A2(n735), .ZN(n706) );
  NOR2_X1 U807 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U808 ( .A(n708), .B(KEYINPUT31), .Z(n750) );
  INV_X1 U809 ( .A(G1996), .ZN(n709) );
  NOR2_X1 U810 ( .A1(n739), .A2(n709), .ZN(n711) );
  XOR2_X1 U811 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n710) );
  XNOR2_X1 U812 ( .A(n711), .B(n710), .ZN(n713) );
  NAND2_X1 U813 ( .A1(n739), .A2(G1341), .ZN(n712) );
  NAND2_X1 U814 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U815 ( .A1(n719), .A2(n956), .ZN(n718) );
  NAND2_X1 U816 ( .A1(G2067), .A2(n723), .ZN(n716) );
  NAND2_X1 U817 ( .A1(G1348), .A2(n739), .ZN(n715) );
  NAND2_X1 U818 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U819 ( .A1(n718), .A2(n717), .ZN(n721) );
  OR2_X1 U820 ( .A1(n956), .A2(n719), .ZN(n720) );
  NAND2_X1 U821 ( .A1(n721), .A2(n720), .ZN(n727) );
  XNOR2_X1 U822 ( .A(n722), .B(KEYINPUT27), .ZN(n725) );
  INV_X1 U823 ( .A(G1956), .ZN(n982) );
  NOR2_X1 U824 ( .A1(n982), .A2(n723), .ZN(n724) );
  NOR2_X1 U825 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U826 ( .A1(n959), .A2(n728), .ZN(n726) );
  NAND2_X1 U827 ( .A1(n727), .A2(n726), .ZN(n732) );
  NOR2_X1 U828 ( .A1(n959), .A2(n728), .ZN(n730) );
  XNOR2_X1 U829 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U830 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U831 ( .A1(n735), .A2(G171), .ZN(n736) );
  INV_X1 U832 ( .A(G8), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n774), .A2(G1971), .ZN(n738) );
  XNOR2_X1 U834 ( .A(KEYINPUT99), .B(n738), .ZN(n742) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U836 ( .A1(G166), .A2(n740), .ZN(n741) );
  NAND2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n743) );
  OR2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U839 ( .A(n745), .ZN(n747) );
  AND2_X1 U840 ( .A1(G286), .A2(G8), .ZN(n746) );
  OR2_X1 U841 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U842 ( .A1(G8), .A2(n749), .ZN(n755) );
  AND2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n770) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U848 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U849 ( .A1(n763), .A2(n758), .ZN(n967) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n962) );
  INV_X1 U851 ( .A(n962), .ZN(n759) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n766) );
  INV_X1 U854 ( .A(n774), .ZN(n780) );
  NAND2_X1 U855 ( .A1(n780), .A2(n763), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n768) );
  XNOR2_X1 U858 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n974) );
  NAND2_X1 U860 ( .A1(n769), .A2(n974), .ZN(n776) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U862 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n770), .A2(n772), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(n777), .ZN(n783) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XNOR2_X1 U868 ( .A(n779), .B(KEYINPUT24), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n800) );
  OR2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U873 ( .A(KEYINPUT87), .B(n788), .Z(n832) );
  XNOR2_X1 U874 ( .A(KEYINPUT37), .B(G2067), .ZN(n830) );
  NAND2_X1 U875 ( .A1(G140), .A2(n626), .ZN(n789) );
  XNOR2_X1 U876 ( .A(n789), .B(KEYINPUT88), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G104), .A2(n883), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U879 ( .A(KEYINPUT34), .B(n792), .ZN(n798) );
  NAND2_X1 U880 ( .A1(n879), .A2(G128), .ZN(n793) );
  XOR2_X1 U881 ( .A(KEYINPUT89), .B(n793), .Z(n795) );
  NAND2_X1 U882 ( .A1(n880), .A2(G116), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U884 ( .A(KEYINPUT35), .B(n796), .Z(n797) );
  NOR2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U886 ( .A(KEYINPUT36), .B(n799), .ZN(n895) );
  NOR2_X1 U887 ( .A1(n830), .A2(n895), .ZN(n948) );
  NAND2_X1 U888 ( .A1(n832), .A2(n948), .ZN(n828) );
  NAND2_X1 U889 ( .A1(n880), .A2(G117), .ZN(n807) );
  NAND2_X1 U890 ( .A1(G129), .A2(n879), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G141), .A2(n626), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n883), .A2(G105), .ZN(n803) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(n803), .Z(n804) );
  NOR2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U897 ( .A(KEYINPUT91), .B(n808), .Z(n900) );
  NAND2_X1 U898 ( .A1(G1996), .A2(n900), .ZN(n809) );
  XOR2_X1 U899 ( .A(KEYINPUT92), .B(n809), .Z(n818) );
  NAND2_X1 U900 ( .A1(n879), .A2(G119), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n810), .B(KEYINPUT90), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G131), .A2(n626), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n816) );
  NAND2_X1 U904 ( .A1(G107), .A2(n880), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G95), .A2(n883), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n894) );
  AND2_X1 U908 ( .A1(G1991), .A2(n894), .ZN(n817) );
  NOR2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n932) );
  INV_X1 U910 ( .A(n832), .ZN(n820) );
  NOR2_X1 U911 ( .A1(n932), .A2(n820), .ZN(n824) );
  XOR2_X1 U912 ( .A(KEYINPUT93), .B(n824), .Z(n819) );
  XOR2_X1 U913 ( .A(G1986), .B(G290), .Z(n963) );
  OR2_X1 U914 ( .A1(n963), .A2(n820), .ZN(n821) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n900), .ZN(n937) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n894), .ZN(n940) );
  NOR2_X1 U918 ( .A1(n822), .A2(n940), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U920 ( .A1(n937), .A2(n825), .ZN(n826) );
  XOR2_X1 U921 ( .A(KEYINPUT39), .B(n826), .Z(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(KEYINPUT103), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n830), .A2(n895), .ZN(n945) );
  NAND2_X1 U925 ( .A1(n831), .A2(n945), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(KEYINPUT40), .B(n835), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U930 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U933 ( .A(n840), .ZN(G319) );
  XNOR2_X1 U934 ( .A(G1996), .B(KEYINPUT41), .ZN(n850) );
  XOR2_X1 U935 ( .A(G1956), .B(G1966), .Z(n842) );
  XNOR2_X1 U936 ( .A(G1991), .B(G1981), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U938 ( .A(G1961), .B(G1971), .Z(n844) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1976), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U941 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT108), .B(G2474), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U944 ( .A(n850), .B(n849), .ZN(G229) );
  XNOR2_X1 U945 ( .A(G2072), .B(G2090), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n851), .B(KEYINPUT105), .ZN(n861) );
  XOR2_X1 U947 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n853) );
  XNOR2_X1 U948 ( .A(G2678), .B(G2100), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U950 ( .A(G2096), .B(G2084), .Z(n855) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2078), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U953 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U954 ( .A(KEYINPUT43), .B(KEYINPUT42), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U957 ( .A1(G124), .A2(n879), .ZN(n862) );
  XNOR2_X1 U958 ( .A(n862), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U959 ( .A1(G112), .A2(n880), .ZN(n863) );
  XOR2_X1 U960 ( .A(KEYINPUT109), .B(n863), .Z(n864) );
  NAND2_X1 U961 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U962 ( .A1(n883), .A2(G100), .ZN(n867) );
  NAND2_X1 U963 ( .A1(G136), .A2(n626), .ZN(n866) );
  NAND2_X1 U964 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U965 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U966 ( .A(n935), .B(G162), .Z(n878) );
  NAND2_X1 U967 ( .A1(n883), .A2(G103), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G139), .A2(n626), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G127), .A2(n879), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G115), .A2(n880), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n928) );
  XNOR2_X1 U975 ( .A(G164), .B(n928), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n902) );
  NAND2_X1 U977 ( .A1(G130), .A2(n879), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G118), .A2(n880), .ZN(n881) );
  NAND2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n889) );
  NAND2_X1 U980 ( .A1(n883), .A2(G106), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G142), .A2(n626), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U983 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  XNOR2_X1 U984 ( .A(KEYINPUT110), .B(n887), .ZN(n888) );
  NOR2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n893) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n891) );
  XNOR2_X1 U987 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U990 ( .A(n895), .B(n894), .Z(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U992 ( .A(G160), .B(n898), .Z(n899) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U994 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U995 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n955), .B(KEYINPUT113), .ZN(n905) );
  XNOR2_X1 U997 ( .A(G171), .B(n956), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n908) );
  XNOR2_X1 U999 ( .A(G286), .B(n906), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1002 ( .A(G2443), .B(G2451), .Z(n911) );
  XNOR2_X1 U1003 ( .A(G2446), .B(G2454), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1005 ( .A(n912), .B(G2427), .Z(n914) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(n914), .B(n913), .ZN(n918) );
  XOR2_X1 U1008 ( .A(G2435), .B(KEYINPUT104), .Z(n916) );
  XNOR2_X1 U1009 ( .A(G2430), .B(G2438), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1011 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1012 ( .A1(G14), .A2(n919), .ZN(n927) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n927), .ZN(n922) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(G225) );
  XOR2_X1 U1019 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1021 ( .A(G120), .ZN(G236) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  INV_X1 U1023 ( .A(G96), .ZN(G221) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(G325) );
  INV_X1 U1026 ( .A(G325), .ZN(G261) );
  INV_X1 U1027 ( .A(n927), .ZN(G401) );
  XOR2_X1 U1028 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n931), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n944) );
  XOR2_X1 U1033 ( .A(G2084), .B(G160), .Z(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(n938), .B(KEYINPUT51), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(n949), .ZN(n951) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n952), .A2(G29), .ZN(n953) );
  XOR2_X1 U1047 ( .A(KEYINPUT115), .B(n953), .Z(n1037) );
  INV_X1 U1048 ( .A(G16), .ZN(n1005) );
  XOR2_X1 U1049 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n954) );
  XNOR2_X1 U1050 ( .A(n1005), .B(n954), .ZN(n980) );
  XNOR2_X1 U1051 ( .A(n955), .B(G1341), .ZN(n972) );
  XNOR2_X1 U1052 ( .A(G1348), .B(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(G1971), .A2(G303), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n969) );
  XNOR2_X1 U1055 ( .A(n959), .B(G1956), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G171), .B(G1961), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(KEYINPUT123), .B(n970), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT124), .B(n973), .ZN(n978) );
  XNOR2_X1 U1065 ( .A(G1966), .B(G168), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT57), .B(n976), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n1007) );
  XNOR2_X1 U1070 ( .A(G5), .B(n981), .ZN(n994) );
  XNOR2_X1 U1071 ( .A(G20), .B(n982), .ZN(n986) );
  XNOR2_X1 U1072 ( .A(G1981), .B(G6), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G19), .B(G1341), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n989) );
  XOR2_X1 U1076 ( .A(KEYINPUT59), .B(G1348), .Z(n987) );
  XNOR2_X1 U1077 ( .A(G4), .B(n987), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1079 ( .A(KEYINPUT60), .B(n990), .Z(n992) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G21), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n1002) );
  XNOR2_X1 U1083 ( .A(G1986), .B(G24), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(G22), .B(G1971), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G1976), .B(KEYINPUT125), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(G23), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(KEYINPUT58), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT61), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1035) );
  XNOR2_X1 U1094 ( .A(G27), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(G2067), .B(G26), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G1996), .B(G32), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(G33), .B(G2072), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT118), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(G28), .ZN(n1019) );
  XOR2_X1 U1103 ( .A(G25), .B(G1991), .Z(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT117), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(KEYINPUT53), .B(n1020), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(n1021), .B(KEYINPUT119), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(G2090), .B(G35), .Z(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT116), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(KEYINPUT120), .B(n1025), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(G34), .B(G2084), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(KEYINPUT54), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1115 ( .A(KEYINPUT55), .B(n1029), .ZN(n1031) );
  INV_X1 U1116 ( .A(G29), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(G11), .ZN(n1033) );
  XOR2_X1 U1119 ( .A(KEYINPUT121), .B(n1033), .Z(n1034) );
  NOR2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1122 ( .A(n1038), .B(KEYINPUT126), .ZN(n1039) );
  XNOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1039), .ZN(G150) );
  INV_X1 U1124 ( .A(G150), .ZN(G311) );
endmodule

