

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746;

  XNOR2_X2 U370 ( .A(n543), .B(KEYINPUT107), .ZN(n538) );
  NOR2_X2 U371 ( .A1(n535), .A2(n545), .ZN(n642) );
  XNOR2_X2 U372 ( .A(n540), .B(n444), .ZN(n746) );
  AND2_X2 U373 ( .A1(n669), .A2(n670), .ZN(n374) );
  INV_X1 U374 ( .A(n588), .ZN(n687) );
  XNOR2_X1 U375 ( .A(n599), .B(KEYINPUT40), .ZN(n744) );
  NAND2_X1 U376 ( .A1(n383), .A2(n382), .ZN(n573) );
  AND2_X1 U377 ( .A1(n385), .A2(n384), .ZN(n383) );
  XNOR2_X1 U378 ( .A(n503), .B(n502), .ZN(n628) );
  XNOR2_X1 U379 ( .A(n420), .B(KEYINPUT66), .ZN(n482) );
  XNOR2_X1 U380 ( .A(n730), .B(n483), .ZN(n359) );
  AND2_X1 U381 ( .A1(n701), .A2(n667), .ZN(n470) );
  XNOR2_X1 U382 ( .A(n423), .B(KEYINPUT83), .ZN(n616) );
  XNOR2_X1 U383 ( .A(n448), .B(n463), .ZN(n375) );
  INV_X1 U384 ( .A(KEYINPUT3), .ZN(n461) );
  XNOR2_X1 U385 ( .A(n430), .B(n402), .ZN(n625) );
  INV_X1 U386 ( .A(KEYINPUT1), .ZN(n402) );
  NOR2_X1 U387 ( .A1(n566), .A2(n403), .ZN(n604) );
  AND2_X1 U388 ( .A1(n413), .A2(n584), .ZN(n412) );
  NAND2_X1 U389 ( .A1(n548), .A2(KEYINPUT34), .ZN(n413) );
  NAND2_X1 U390 ( .A1(n374), .A2(G478), .ZN(n429) );
  NAND2_X1 U391 ( .A1(n374), .A2(G475), .ZN(n409) );
  NOR2_X1 U392 ( .A1(n746), .A2(KEYINPUT84), .ZN(n442) );
  NOR2_X1 U393 ( .A1(n441), .A2(n741), .ZN(n541) );
  NAND2_X1 U394 ( .A1(n380), .A2(n379), .ZN(n441) );
  AND2_X1 U395 ( .A1(n443), .A2(n381), .ZN(n380) );
  NAND2_X1 U396 ( .A1(n368), .A2(n442), .ZN(n379) );
  NAND2_X1 U397 ( .A1(n639), .A2(n386), .ZN(n384) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n525) );
  XNOR2_X1 U399 ( .A(n516), .B(n417), .ZN(n730) );
  XNOR2_X1 U400 ( .A(n482), .B(n418), .ZN(n417) );
  XNOR2_X1 U401 ( .A(n419), .B(G131), .ZN(n418) );
  INV_X1 U402 ( .A(G137), .ZN(n419) );
  XNOR2_X1 U403 ( .A(n364), .B(KEYINPUT78), .ZN(n363) );
  INV_X1 U404 ( .A(G101), .ZN(n364) );
  INV_X1 U405 ( .A(KEYINPUT2), .ZN(n666) );
  NOR2_X1 U406 ( .A1(G237), .A2(G902), .ZN(n456) );
  NOR2_X1 U407 ( .A1(n716), .A2(G902), .ZN(n503) );
  XNOR2_X1 U408 ( .A(n437), .B(n492), .ZN(n436) );
  XNOR2_X1 U409 ( .A(n490), .B(KEYINPUT95), .ZN(n437) );
  INV_X1 U410 ( .A(KEYINPUT24), .ZN(n490) );
  XOR2_X1 U411 ( .A(G128), .B(G119), .Z(n449) );
  XNOR2_X1 U412 ( .A(n491), .B(n434), .ZN(n731) );
  XNOR2_X1 U413 ( .A(G140), .B(KEYINPUT10), .ZN(n434) );
  XNOR2_X1 U414 ( .A(n445), .B(n720), .ZN(n701) );
  XNOR2_X1 U415 ( .A(n482), .B(n469), .ZN(n446) );
  XNOR2_X1 U416 ( .A(n597), .B(n353), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n610), .B(n373), .ZN(n372) );
  INV_X1 U418 ( .A(KEYINPUT112), .ZN(n373) );
  XNOR2_X1 U419 ( .A(n508), .B(n507), .ZN(n653) );
  NAND2_X1 U420 ( .A1(n627), .A2(n628), .ZN(n624) );
  XNOR2_X1 U421 ( .A(n352), .B(n404), .ZN(n430) );
  INV_X1 U422 ( .A(G469), .ZN(n404) );
  XOR2_X1 U423 ( .A(KEYINPUT6), .B(n631), .Z(n572) );
  XNOR2_X1 U424 ( .A(n514), .B(n398), .ZN(n714) );
  XNOR2_X1 U425 ( .A(n515), .B(n399), .ZN(n398) );
  XNOR2_X1 U426 ( .A(G107), .B(G116), .ZN(n512) );
  AND2_X1 U427 ( .A1(n392), .A2(n668), .ZN(n669) );
  INV_X1 U428 ( .A(KEYINPUT84), .ZN(n440) );
  INV_X1 U429 ( .A(KEYINPUT85), .ZN(n386) );
  XNOR2_X1 U430 ( .A(n422), .B(G128), .ZN(n481) );
  INV_X1 U431 ( .A(G143), .ZN(n422) );
  XNOR2_X1 U432 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n458) );
  XNOR2_X1 U433 ( .A(n481), .B(n421), .ZN(n516) );
  INV_X1 U434 ( .A(G134), .ZN(n421) );
  XNOR2_X1 U435 ( .A(G122), .B(KEYINPUT11), .ZN(n521) );
  XNOR2_X1 U436 ( .A(G143), .B(G131), .ZN(n519) );
  XOR2_X1 U437 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n527) );
  XNOR2_X1 U438 ( .A(n554), .B(KEYINPUT45), .ZN(n556) );
  INV_X1 U439 ( .A(KEYINPUT4), .ZN(n420) );
  XNOR2_X1 U440 ( .A(n389), .B(KEYINPUT68), .ZN(n570) );
  XNOR2_X1 U441 ( .A(n365), .B(KEYINPUT74), .ZN(n546) );
  NOR2_X1 U442 ( .A1(n625), .A2(n624), .ZN(n365) );
  NOR2_X1 U443 ( .A1(n624), .A2(n432), .ZN(n431) );
  NAND2_X1 U444 ( .A1(n476), .A2(n475), .ZN(n367) );
  XNOR2_X1 U445 ( .A(n359), .B(n450), .ZN(n672) );
  XNOR2_X1 U446 ( .A(n504), .B(KEYINPUT5), .ZN(n400) );
  INV_X1 U447 ( .A(n556), .ZN(n725) );
  INV_X1 U448 ( .A(n516), .ZN(n399) );
  XNOR2_X1 U449 ( .A(n396), .B(n511), .ZN(n513) );
  XNOR2_X1 U450 ( .A(n510), .B(n397), .ZN(n396) );
  INV_X1 U451 ( .A(KEYINPUT7), .ZN(n397) );
  XOR2_X1 U452 ( .A(G902), .B(KEYINPUT15), .Z(n457) );
  XNOR2_X1 U453 ( .A(n732), .B(n356), .ZN(n665) );
  XNOR2_X1 U454 ( .A(n361), .B(n359), .ZN(n705) );
  XNOR2_X1 U455 ( .A(n480), .B(n362), .ZN(n361) );
  XNOR2_X1 U456 ( .A(n479), .B(n363), .ZN(n362) );
  INV_X1 U457 ( .A(G953), .ZN(n663) );
  XOR2_X1 U458 ( .A(KEYINPUT90), .B(n473), .Z(n639) );
  BUF_X1 U459 ( .A(n613), .Z(n395) );
  XNOR2_X1 U460 ( .A(n518), .B(n517), .ZN(n544) );
  XNOR2_X1 U461 ( .A(n466), .B(n375), .ZN(n720) );
  XNOR2_X1 U462 ( .A(KEYINPUT16), .B(G122), .ZN(n465) );
  XNOR2_X1 U463 ( .A(n435), .B(n731), .ZN(n498) );
  XNOR2_X1 U464 ( .A(n489), .B(n436), .ZN(n435) );
  XNOR2_X1 U465 ( .A(KEYINPUT42), .B(n605), .ZN(n742) );
  NAND2_X1 U466 ( .A1(n360), .A2(n690), .ZN(n599) );
  XNOR2_X1 U467 ( .A(n370), .B(n369), .ZN(n575) );
  INV_X1 U468 ( .A(KEYINPUT36), .ZN(n369) );
  XNOR2_X1 U469 ( .A(n366), .B(n534), .ZN(n741) );
  NAND2_X1 U470 ( .A1(n347), .A2(n410), .ZN(n366) );
  OR2_X1 U471 ( .A1(n653), .A2(n414), .ZN(n410) );
  INV_X1 U472 ( .A(KEYINPUT32), .ZN(n444) );
  AND2_X1 U473 ( .A1(n349), .A2(n574), .ZN(n390) );
  INV_X1 U474 ( .A(n624), .ZN(n401) );
  NAND2_X1 U475 ( .A1(n427), .A2(n407), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n429), .B(n428), .ZN(n427) );
  INV_X1 U477 ( .A(n714), .ZN(n428) );
  INV_X1 U478 ( .A(KEYINPUT60), .ZN(n405) );
  NAND2_X1 U479 ( .A1(n408), .A2(n407), .ZN(n406) );
  XNOR2_X1 U480 ( .A(n409), .B(n354), .ZN(n408) );
  AND2_X1 U481 ( .A1(n411), .A2(n412), .ZN(n347) );
  NAND2_X1 U482 ( .A1(n642), .A2(n627), .ZN(n348) );
  NOR2_X1 U483 ( .A1(n572), .A2(n628), .ZN(n349) );
  OR2_X1 U484 ( .A1(n639), .A2(n386), .ZN(n350) );
  AND2_X1 U485 ( .A1(n382), .A2(n474), .ZN(n351) );
  NOR2_X1 U486 ( .A1(n705), .A2(G902), .ZN(n352) );
  XOR2_X1 U487 ( .A(KEYINPUT39), .B(KEYINPUT72), .Z(n353) );
  INV_X1 U488 ( .A(KEYINPUT34), .ZN(n416) );
  XOR2_X1 U489 ( .A(n713), .B(n712), .Z(n354) );
  XOR2_X1 U490 ( .A(n672), .B(n671), .Z(n355) );
  AND2_X1 U491 ( .A1(n666), .A2(KEYINPUT76), .ZN(n356) );
  XOR2_X1 U492 ( .A(KEYINPUT86), .B(n674), .Z(n357) );
  XOR2_X1 U493 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n358) );
  INV_X1 U494 ( .A(G146), .ZN(n483) );
  INV_X1 U495 ( .A(n718), .ZN(n407) );
  AND2_X1 U496 ( .A1(n360), .A2(n692), .ZN(n698) );
  AND2_X1 U497 ( .A1(n546), .A2(n572), .ZN(n508) );
  NAND2_X1 U498 ( .A1(n367), .A2(n477), .ZN(n438) );
  NAND2_X1 U499 ( .A1(n604), .A2(n367), .ZN(n588) );
  INV_X1 U500 ( .A(n368), .ZN(n683) );
  NAND2_X1 U501 ( .A1(n538), .A2(n377), .ZN(n368) );
  NAND2_X1 U502 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U503 ( .A(n573), .ZN(n371) );
  NAND2_X1 U504 ( .A1(n571), .A2(n572), .ZN(n610) );
  NAND2_X1 U505 ( .A1(n374), .A2(G210), .ZN(n703) );
  NAND2_X1 U506 ( .A1(n374), .A2(G472), .ZN(n673) );
  NAND2_X1 U507 ( .A1(n374), .A2(G469), .ZN(n708) );
  NAND2_X1 U508 ( .A1(n374), .A2(G217), .ZN(n715) );
  XNOR2_X1 U509 ( .A(n375), .B(n400), .ZN(n450) );
  NAND2_X1 U510 ( .A1(n538), .A2(n376), .ZN(n381) );
  AND2_X1 U511 ( .A1(n439), .A2(n562), .ZN(n376) );
  NOR2_X1 U512 ( .A1(n631), .A2(n378), .ZN(n377) );
  INV_X1 U513 ( .A(n562), .ZN(n378) );
  NAND2_X1 U514 ( .A1(n351), .A2(n383), .ZN(n475) );
  OR2_X1 U515 ( .A1(n613), .A2(n350), .ZN(n382) );
  NAND2_X1 U516 ( .A1(n613), .A2(n386), .ZN(n385) );
  XNOR2_X1 U517 ( .A(n406), .B(n405), .ZN(G60) );
  XNOR2_X1 U518 ( .A(n387), .B(n357), .ZN(G57) );
  NAND2_X1 U519 ( .A1(n394), .A2(n407), .ZN(n387) );
  NAND2_X1 U520 ( .A1(n415), .A2(n416), .ZN(n414) );
  NAND2_X1 U521 ( .A1(n388), .A2(KEYINPUT47), .ZN(n569) );
  NAND2_X1 U522 ( .A1(n687), .A2(n567), .ZN(n388) );
  NAND2_X1 U523 ( .A1(n563), .A2(n627), .ZN(n389) );
  NAND2_X1 U524 ( .A1(n573), .A2(KEYINPUT19), .ZN(n476) );
  NAND2_X1 U525 ( .A1(n539), .A2(n390), .ZN(n540) );
  XOR2_X1 U526 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n494) );
  XNOR2_X1 U527 ( .A(n391), .B(n425), .ZN(n424) );
  NAND2_X1 U528 ( .A1(n608), .A2(n609), .ZN(n391) );
  NAND2_X1 U529 ( .A1(n509), .A2(G221), .ZN(n496) );
  XNOR2_X1 U530 ( .A(n495), .B(KEYINPUT81), .ZN(n509) );
  NAND2_X2 U531 ( .A1(n616), .A2(n615), .ZN(n732) );
  XNOR2_X1 U532 ( .A(n438), .B(KEYINPUT0), .ZN(n536) );
  NAND2_X1 U533 ( .A1(n725), .A2(n666), .ZN(n392) );
  XNOR2_X1 U534 ( .A(n470), .B(n471), .ZN(n613) );
  XNOR2_X1 U535 ( .A(n393), .B(n358), .ZN(G51) );
  NAND2_X1 U536 ( .A1(n704), .A2(n407), .ZN(n393) );
  XNOR2_X1 U537 ( .A(n673), .B(n355), .ZN(n394) );
  NAND2_X1 U538 ( .A1(n744), .A2(n742), .ZN(n607) );
  NAND2_X1 U539 ( .A1(n631), .A2(n576), .ZN(n578) );
  XNOR2_X2 U540 ( .A(n505), .B(n506), .ZN(n631) );
  AND2_X1 U541 ( .A1(n430), .A2(n401), .ZN(n433) );
  INV_X1 U542 ( .A(n430), .ZN(n403) );
  NAND2_X1 U543 ( .A1(n653), .A2(KEYINPUT34), .ZN(n411) );
  INV_X1 U544 ( .A(n548), .ZN(n415) );
  XNOR2_X1 U545 ( .A(n426), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U546 ( .A(n460), .B(n459), .ZN(n448) );
  NAND2_X1 U547 ( .A1(n424), .A2(n699), .ZN(n423) );
  INV_X1 U548 ( .A(KEYINPUT48), .ZN(n425) );
  NAND2_X1 U549 ( .A1(n431), .A2(n430), .ZN(n580) );
  INV_X1 U550 ( .A(n579), .ZN(n432) );
  NAND2_X1 U551 ( .A1(n415), .A2(n433), .ZN(n549) );
  NOR2_X2 U552 ( .A1(n536), .A2(n348), .ZN(n537) );
  NOR2_X1 U553 ( .A1(n631), .A2(n440), .ZN(n439) );
  NAND2_X1 U554 ( .A1(n746), .A2(KEYINPUT84), .ZN(n443) );
  XNOR2_X1 U555 ( .A(n447), .B(n446), .ZN(n445) );
  XNOR2_X1 U556 ( .A(n468), .B(n491), .ZN(n447) );
  BUF_X1 U557 ( .A(n556), .Z(n664) );
  INV_X1 U558 ( .A(n628), .ZN(n562) );
  XNOR2_X1 U559 ( .A(n481), .B(n467), .ZN(n468) );
  INV_X1 U560 ( .A(n698), .ZN(n615) );
  XNOR2_X1 U561 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U562 ( .A(n478), .B(n465), .ZN(n466) );
  NOR2_X1 U563 ( .A1(G952), .A2(n663), .ZN(n718) );
  XNOR2_X1 U564 ( .A(n662), .B(n661), .ZN(G75) );
  NAND2_X1 U565 ( .A1(G237), .A2(G234), .ZN(n451) );
  XNOR2_X1 U566 ( .A(n451), .B(KEYINPUT14), .ZN(n453) );
  NAND2_X1 U567 ( .A1(G902), .A2(n453), .ZN(n557) );
  XOR2_X1 U568 ( .A(G898), .B(KEYINPUT92), .Z(n724) );
  NAND2_X1 U569 ( .A1(G953), .A2(n724), .ZN(n719) );
  NOR2_X1 U570 ( .A1(n557), .A2(n719), .ZN(n452) );
  XNOR2_X1 U571 ( .A(KEYINPUT93), .B(n452), .ZN(n455) );
  NAND2_X1 U572 ( .A1(G952), .A2(n453), .ZN(n652) );
  NOR2_X1 U573 ( .A1(n652), .A2(G953), .ZN(n454) );
  XNOR2_X1 U574 ( .A(n454), .B(KEYINPUT91), .ZN(n560) );
  NAND2_X1 U575 ( .A1(n455), .A2(n560), .ZN(n477) );
  XNOR2_X1 U576 ( .A(n456), .B(KEYINPUT75), .ZN(n472) );
  AND2_X1 U577 ( .A1(n472), .A2(G210), .ZN(n471) );
  XNOR2_X1 U578 ( .A(KEYINPUT89), .B(n457), .ZN(n667) );
  INV_X1 U579 ( .A(n458), .ZN(n460) );
  XNOR2_X1 U580 ( .A(G119), .B(G101), .ZN(n459) );
  XNOR2_X1 U581 ( .A(G116), .B(G113), .ZN(n462) );
  XNOR2_X1 U582 ( .A(G107), .B(G110), .ZN(n464) );
  XNOR2_X1 U583 ( .A(n464), .B(G104), .ZN(n478) );
  XOR2_X1 U584 ( .A(G146), .B(G125), .Z(n491) );
  XOR2_X1 U585 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n467) );
  NAND2_X1 U586 ( .A1(G224), .A2(n663), .ZN(n469) );
  NAND2_X1 U587 ( .A1(n472), .A2(G214), .ZN(n473) );
  INV_X1 U588 ( .A(KEYINPUT19), .ZN(n474) );
  BUF_X1 U589 ( .A(n536), .Z(n548) );
  XOR2_X1 U590 ( .A(G140), .B(n478), .Z(n480) );
  NAND2_X1 U591 ( .A1(G227), .A2(n663), .ZN(n479) );
  XOR2_X1 U592 ( .A(KEYINPUT21), .B(KEYINPUT98), .Z(n486) );
  NAND2_X1 U593 ( .A1(G234), .A2(n667), .ZN(n484) );
  XNOR2_X1 U594 ( .A(KEYINPUT20), .B(n484), .ZN(n499) );
  NAND2_X1 U595 ( .A1(n499), .A2(G221), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n486), .B(n485), .ZN(n627) );
  XOR2_X1 U597 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n488) );
  XNOR2_X1 U598 ( .A(G137), .B(G110), .ZN(n487) );
  XNOR2_X1 U599 ( .A(n488), .B(n487), .ZN(n489) );
  INV_X1 U600 ( .A(KEYINPUT96), .ZN(n492) );
  NAND2_X1 U601 ( .A1(G234), .A2(n663), .ZN(n493) );
  XNOR2_X1 U602 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U603 ( .A(n496), .B(n449), .ZN(n497) );
  XNOR2_X1 U604 ( .A(n497), .B(n498), .ZN(n716) );
  XOR2_X1 U605 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n501) );
  NAND2_X1 U606 ( .A1(n499), .A2(G217), .ZN(n500) );
  XNOR2_X1 U607 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U608 ( .A(KEYINPUT99), .B(G472), .ZN(n506) );
  NAND2_X1 U609 ( .A1(n525), .A2(G210), .ZN(n504) );
  NOR2_X1 U610 ( .A1(G902), .A2(n672), .ZN(n505) );
  XOR2_X1 U611 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n507) );
  XNOR2_X1 U612 ( .A(G478), .B(KEYINPUT106), .ZN(n518) );
  NAND2_X1 U613 ( .A1(n509), .A2(G217), .ZN(n515) );
  XOR2_X1 U614 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n511) );
  XNOR2_X1 U615 ( .A(G122), .B(KEYINPUT9), .ZN(n510) );
  XNOR2_X1 U616 ( .A(n513), .B(n512), .ZN(n514) );
  NOR2_X1 U617 ( .A1(n714), .A2(G902), .ZN(n517) );
  INV_X1 U618 ( .A(n544), .ZN(n535) );
  XOR2_X1 U619 ( .A(G104), .B(G113), .Z(n520) );
  XNOR2_X1 U620 ( .A(n520), .B(n519), .ZN(n524) );
  XOR2_X1 U621 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n522) );
  XNOR2_X1 U622 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U623 ( .A(n524), .B(n523), .ZN(n529) );
  NAND2_X1 U624 ( .A1(G214), .A2(n525), .ZN(n526) );
  XNOR2_X1 U625 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U626 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U627 ( .A(n731), .B(n530), .ZN(n711) );
  NOR2_X1 U628 ( .A1(G902), .A2(n711), .ZN(n532) );
  XNOR2_X1 U629 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n531) );
  XNOR2_X1 U630 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U631 ( .A(G475), .B(n533), .Z(n545) );
  AND2_X1 U632 ( .A1(n535), .A2(n545), .ZN(n584) );
  XOR2_X1 U633 ( .A(KEYINPUT35), .B(KEYINPUT79), .Z(n534) );
  INV_X1 U634 ( .A(n642), .ZN(n600) );
  XNOR2_X1 U635 ( .A(n537), .B(KEYINPUT22), .ZN(n539) );
  NAND2_X1 U636 ( .A1(n539), .A2(n625), .ZN(n543) );
  XNOR2_X1 U637 ( .A(n625), .B(KEYINPUT87), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n541), .B(KEYINPUT44), .ZN(n553) );
  OR2_X1 U639 ( .A1(n562), .A2(n572), .ZN(n542) );
  NOR2_X1 U640 ( .A1(n543), .A2(n542), .ZN(n675) );
  NAND2_X1 U641 ( .A1(n545), .A2(n544), .ZN(n598) );
  INV_X1 U642 ( .A(n598), .ZN(n690) );
  NOR2_X1 U643 ( .A1(n545), .A2(n544), .ZN(n692) );
  NOR2_X1 U644 ( .A1(n690), .A2(n692), .ZN(n640) );
  NAND2_X1 U645 ( .A1(n631), .A2(n546), .ZN(n635) );
  NOR2_X1 U646 ( .A1(n548), .A2(n635), .ZN(n547) );
  XOR2_X1 U647 ( .A(KEYINPUT31), .B(n547), .Z(n693) );
  NOR2_X1 U648 ( .A1(n631), .A2(n549), .ZN(n678) );
  NOR2_X1 U649 ( .A1(n693), .A2(n678), .ZN(n550) );
  NOR2_X1 U650 ( .A1(n640), .A2(n550), .ZN(n551) );
  NOR2_X1 U651 ( .A1(n675), .A2(n551), .ZN(n552) );
  NAND2_X1 U652 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U653 ( .A(KEYINPUT82), .B(n664), .ZN(n555) );
  NAND2_X1 U654 ( .A1(n555), .A2(n666), .ZN(n620) );
  NAND2_X1 U655 ( .A1(KEYINPUT80), .A2(n640), .ZN(n567) );
  NOR2_X1 U656 ( .A1(G900), .A2(n557), .ZN(n558) );
  NAND2_X1 U657 ( .A1(G953), .A2(n558), .ZN(n559) );
  XNOR2_X1 U658 ( .A(n559), .B(KEYINPUT108), .ZN(n561) );
  NAND2_X1 U659 ( .A1(n561), .A2(n560), .ZN(n579) );
  AND2_X1 U660 ( .A1(n562), .A2(n579), .ZN(n563) );
  INV_X1 U661 ( .A(n570), .ZN(n564) );
  NAND2_X1 U662 ( .A1(n564), .A2(n631), .ZN(n565) );
  XNOR2_X1 U663 ( .A(n565), .B(KEYINPUT28), .ZN(n566) );
  OR2_X1 U664 ( .A1(KEYINPUT47), .A2(KEYINPUT80), .ZN(n568) );
  NAND2_X1 U665 ( .A1(n569), .A2(n568), .ZN(n587) );
  NOR2_X1 U666 ( .A1(n570), .A2(n598), .ZN(n571) );
  NAND2_X1 U667 ( .A1(n575), .A2(n574), .ZN(n695) );
  INV_X1 U668 ( .A(n639), .ZN(n576) );
  XNOR2_X1 U669 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n577) );
  XNOR2_X1 U670 ( .A(n578), .B(n577), .ZN(n582) );
  XNOR2_X1 U671 ( .A(n580), .B(KEYINPUT77), .ZN(n581) );
  NAND2_X1 U672 ( .A1(n582), .A2(n581), .ZN(n596) );
  NOR2_X1 U673 ( .A1(n395), .A2(n596), .ZN(n583) );
  XNOR2_X1 U674 ( .A(KEYINPUT110), .B(n583), .ZN(n585) );
  NAND2_X1 U675 ( .A1(n585), .A2(n584), .ZN(n686) );
  NAND2_X1 U676 ( .A1(n695), .A2(n686), .ZN(n586) );
  NOR2_X1 U677 ( .A1(n587), .A2(n586), .ZN(n594) );
  INV_X1 U678 ( .A(KEYINPUT80), .ZN(n590) );
  NOR2_X1 U679 ( .A1(n588), .A2(KEYINPUT47), .ZN(n589) );
  NOR2_X1 U680 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U681 ( .A1(n640), .A2(n591), .ZN(n592) );
  INV_X1 U682 ( .A(n592), .ZN(n593) );
  AND2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n609) );
  XNOR2_X1 U684 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n595) );
  XNOR2_X1 U685 ( .A(n395), .B(n595), .ZN(n644) );
  NOR2_X1 U686 ( .A1(n596), .A2(n644), .ZN(n597) );
  XOR2_X1 U687 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n603) );
  NOR2_X1 U688 ( .A1(n639), .A2(n600), .ZN(n646) );
  INV_X1 U689 ( .A(n644), .ZN(n601) );
  NAND2_X1 U690 ( .A1(n646), .A2(n601), .ZN(n602) );
  XNOR2_X1 U691 ( .A(n603), .B(n602), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n623), .A2(n604), .ZN(n605) );
  XOR2_X1 U693 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n606) );
  XNOR2_X1 U694 ( .A(n607), .B(n606), .ZN(n608) );
  NOR2_X1 U695 ( .A1(n639), .A2(n610), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n625), .A2(n611), .ZN(n612) );
  XNOR2_X1 U697 ( .A(n612), .B(KEYINPUT43), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n614), .A2(n395), .ZN(n699) );
  NOR2_X1 U699 ( .A1(n725), .A2(n732), .ZN(n617) );
  NOR2_X1 U700 ( .A1(n666), .A2(n617), .ZN(n618) );
  NAND2_X1 U701 ( .A1(KEYINPUT82), .A2(n618), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n666), .A2(n732), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n658) );
  INV_X1 U705 ( .A(n623), .ZN(n654) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U707 ( .A(KEYINPUT50), .B(n626), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT49), .B(n629), .Z(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n634), .B(KEYINPUT118), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U714 ( .A(KEYINPUT51), .B(n637), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n654), .A2(n638), .ZN(n649) );
  NOR2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U720 ( .A1(n647), .A2(n653), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n650), .B(KEYINPUT52), .ZN(n651) );
  NOR2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U727 ( .A1(G953), .A2(n659), .ZN(n662) );
  INV_X1 U728 ( .A(KEYINPUT53), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(KEYINPUT119), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n670) );
  INV_X1 U731 ( .A(n667), .ZN(n668) );
  XOR2_X1 U732 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n671) );
  XOR2_X1 U733 ( .A(KEYINPUT63), .B(KEYINPUT88), .Z(n674) );
  XOR2_X1 U734 ( .A(G101), .B(n675), .Z(n676) );
  XNOR2_X1 U735 ( .A(KEYINPUT114), .B(n676), .ZN(G3) );
  NAND2_X1 U736 ( .A1(n678), .A2(n690), .ZN(n677) );
  XNOR2_X1 U737 ( .A(n677), .B(G104), .ZN(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n680) );
  NAND2_X1 U739 ( .A1(n678), .A2(n692), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n680), .B(n679), .ZN(n682) );
  XOR2_X1 U741 ( .A(G107), .B(KEYINPUT27), .Z(n681) );
  XNOR2_X1 U742 ( .A(n682), .B(n681), .ZN(G9) );
  XOR2_X1 U743 ( .A(G110), .B(n683), .Z(G12) );
  XOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .Z(n685) );
  NAND2_X1 U745 ( .A1(n687), .A2(n692), .ZN(n684) );
  XNOR2_X1 U746 ( .A(n685), .B(n684), .ZN(G30) );
  XNOR2_X1 U747 ( .A(G143), .B(n686), .ZN(G45) );
  NAND2_X1 U748 ( .A1(n687), .A2(n690), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(KEYINPUT116), .ZN(n689) );
  XNOR2_X1 U750 ( .A(G146), .B(n689), .ZN(G48) );
  NAND2_X1 U751 ( .A1(n693), .A2(n690), .ZN(n691) );
  XNOR2_X1 U752 ( .A(n691), .B(G113), .ZN(G15) );
  NAND2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U754 ( .A(n694), .B(G116), .ZN(G18) );
  XNOR2_X1 U755 ( .A(KEYINPUT37), .B(KEYINPUT117), .ZN(n696) );
  XNOR2_X1 U756 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U757 ( .A(G125), .B(n697), .ZN(G27) );
  XOR2_X1 U758 ( .A(G134), .B(n698), .Z(G36) );
  XNOR2_X1 U759 ( .A(G140), .B(n699), .ZN(G42) );
  XOR2_X1 U760 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n700) );
  XNOR2_X1 U761 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U762 ( .A(n703), .B(n702), .ZN(n704) );
  XOR2_X1 U763 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n707) );
  XNOR2_X1 U764 ( .A(n705), .B(KEYINPUT121), .ZN(n706) );
  XNOR2_X1 U765 ( .A(n707), .B(n706), .ZN(n709) );
  XOR2_X1 U766 ( .A(n709), .B(n708), .Z(n710) );
  NOR2_X1 U767 ( .A1(n718), .A2(n710), .ZN(G54) );
  XNOR2_X1 U768 ( .A(KEYINPUT59), .B(KEYINPUT65), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n711), .B(KEYINPUT122), .ZN(n712) );
  XNOR2_X1 U770 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U771 ( .A1(n718), .A2(n717), .ZN(G66) );
  NAND2_X1 U772 ( .A1(n720), .A2(n719), .ZN(n729) );
  XOR2_X1 U773 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n722) );
  NAND2_X1 U774 ( .A1(G224), .A2(G953), .ZN(n721) );
  XNOR2_X1 U775 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n727) );
  NOR2_X1 U777 ( .A1(G953), .A2(n725), .ZN(n726) );
  NOR2_X1 U778 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n729), .B(n728), .ZN(G69) );
  XNOR2_X1 U780 ( .A(n730), .B(n731), .ZN(n736) );
  INV_X1 U781 ( .A(n736), .ZN(n733) );
  XNOR2_X1 U782 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U783 ( .A1(G953), .A2(n734), .ZN(n735) );
  XNOR2_X1 U784 ( .A(KEYINPUT125), .B(n735), .ZN(n740) );
  XNOR2_X1 U785 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U787 ( .A1(n738), .A2(G953), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n740), .A2(n739), .ZN(G72) );
  XOR2_X1 U789 ( .A(n741), .B(G122), .Z(G24) );
  XNOR2_X1 U790 ( .A(G137), .B(n742), .ZN(n743) );
  XNOR2_X1 U791 ( .A(n743), .B(KEYINPUT126), .ZN(G39) );
  XOR2_X1 U792 ( .A(n744), .B(G131), .Z(n745) );
  XNOR2_X1 U793 ( .A(KEYINPUT127), .B(n745), .ZN(G33) );
  XOR2_X1 U794 ( .A(n746), .B(G119), .Z(G21) );
endmodule

