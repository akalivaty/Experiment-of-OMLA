//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G50), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT65), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n211), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n203), .A2(new_n204), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n225), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT75), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  OAI211_X1 g0060(.A(KEYINPUT7), .B(new_n230), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n253), .B1(new_n262), .B2(G68), .ZN(new_n263));
  AOI211_X1 g0063(.A(KEYINPUT75), .B(new_n214), .C1(new_n256), .C2(new_n261), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT70), .A2(G58), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT70), .A2(G58), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n213), .A2(new_n215), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n202), .ZN(new_n269));
  NOR3_X1   g0069(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n230), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G159), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT76), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n212), .A2(G68), .ZN(new_n279));
  OR2_X1    g0079(.A1(KEYINPUT70), .A2(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT70), .A2(G58), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n278), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(G20), .B1(new_n282), .B2(new_n203), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT76), .ZN(new_n284));
  INV_X1    g0084(.A(new_n276), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n277), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n265), .A2(new_n287), .A3(KEYINPUT16), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n229), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n255), .A2(new_n254), .A3(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n257), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT7), .B1(new_n295), .B2(new_n230), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n283), .B(new_n285), .C1(new_n297), .C2(new_n216), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT16), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n291), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT8), .A2(G58), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n267), .A2(new_n266), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n304), .B2(KEYINPUT8), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(KEYINPUT69), .A2(G1), .ZN(new_n307));
  NAND2_X1  g0107(.A1(KEYINPUT69), .A2(G1), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n307), .A2(G13), .A3(G20), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT69), .A2(G1), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT69), .A2(G1), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n290), .B1(new_n313), .B2(G20), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n305), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n301), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT77), .ZN(new_n319));
  INV_X1    g0119(.A(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n288), .B2(new_n300), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT77), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G87), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT78), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n293), .A2(new_n294), .A3(G226), .A4(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n293), .A2(new_n294), .A3(G223), .A4(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G41), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G1), .A3(G13), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n332), .A2(G274), .ZN(new_n335));
  INV_X1    g0135(.A(G1), .ZN(new_n336));
  OR2_X1    g0136(.A1(KEYINPUT68), .A2(G41), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT68), .A2(G41), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n335), .B(new_n336), .C1(G45), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n313), .A2(G41), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n307), .A2(G45), .A3(new_n308), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(G232), .A3(new_n332), .A4(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n334), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(G169), .B2(new_n344), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n319), .A2(new_n323), .A3(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n340), .A2(new_n343), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n350), .A2(KEYINPUT79), .A3(new_n351), .A4(new_n334), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT79), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n344), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n344), .A2(G190), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n321), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n301), .A2(new_n357), .A3(new_n317), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(KEYINPUT80), .B2(KEYINPUT17), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n349), .A2(KEYINPUT18), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n216), .A2(G20), .B1(G50), .B2(new_n273), .ZN(new_n364));
  INV_X1    g0164(.A(G77), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n230), .A2(G33), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT71), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n366), .B(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n364), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT11), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n369), .A2(new_n370), .A3(new_n290), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(new_n369), .B2(new_n290), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n371), .A2(new_n372), .B1(new_n214), .B2(new_n315), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT12), .B1(new_n217), .B2(new_n309), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT74), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n309), .A2(KEYINPUT12), .A3(G68), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n295), .A2(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G226), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n295), .A2(new_n328), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G232), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n333), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT13), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n341), .A2(G238), .A3(new_n332), .A4(new_n342), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n340), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n386), .B1(new_n385), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(G200), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n391), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(G190), .A3(new_n389), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n378), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G169), .B1(new_n390), .B2(new_n391), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(G179), .A3(new_n389), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(G169), .C1(new_n390), .C2(new_n391), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n378), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n396), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n322), .B1(new_n301), .B2(new_n317), .ZN(new_n405));
  AOI211_X1 g0205(.A(KEYINPUT77), .B(new_n320), .C1(new_n288), .C2(new_n300), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n405), .A2(new_n406), .A3(new_n347), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n363), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT8), .B(G58), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n411), .A2(new_n274), .B1(new_n230), .B2(new_n365), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n366), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n290), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n314), .A2(G77), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n415), .B(new_n416), .C1(G77), .C2(new_n309), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n379), .A2(KEYINPUT72), .A3(G232), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT72), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n255), .A2(new_n328), .ZN(new_n420));
  INV_X1    g0220(.A(G232), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n381), .A2(G238), .B1(G107), .B2(new_n295), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n332), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G244), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n341), .A2(new_n332), .A3(new_n342), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n340), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n417), .B1(new_n429), .B2(G190), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n425), .B2(new_n428), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n345), .ZN(new_n433));
  INV_X1    g0233(.A(G169), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n425), .B2(new_n428), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n417), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n205), .A2(G20), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n273), .A2(G150), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n438), .B(new_n439), .C1(new_n306), .C2(new_n368), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n290), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n309), .A2(G50), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(G50), .B2(new_n314), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n381), .A2(G223), .B1(G77), .B2(new_n295), .ZN(new_n446));
  INV_X1    g0246(.A(G222), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(new_n420), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n333), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n341), .A2(G226), .A3(new_n332), .A4(new_n342), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n340), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n445), .B1(new_n434), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(new_n345), .A3(new_n451), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n452), .A2(new_n351), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(G200), .B2(new_n452), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n444), .A2(KEYINPUT9), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT9), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n441), .A2(new_n459), .A3(new_n443), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT10), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n457), .B2(new_n461), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n437), .B(new_n455), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n465), .A2(KEYINPUT73), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(KEYINPUT73), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n410), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n255), .A2(G257), .A3(new_n328), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n295), .A2(G303), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n255), .A2(G1698), .ZN(new_n472));
  INV_X1    g0272(.A(G264), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n333), .ZN(new_n475));
  INV_X1    g0275(.A(G41), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT5), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n307), .A2(new_n477), .A3(G45), .A4(new_n308), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT5), .B1(new_n337), .B2(new_n338), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n335), .ZN(new_n481));
  OAI211_X1 g0281(.A(G270), .B(new_n332), .C1(new_n478), .C2(new_n479), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G200), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n309), .A2(G116), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n307), .A2(G33), .A3(new_n308), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n309), .A2(new_n291), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n487), .B2(G116), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT81), .B(G97), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n230), .B(new_n489), .C1(new_n490), .C2(G33), .ZN(new_n491));
  INV_X1    g0291(.A(G116), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n289), .A2(new_n229), .B1(G20), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(KEYINPUT20), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT20), .B1(new_n491), .B2(new_n493), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n488), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT86), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n484), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n484), .B2(new_n498), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n483), .A2(new_n351), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n497), .A2(new_n483), .A3(G169), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n497), .A2(new_n483), .A3(KEYINPUT21), .A4(G169), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G179), .A3(new_n497), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n309), .A2(G97), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n487), .B2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT6), .B1(new_n490), .B2(G107), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G97), .A2(G107), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n209), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n516), .B1(new_n515), .B2(new_n519), .ZN(new_n522));
  OAI21_X1  g0322(.A(G20), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n262), .A2(G107), .B1(G77), .B2(new_n273), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n514), .B1(new_n525), .B2(new_n290), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n207), .A2(KEYINPUT81), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT81), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G97), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n517), .B1(new_n530), .B2(new_n208), .ZN(new_n531));
  INV_X1    g0331(.A(new_n519), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT82), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n230), .B1(new_n533), .B2(new_n520), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n273), .A2(G77), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n297), .B2(new_n208), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n514), .B(new_n290), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n513), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(new_n332), .C1(new_n478), .C2(new_n479), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n481), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n255), .A2(G250), .A3(G1698), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n542), .A2(new_n489), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n293), .A2(new_n294), .A3(G244), .A4(new_n328), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT4), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(KEYINPUT84), .A3(new_n545), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT84), .B1(new_n544), .B2(new_n545), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n543), .B(new_n546), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n541), .B1(new_n550), .B2(new_n333), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G179), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n434), .B2(new_n551), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n539), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G87), .A2(G107), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n490), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n230), .B1(new_n383), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n255), .A2(new_n230), .A3(G68), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n490), .B2(new_n366), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n309), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(new_n290), .B1(new_n563), .B2(new_n413), .ZN(new_n564));
  INV_X1    g0364(.A(new_n413), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n487), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n293), .A2(new_n294), .A3(G244), .A4(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n293), .A2(new_n294), .A3(G238), .A4(new_n328), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n259), .C2(new_n492), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n333), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n342), .A2(G250), .A3(new_n332), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n313), .A2(new_n332), .A3(G45), .A4(G274), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n434), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n573), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n333), .B2(new_n570), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n345), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n567), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n354), .B1(new_n571), .B2(new_n574), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n487), .A2(G87), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n571), .A2(new_n574), .A3(G190), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n582), .A2(new_n564), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G264), .B(new_n332), .C1(new_n478), .C2(new_n479), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n293), .A2(new_n294), .A3(G257), .A4(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n293), .A2(new_n294), .A3(G250), .A4(new_n328), .ZN(new_n589));
  XOR2_X1   g0389(.A(KEYINPUT88), .B(G294), .Z(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n259), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n333), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT89), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n481), .B(new_n587), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT89), .B1(new_n591), .B2(new_n333), .ZN(new_n595));
  OAI21_X1  g0395(.A(G169), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n592), .A2(new_n481), .A3(new_n587), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n597), .A2(new_n345), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n255), .A2(new_n230), .A3(G87), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT22), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(KEYINPUT87), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n602), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n255), .A2(new_n604), .A3(new_n230), .A4(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT24), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n366), .A2(new_n492), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT23), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n230), .B2(G107), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n208), .A2(KEYINPUT23), .A3(G20), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n607), .B1(new_n606), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n290), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT25), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n309), .B2(G107), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n563), .A2(KEYINPUT25), .A3(new_n208), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n617), .A2(new_n618), .B1(new_n487), .B2(G107), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n599), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n594), .A2(G190), .A3(new_n595), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n597), .A2(new_n354), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n615), .B(new_n619), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n586), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n513), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n290), .B1(new_n534), .B2(new_n536), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT83), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n626), .B1(new_n628), .B2(new_n537), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n551), .A2(G190), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n550), .A2(new_n333), .ZN(new_n632));
  INV_X1    g0432(.A(new_n541), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n630), .A2(new_n631), .B1(new_n634), .B2(G200), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n551), .A2(KEYINPUT85), .A3(G190), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n511), .A2(new_n554), .A3(new_n625), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n469), .A2(new_n638), .ZN(G372));
  NAND3_X1  g0439(.A1(new_n318), .A2(new_n408), .A3(new_n348), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT18), .B1(new_n321), .B2(new_n347), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n436), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n402), .A2(new_n403), .B1(new_n644), .B2(new_n395), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n362), .A2(new_n360), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n643), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n463), .A2(new_n464), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n648), .A2(new_n650), .B1(new_n454), .B2(new_n453), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT90), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n578), .B2(G169), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n575), .A2(KEYINPUT90), .A3(new_n434), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n564), .A2(new_n566), .B1(new_n578), .B2(new_n345), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n581), .B1(G190), .B2(new_n578), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n564), .A2(new_n583), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n655), .A2(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n624), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n509), .A2(new_n507), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n621), .A2(new_n661), .A3(new_n506), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n554), .A2(new_n660), .A3(new_n637), .A4(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n539), .A2(new_n659), .A3(new_n664), .A4(new_n553), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n655), .A2(new_n656), .ZN(new_n666));
  AOI211_X1 g0466(.A(new_n345), .B(new_n541), .C1(new_n550), .C2(new_n333), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n434), .B1(new_n632), .B2(new_n633), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n580), .A2(new_n585), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n629), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n665), .B(new_n666), .C1(new_n671), .C2(new_n664), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n651), .B1(new_n469), .B2(new_n673), .ZN(G369));
  AND2_X1   g0474(.A1(new_n230), .A2(G13), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n313), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n676), .A2(KEYINPUT91), .A3(KEYINPUT27), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT91), .B1(new_n676), .B2(KEYINPUT27), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(G213), .B1(new_n676), .B2(KEYINPUT27), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n511), .B1(new_n498), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n510), .A2(new_n497), .A3(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n621), .B2(new_n685), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n596), .A2(new_n598), .B1(new_n615), .B2(new_n619), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(KEYINPUT93), .A3(new_n684), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n620), .A2(new_n684), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n620), .A2(KEYINPUT92), .A3(new_n684), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(new_n621), .A3(new_n624), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n690), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n510), .A2(new_n685), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n695), .B2(new_n700), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n621), .A2(new_n684), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n226), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n339), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n556), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(G1), .ZN(new_n712));
  INV_X1    g0512(.A(new_n232), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n710), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n685), .B1(new_n663), .B2(new_n672), .ZN(new_n716));
  XNOR2_X1  g0516(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT96), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n660), .A2(new_n637), .A3(new_n554), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT97), .B1(new_n510), .B2(new_n693), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT97), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n621), .A2(new_n661), .A3(new_n723), .A4(new_n506), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n659), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT26), .B1(new_n554), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n629), .A2(new_n669), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n664), .A3(new_n586), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n666), .A3(new_n730), .ZN(new_n731));
  OAI211_X1 g0531(.A(KEYINPUT29), .B(new_n685), .C1(new_n726), .C2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n716), .A2(KEYINPUT96), .A3(new_n717), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n720), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  AND4_X1   g0535(.A1(new_n571), .A2(new_n592), .A3(new_n574), .A4(new_n587), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n551), .A2(new_n508), .A3(G179), .A4(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT94), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n737), .B2(new_n738), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n483), .A2(new_n345), .A3(new_n575), .A4(new_n597), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n551), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n735), .B1(new_n744), .B2(new_n685), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n741), .A2(new_n743), .ZN(new_n746));
  OAI211_X1 g0546(.A(KEYINPUT31), .B(new_n684), .C1(new_n746), .C2(new_n740), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n745), .B(new_n747), .C1(new_n638), .C2(new_n684), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n734), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n715), .B1(new_n751), .B2(G1), .ZN(G364));
  AOI21_X1  g0552(.A(new_n229), .B1(G20), .B2(new_n434), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n230), .B1(new_n755), .B2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n590), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n230), .A2(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n354), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n755), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G283), .A2(new_n761), .B1(new_n763), .B2(G329), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n345), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n230), .A2(new_n351), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n766), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n764), .B1(new_n765), .B2(new_n767), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n351), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n757), .B(new_n771), .C1(G326), .C2(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n769), .A2(new_n759), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT99), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT99), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G303), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n295), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT101), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n772), .A2(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n784), .B2(KEYINPUT102), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(KEYINPUT102), .B2(new_n784), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n774), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n756), .A2(new_n207), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n782), .B2(G68), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT100), .Z(new_n790));
  NAND2_X1  g0590(.A1(new_n763), .A2(G159), .ZN(new_n791));
  INV_X1    g0591(.A(new_n773), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(KEYINPUT32), .B1(new_n204), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(KEYINPUT32), .B2(new_n791), .ZN(new_n794));
  INV_X1    g0594(.A(new_n778), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G87), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n760), .A2(new_n208), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n255), .B1(new_n767), .B2(new_n365), .ZN(new_n798));
  INV_X1    g0598(.A(new_n770), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n797), .B(new_n798), .C1(new_n304), .C2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n790), .A2(new_n794), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n754), .B1(new_n787), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n753), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n251), .A2(G45), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT98), .Z(new_n809));
  NOR2_X1   g0609(.A1(new_n708), .A2(new_n255), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(G45), .C2(new_n713), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n708), .A2(new_n295), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n812), .A2(G355), .B1(new_n492), .B2(new_n708), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n807), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n336), .B1(new_n675), .B2(G45), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n709), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n802), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n805), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n688), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n689), .A2(new_n818), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n688), .A2(G330), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT103), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n684), .A2(new_n417), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n432), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n436), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n644), .A2(new_n685), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n716), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n685), .B(new_n832), .C1(new_n663), .C2(new_n672), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n749), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT105), .Z(new_n836));
  AOI21_X1  g0636(.A(new_n817), .B1(new_n834), .B2(new_n749), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n767), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G116), .A2(new_n839), .B1(new_n761), .B2(G87), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n841), .B2(new_n770), .C1(new_n778), .C2(new_n208), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n295), .B1(new_n762), .B2(new_n765), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n783), .A2(new_n844), .B1(new_n792), .B2(new_n779), .ZN(new_n845));
  NOR4_X1   g0645(.A1(new_n842), .A2(new_n788), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT104), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G143), .A2(new_n799), .B1(new_n839), .B2(G159), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n773), .A2(G137), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n783), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n795), .A2(G50), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n761), .A2(G68), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n763), .A2(G132), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n255), .ZN(new_n858));
  INV_X1    g0658(.A(new_n756), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n304), .B2(new_n859), .ZN(new_n860));
  AND4_X1   g0660(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n753), .B1(new_n847), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n753), .A2(new_n803), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n818), .B1(new_n365), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n862), .B(new_n864), .C1(new_n832), .C2(new_n804), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n838), .A2(new_n865), .ZN(G384));
  OAI211_X1 g0666(.A(new_n403), .B(new_n684), .C1(new_n402), .C2(new_n396), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n401), .A2(new_n399), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n393), .A2(new_n389), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n400), .B1(new_n869), .B2(G169), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n403), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n403), .A2(new_n684), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n395), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n830), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n748), .A2(new_n874), .A3(KEYINPUT40), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT106), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n361), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n318), .A2(new_n348), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n321), .A2(KEYINPUT106), .A3(new_n357), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n405), .A2(new_n406), .A3(new_n682), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT107), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n361), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n405), .A2(new_n406), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n348), .ZN(new_n888));
  INV_X1    g0688(.A(new_n881), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT107), .B(KEYINPUT37), .C1(new_n880), .C2(new_n881), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n884), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n321), .A2(new_n357), .A3(new_n359), .ZN(new_n893));
  NOR2_X1   g0693(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n321), .B2(new_n357), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n641), .B(new_n640), .C1(new_n893), .C2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n896), .A2(KEYINPUT108), .A3(new_n881), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT108), .B1(new_n896), .B2(new_n881), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n892), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n288), .A2(new_n290), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT16), .B1(new_n265), .B2(new_n287), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n317), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n681), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n646), .B1(new_n407), .B2(new_n408), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n349), .A2(KEYINPUT18), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n348), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n906), .A3(new_n361), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n890), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(new_n914), .A3(KEYINPUT38), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n875), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT109), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n748), .A2(new_n874), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n906), .B1(new_n363), .B2(new_n409), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n888), .A2(new_n889), .B1(new_n912), .B2(KEYINPUT37), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n901), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n918), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n917), .B1(new_n922), .B2(KEYINPUT40), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n748), .A2(new_n874), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n919), .A2(new_n920), .A3(new_n901), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n910), .B2(new_n914), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(KEYINPUT109), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n916), .B1(new_n923), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n468), .A2(new_n748), .ZN(new_n932));
  OAI21_X1  g0732(.A(G330), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n867), .A2(new_n873), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n833), .A2(new_n829), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n925), .C2(new_n926), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n643), .B2(new_n681), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT39), .B1(new_n925), .B2(new_n926), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n892), .B2(new_n899), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n915), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n402), .A2(new_n403), .A3(new_n685), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n938), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n468), .A2(new_n720), .A3(new_n732), .A4(new_n733), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n947), .A2(new_n651), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n946), .B(new_n948), .Z(new_n949));
  OAI22_X1  g0749(.A1(new_n934), .A2(new_n949), .B1(new_n313), .B2(new_n675), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n934), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n521), .A2(new_n522), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT35), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(KEYINPUT35), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(G116), .A4(new_n231), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT36), .Z(new_n957));
  NAND3_X1  g0757(.A1(new_n232), .A2(G77), .A3(new_n268), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n204), .A2(G68), .ZN(new_n959));
  AOI211_X1 g0759(.A(G13), .B(new_n313), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n951), .A2(new_n957), .A3(new_n960), .ZN(G367));
  INV_X1    g0761(.A(new_n810), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n806), .B1(new_n226), .B2(new_n413), .C1(new_n243), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n817), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n795), .A2(new_n304), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n255), .B1(new_n770), .B2(new_n850), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G159), .B2(new_n782), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n859), .A2(G68), .B1(G143), .B2(new_n773), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n760), .A2(new_n365), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n767), .A2(new_n204), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(G137), .C2(new_n763), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n965), .A2(new_n967), .A3(new_n968), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n795), .A2(G116), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT46), .ZN(new_n974));
  INV_X1    g0774(.A(new_n590), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n973), .A2(new_n974), .B1(new_n975), .B2(new_n782), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n974), .B2(new_n973), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT116), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n799), .A2(G303), .B1(new_n761), .B2(new_n530), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n844), .B2(new_n767), .ZN(new_n981));
  XOR2_X1   g0781(.A(KEYINPUT115), .B(G311), .Z(new_n982));
  NOR2_X1   g0782(.A1(new_n792), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n255), .B1(new_n763), .B2(G317), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n208), .B2(new_n756), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n981), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n977), .B2(new_n978), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n972), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT117), .B(KEYINPUT47), .Z(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n964), .B1(new_n990), .B2(new_n753), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n685), .A2(new_n658), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(new_n656), .A3(new_n655), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n727), .B2(new_n992), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(new_n820), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT110), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n554), .B2(new_n685), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n729), .A2(KEYINPUT110), .A3(new_n684), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n554), .B(new_n637), .C1(new_n629), .C2(new_n685), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(KEYINPUT111), .A3(new_n704), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT111), .B1(new_n1002), .B2(new_n704), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT42), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1005), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT42), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n1008), .A3(new_n1003), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n554), .B1(new_n1010), .B2(new_n621), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n685), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1006), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT112), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1014), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1016), .A2(new_n1017), .B1(KEYINPUT43), .B2(new_n994), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT112), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n702), .A2(new_n1010), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1018), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT114), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT113), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n701), .B1(new_n510), .B2(new_n685), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n704), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(new_n689), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n751), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n749), .A3(new_n734), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n706), .A2(new_n1002), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT45), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1010), .B(KEYINPUT44), .C1(new_n704), .C2(new_n705), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT44), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n706), .B2(new_n1002), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n702), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n751), .B1(new_n1038), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n709), .B(KEYINPUT41), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n816), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1029), .A2(new_n1030), .A3(new_n1051), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n1018), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1025), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n815), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT114), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n996), .B1(new_n1052), .B2(new_n1058), .ZN(G387));
  NAND3_X1  g0859(.A1(new_n695), .A2(new_n700), .A3(new_n805), .ZN(new_n1060));
  INV_X1    g0860(.A(G45), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n810), .B1(new_n240), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n812), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1062), .B1(new_n711), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n411), .A2(G50), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT50), .ZN(new_n1066));
  AOI21_X1  g0866(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n711), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1064), .A2(new_n1068), .B1(new_n208), .B2(new_n708), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n817), .B1(new_n1069), .B2(new_n807), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G317), .A2(new_n799), .B1(new_n839), .B2(G303), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n783), .B2(new_n982), .C1(new_n768), .C2(new_n792), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n795), .A2(new_n975), .B1(G283), .B2(new_n859), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n760), .A2(new_n492), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n255), .B(new_n1081), .C1(G326), .C2(new_n763), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n305), .A2(new_n782), .B1(G68), .B2(new_n839), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT118), .Z(new_n1085));
  NOR2_X1   g0885(.A1(new_n756), .A2(new_n413), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G97), .A2(new_n761), .B1(new_n763), .B2(G150), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1087), .B(new_n255), .C1(new_n204), .C2(new_n770), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(G159), .C2(new_n773), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n365), .B2(new_n778), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1083), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1070), .B1(new_n1091), .B2(new_n753), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1034), .A2(new_n816), .B1(new_n1060), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n710), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT119), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1094), .A2(new_n1095), .B1(new_n751), .B2(new_n1034), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(G393));
  OR2_X1    g0898(.A1(new_n1048), .A2(new_n815), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n248), .A2(new_n810), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n806), .B1(new_n226), .B2(new_n490), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n817), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n799), .A2(G311), .B1(G317), .B2(new_n773), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT121), .B(KEYINPUT52), .Z(new_n1104));
  XNOR2_X1  g0904(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n783), .A2(new_n779), .B1(new_n756), .B2(new_n492), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n767), .A2(new_n841), .B1(new_n762), .B2(new_n768), .ZN(new_n1107));
  NOR4_X1   g0907(.A1(new_n1106), .A2(new_n1107), .A3(new_n255), .A4(new_n797), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1105), .B(new_n1108), .C1(new_n844), .C2(new_n778), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n763), .A2(G143), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n295), .B1(new_n761), .B2(G87), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n778), .C2(new_n216), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT120), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n799), .A2(G159), .B1(G150), .B2(new_n773), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT51), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n859), .A2(G77), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n411), .B2(new_n767), .C1(new_n783), .C2(new_n204), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1109), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1102), .B1(new_n1119), .B2(new_n753), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1002), .B2(new_n820), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1099), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1038), .A2(new_n1048), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT122), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT122), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1038), .A2(new_n1048), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1038), .A2(new_n1048), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(new_n710), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1122), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(G390));
  INV_X1    g0931(.A(new_n863), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G107), .A2(new_n782), .B1(new_n773), .B2(G283), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n856), .A2(new_n1133), .A3(new_n1116), .A4(new_n295), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G116), .A2(new_n799), .B1(new_n839), .B2(new_n530), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n841), .B2(new_n762), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G87), .C2(new_n795), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G50), .A2(new_n761), .B1(new_n763), .B2(G125), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n295), .B1(new_n799), .B2(G132), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n778), .A2(new_n850), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT53), .Z(new_n1142));
  AOI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(G128), .C2(new_n773), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n767), .A2(new_n1144), .B1(new_n756), .B2(new_n275), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G137), .B2(new_n782), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT124), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1137), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n817), .B1(new_n305), .B2(new_n1132), .C1(new_n1148), .C2(new_n754), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n943), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n803), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n936), .A2(new_n935), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n944), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n939), .B(new_n1154), .C1(new_n940), .C2(new_n942), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n748), .A2(G330), .A3(new_n832), .A4(new_n935), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT123), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n685), .B1(new_n726), .B2(new_n731), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n828), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n829), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n935), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(new_n944), .C1(new_n925), .C2(new_n940), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1155), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1158), .B1(new_n1155), .B2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1152), .B1(new_n1166), .B2(new_n815), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n468), .A2(G330), .A3(new_n748), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n947), .A2(new_n651), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n935), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n749), .B2(new_n830), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1156), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n936), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n829), .A3(new_n1174), .A4(new_n1156), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1169), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n710), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1167), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(G378));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1169), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(KEYINPUT40), .B(new_n924), .C1(new_n940), .C2(new_n925), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT109), .B1(new_n927), .B2(new_n928), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n922), .A2(new_n917), .A3(KEYINPUT40), .ZN(new_n1187));
  OAI211_X1 g0987(.A(G330), .B(new_n1185), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n650), .A2(new_n455), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n445), .A2(new_n682), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1189), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1188), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n930), .A2(G330), .A3(new_n1194), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1196), .A2(new_n946), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n946), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1184), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n946), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n929), .A2(new_n923), .ZN(new_n1202));
  AND4_X1   g1002(.A1(G330), .A2(new_n1202), .A3(new_n1185), .A4(new_n1194), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1194), .B1(new_n930), .B2(G330), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1196), .A2(new_n946), .A3(new_n1197), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1205), .A2(new_n1206), .B1(new_n1183), .B2(new_n1179), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n709), .B(new_n1200), .C1(new_n1207), .C2(KEYINPUT57), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1195), .A2(new_n803), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n817), .B1(G50), .B2(new_n1132), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n339), .A2(new_n255), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G50), .B(new_n1211), .C1(new_n259), .C2(new_n476), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n783), .A2(new_n207), .B1(new_n792), .B2(new_n492), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n844), .B2(new_n762), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G68), .C2(new_n859), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n767), .A2(new_n413), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n760), .A2(new_n303), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G107), .C2(new_n799), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1215), .B(new_n1218), .C1(new_n365), .C2(new_n778), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT58), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1212), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1144), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n795), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n782), .A2(G132), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G128), .A2(new_n799), .B1(new_n839), .B2(G137), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n859), .A2(G150), .B1(G125), .B2(new_n773), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n259), .B(new_n476), .C1(new_n760), .C2(new_n275), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G124), .B2(new_n763), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1221), .B1(new_n1220), .B2(new_n1219), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1210), .B1(new_n1233), .B2(new_n753), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1209), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(new_n816), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1208), .A2(new_n1238), .ZN(G375));
  NAND2_X1  g1039(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1169), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n1177), .A3(new_n1050), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1170), .A2(new_n803), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n817), .B1(G68), .B2(new_n1132), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G107), .A2(new_n839), .B1(new_n763), .B2(G303), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n844), .B2(new_n770), .C1(new_n778), .C2(new_n207), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n295), .B1(new_n760), .B2(new_n365), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n783), .A2(new_n492), .B1(new_n792), .B2(new_n841), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1247), .A2(new_n1086), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1251), .A2(KEYINPUT125), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n795), .A2(G159), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n295), .B(new_n1217), .C1(G50), .C2(new_n859), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1222), .A2(new_n782), .B1(G132), .B2(new_n773), .ZN(new_n1255));
  INV_X1    g1055(.A(G128), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n767), .A2(new_n850), .B1(new_n762), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G137), .B2(new_n799), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1251), .A2(KEYINPUT125), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1252), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1245), .B1(new_n1261), .B2(new_n753), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1240), .A2(new_n816), .B1(new_n1244), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1243), .A2(new_n1263), .ZN(G381));
  OR4_X1    g1064(.A1(G384), .A2(G390), .A3(G378), .A4(G381), .ZN(new_n1265));
  OR2_X1    g1065(.A1(G393), .A2(G396), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G387), .A2(new_n1265), .A3(G375), .A4(new_n1266), .ZN(G407));
  NAND2_X1  g1067(.A1(new_n683), .A2(G213), .ZN(new_n1268));
  OR3_X1    g1068(.A1(G375), .A2(G378), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(G407), .A2(G213), .A3(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1242), .B1(new_n1271), .B2(new_n1176), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1241), .A2(KEYINPUT60), .A3(new_n1169), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n709), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1263), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n865), .A3(new_n838), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(G384), .A3(new_n1263), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1208), .A2(G378), .A3(new_n1238), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1236), .B1(new_n1207), .B2(new_n1050), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1205), .A2(KEYINPUT126), .A3(new_n1206), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n816), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1268), .B(new_n1279), .C1(new_n1280), .C2(new_n1286), .ZN(new_n1287));
  XOR2_X1   g1087(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1268), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n683), .A2(G213), .A3(G2897), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1278), .B(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1283), .A2(new_n816), .A3(new_n1284), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1237), .A2(new_n1050), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1235), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1180), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1208), .A2(G378), .A3(new_n1238), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1268), .A4(new_n1279), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1289), .A2(new_n1293), .A3(new_n1294), .A4(new_n1303), .ZN(new_n1304));
  XOR2_X1   g1104(.A(G393), .B(G396), .Z(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1030), .B1(new_n1029), .B2(new_n1051), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1055), .A2(new_n1057), .A3(KEYINPUT114), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G390), .B1(new_n1309), .B2(new_n996), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n996), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1311), .B(new_n1130), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1306), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G387), .A2(new_n1130), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1309), .A2(new_n996), .A3(G390), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1305), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1304), .A2(new_n1317), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1287), .A2(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1301), .A2(KEYINPUT63), .A3(new_n1268), .A4(new_n1279), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1319), .A2(new_n1320), .A3(new_n1322), .A4(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1318), .A2(new_n1324), .ZN(G405));
  NAND2_X1  g1125(.A1(G375), .A2(new_n1180), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1326), .A2(new_n1278), .A3(new_n1300), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1278), .B1(new_n1326), .B2(new_n1300), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1319), .B(new_n1329), .ZN(G402));
endmodule


