//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G77), .B2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT65), .B(G238), .Z(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT66), .Z(new_n225));
  NOR3_X1   g0025(.A1(new_n220), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n205), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n204), .ZN(new_n235));
  NOR2_X1   g0035(.A1(G58), .A2(G68), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G50), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  AOI211_X1 g0039(.A(new_n210), .B(new_n228), .C1(new_n235), .C2(new_n239), .ZN(G361));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n219), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G270), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(KEYINPUT68), .B(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G68), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G222), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n262), .B(new_n264), .C1(new_n265), .C2(new_n263), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n231), .A2(new_n232), .B1(G33), .B2(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n266), .B(new_n267), .C1(G77), .C2(new_n262), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n269), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n268), .B(new_n272), .C1(new_n217), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G200), .ZN(new_n277));
  INV_X1    g0077(.A(G190), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n231), .A2(new_n232), .A3(new_n280), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n206), .A2(new_n204), .A3(G1), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(new_n204), .B2(G1), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n203), .A2(KEYINPUT69), .A3(G20), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n216), .ZN(new_n289));
  OAI21_X1  g0089(.A(G20), .B1(new_n237), .B2(G50), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n204), .A2(new_n259), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n204), .A2(G33), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n290), .B1(new_n291), .B2(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n281), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n288), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n279), .B1(new_n297), .B2(KEYINPUT9), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n297), .A2(KEYINPUT71), .A3(KEYINPUT9), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT71), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n288), .A2(new_n289), .A3(new_n296), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n277), .B(new_n298), .C1(new_n299), .C2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT10), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n276), .A2(G179), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n276), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G77), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n293), .A2(new_n292), .B1(new_n204), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT70), .ZN(new_n312));
  XOR2_X1   g0112(.A(KEYINPUT15), .B(G87), .Z(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(new_n294), .B2(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n281), .B1(new_n310), .B2(new_n282), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n221), .A2(new_n263), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n262), .B1(new_n213), .B2(G1698), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n267), .B1(G107), .B2(new_n262), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n275), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G244), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n272), .A3(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n322), .A2(new_n278), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(G200), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n287), .A2(G77), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n316), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n316), .A2(new_n325), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n307), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n327), .B(new_n328), .C1(G179), .C2(new_n322), .ZN(new_n329));
  AND4_X1   g0129(.A1(new_n305), .A2(new_n309), .A3(new_n326), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n282), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n293), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n287), .B2(new_n293), .ZN(new_n333));
  AND3_X1   g0133(.A1(KEYINPUT76), .A2(G58), .A3(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT76), .B1(G58), .B2(G68), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n334), .A2(new_n335), .A3(new_n236), .ZN(new_n336));
  INV_X1    g0136(.A(G159), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n336), .A2(new_n204), .B1(new_n337), .B2(new_n292), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n260), .A2(new_n204), .A3(new_n261), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n261), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G68), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n339), .A2(new_n345), .A3(KEYINPUT16), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n281), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(KEYINPUT77), .A3(new_n343), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n343), .A2(KEYINPUT77), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(G68), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT16), .B1(new_n350), .B2(new_n339), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n333), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G179), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT79), .B1(new_n275), .B2(new_n213), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT79), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n274), .A2(new_n269), .A3(new_n355), .A4(G232), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n272), .A3(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n260), .A2(new_n261), .B1(new_n217), .B2(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n265), .A2(new_n263), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n358), .A2(new_n359), .B1(G33), .B2(G87), .ZN(new_n360));
  INV_X1    g0160(.A(new_n267), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT78), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(KEYINPUT3), .A2(G33), .ZN(new_n363));
  NOR2_X1   g0163(.A1(KEYINPUT3), .A2(G33), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n359), .B1(G226), .B2(new_n263), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G87), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT78), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n267), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n357), .B1(new_n362), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n357), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n267), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n353), .A2(new_n370), .B1(new_n373), .B2(new_n307), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n352), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT18), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n347), .A2(new_n351), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n370), .A2(new_n278), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n377), .A2(new_n381), .A3(KEYINPUT17), .A4(new_n333), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n352), .A2(new_n374), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT17), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n278), .A2(new_n370), .B1(new_n373), .B2(new_n379), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n352), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n376), .A2(new_n382), .A3(new_n384), .A4(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(G232), .B(G1698), .C1(new_n363), .C2(new_n364), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT72), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n262), .A2(new_n392), .A3(G232), .A4(G1698), .ZN(new_n393));
  AND3_X1   g0193(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n262), .A2(G226), .A3(new_n263), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n391), .A2(new_n393), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT74), .ZN(new_n400));
  AOI21_X1  g0200(.A(G1698), .B1(new_n260), .B2(new_n261), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n396), .B1(new_n401), .B2(G226), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT74), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n391), .A4(new_n393), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n267), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n271), .B1(new_n320), .B2(G238), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G190), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n294), .A2(new_n310), .B1(new_n204), .B2(G68), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT75), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n292), .A2(new_n216), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n281), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XOR2_X1   g0215(.A(new_n415), .B(KEYINPUT11), .Z(new_n416));
  NAND2_X1  g0216(.A1(new_n282), .A2(new_n222), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT12), .ZN(new_n418));
  INV_X1    g0218(.A(new_n287), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(new_n222), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(G200), .B1(new_n408), .B2(new_n409), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n411), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n421), .ZN(new_n425));
  OAI21_X1  g0225(.A(G169), .B1(new_n408), .B2(new_n409), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT14), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n410), .A2(G179), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(G169), .C1(new_n408), .C2(new_n409), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n424), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n330), .A2(new_n389), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G116), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n259), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n204), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n204), .A2(G107), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT23), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n204), .B(G87), .C1(new_n363), .C2(new_n364), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n439), .A2(KEYINPUT22), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(KEYINPUT22), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n436), .B(new_n438), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT85), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n439), .B(KEYINPUT22), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(KEYINPUT85), .A3(new_n436), .A4(new_n438), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(KEYINPUT24), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT24), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n281), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n283), .B1(G1), .B2(new_n259), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(new_n218), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT25), .ZN(new_n453));
  AOI211_X1 g0253(.A(G107), .B(new_n331), .C1(KEYINPUT86), .C2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(KEYINPUT86), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n450), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(G250), .A2(G1698), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n262), .B(new_n458), .C1(G257), .C2(new_n263), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G294), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n267), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT5), .B(G41), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n464), .A2(new_n270), .A3(G1), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n274), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n464), .A2(G1), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G264), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n462), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G169), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n353), .B2(new_n471), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n457), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n283), .B(G116), .C1(G1), .C2(new_n259), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n331), .A2(G116), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n434), .A2(G20), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  INV_X1    g0279(.A(G97), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n479), .B(new_n204), .C1(G33), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n281), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT20), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n482), .A2(new_n483), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n475), .B(new_n477), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n263), .A2(G257), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G264), .A2(G1698), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(new_n363), .C2(new_n364), .ZN(new_n489));
  INV_X1    g0289(.A(G303), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n260), .A2(new_n490), .A3(new_n261), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(KEYINPUT84), .A3(new_n491), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n267), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n469), .A2(G270), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n466), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n486), .A2(new_n498), .A3(G169), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT21), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(G179), .A3(new_n486), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n486), .A2(new_n498), .A3(KEYINPUT21), .A4(G169), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n474), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n498), .A2(new_n278), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n486), .B(new_n508), .C1(G200), .C2(new_n498), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(new_n263), .C1(new_n363), .C2(new_n364), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n512), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n262), .A2(G244), .A3(new_n263), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n262), .A2(G250), .A3(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n513), .A2(new_n515), .A3(new_n479), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n267), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n469), .A2(G257), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n466), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G169), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n518), .A2(G179), .A3(new_n466), .A4(new_n519), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n282), .A2(new_n480), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n451), .B2(new_n480), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n348), .A2(G107), .A3(new_n349), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n218), .A2(KEYINPUT6), .A3(G97), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n480), .A2(new_n218), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G97), .A2(G107), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n530), .B2(KEYINPUT6), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G20), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n204), .A2(new_n259), .A3(G77), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n526), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n525), .B1(new_n534), .B2(new_n281), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT81), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI211_X1 g0337(.A(KEYINPUT81), .B(new_n525), .C1(new_n534), .C2(new_n281), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n523), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n520), .A2(G200), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n518), .A2(G190), .A3(new_n466), .A4(new_n519), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n535), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G244), .B(G1698), .C1(new_n363), .C2(new_n364), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n435), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(KEYINPUT82), .A2(new_n543), .B1(new_n401), .B2(G238), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n361), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(G250), .B1(new_n464), .B2(G1), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n274), .B1(new_n550), .B2(new_n465), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n307), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n401), .A2(G238), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n544), .B2(new_n545), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n543), .A2(KEYINPUT82), .B1(new_n259), .B2(new_n434), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n267), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n353), .A3(new_n551), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n331), .A2(new_n313), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n283), .B(new_n313), .C1(G1), .C2(new_n259), .ZN(new_n561));
  NOR3_X1   g0361(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT73), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(KEYINPUT19), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n562), .B1(new_n567), .B2(new_n204), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n204), .B(G68), .C1(new_n363), .C2(new_n364), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n294), .A2(new_n480), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(KEYINPUT19), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n281), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n560), .B(new_n561), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n553), .A2(new_n558), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G87), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n259), .A2(G1), .ZN(new_n578));
  NOR4_X1   g0378(.A1(new_n281), .A2(new_n282), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n571), .A2(KEYINPUT19), .ZN(new_n580));
  AOI21_X1  g0380(.A(G20), .B1(new_n396), .B2(KEYINPUT19), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n569), .B(new_n580), .C1(new_n581), .C2(new_n562), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n559), .B(new_n579), .C1(new_n582), .C2(new_n281), .ZN(new_n583));
  OAI21_X1  g0383(.A(G200), .B1(new_n548), .B2(new_n552), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n557), .A2(G190), .A3(new_n551), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n542), .A2(new_n576), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT83), .B1(new_n539), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n542), .A2(new_n576), .A3(new_n586), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n534), .A2(new_n281), .ZN(new_n591));
  INV_X1    g0391(.A(new_n525), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n521), .A2(new_n522), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n535), .A2(new_n536), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n589), .A2(new_n590), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n588), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n462), .A2(new_n470), .A3(new_n278), .A4(new_n466), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n471), .B2(G200), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n450), .A2(new_n452), .A3(new_n456), .A4(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n433), .A2(new_n510), .A3(new_n599), .A4(new_n602), .ZN(G372));
  NAND2_X1  g0403(.A1(new_n431), .A2(new_n425), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n424), .B1(new_n604), .B2(new_n329), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n387), .A3(new_n382), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n376), .A2(new_n384), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n305), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n309), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n433), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n586), .A2(new_n576), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n597), .A2(new_n613), .A3(new_n542), .A4(new_n602), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n505), .B1(new_n457), .B2(new_n473), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n576), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT87), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n595), .A2(new_n586), .A3(new_n576), .A4(new_n593), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n539), .A2(KEYINPUT26), .A3(new_n613), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n539), .A2(KEYINPUT87), .A3(KEYINPUT26), .A4(new_n613), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n616), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n611), .B1(new_n612), .B2(new_n625), .ZN(G369));
  NOR2_X1   g0426(.A1(new_n206), .A2(G20), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n203), .ZN(new_n628));
  XNOR2_X1  g0428(.A(KEYINPUT88), .B(KEYINPUT27), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G343), .ZN(new_n633));
  XOR2_X1   g0433(.A(new_n633), .B(KEYINPUT89), .Z(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n486), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n505), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n505), .ZN(new_n638));
  OR3_X1    g0438(.A1(new_n637), .A2(new_n638), .A3(new_n509), .ZN(new_n639));
  INV_X1    g0439(.A(G330), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n457), .A2(new_n635), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(KEYINPUT90), .A3(new_n602), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n643), .B(new_n474), .C1(KEYINPUT90), .C2(new_n642), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n457), .A2(new_n473), .A3(new_n634), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n645), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n505), .A2(new_n634), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT91), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n644), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n652), .ZN(G399));
  NAND2_X1  g0453(.A1(new_n562), .A2(new_n434), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT92), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n207), .A2(G41), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n655), .A2(new_n203), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n239), .B2(new_n656), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT28), .Z(new_n659));
  INV_X1    g0459(.A(KEYINPUT94), .ZN(new_n660));
  INV_X1    g0460(.A(new_n576), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n589), .A2(new_n597), .A3(new_n602), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n507), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n586), .A2(new_n576), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n597), .A2(new_n619), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n624), .B1(new_n665), .B2(new_n620), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n635), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n660), .B1(new_n667), .B2(KEYINPUT29), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT29), .ZN(new_n669));
  OAI211_X1 g0469(.A(KEYINPUT94), .B(new_n669), .C1(new_n625), .C2(new_n635), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n507), .A2(new_n589), .A3(new_n597), .A4(new_n602), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n537), .A2(new_n538), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n613), .A3(new_n619), .A4(new_n595), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n618), .A2(KEYINPUT26), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n676), .A3(new_n576), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT95), .B1(new_n677), .B2(new_n634), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  OAI211_X1 g0479(.A(KEYINPUT95), .B(new_n634), .C1(new_n616), .C2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT29), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n671), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n599), .A2(new_n510), .A3(new_n602), .A4(new_n634), .ZN(new_n684));
  INV_X1    g0484(.A(new_n471), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n520), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n548), .A2(new_n552), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G179), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n498), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n686), .A2(new_n688), .A3(KEYINPUT93), .A4(new_n498), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n687), .A2(new_n462), .A3(new_n470), .ZN(new_n694));
  INV_X1    g0494(.A(new_n522), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n502), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n694), .A2(new_n502), .A3(KEYINPUT30), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n635), .B1(new_n693), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n689), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT31), .B(new_n635), .C1(new_n700), .C2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n684), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n683), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n659), .B1(new_n709), .B2(G1), .ZN(G364));
  INV_X1    g0510(.A(new_n641), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n203), .B1(new_n627), .B2(G45), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n656), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT96), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n639), .A2(new_n640), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n711), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT97), .Z(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n639), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n234), .B1(G20), .B2(new_n307), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n204), .A2(G190), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n353), .A2(G200), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G311), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n204), .A2(new_n278), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n379), .A2(G179), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT98), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT98), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G303), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n725), .A2(new_n731), .ZN(new_n738));
  INV_X1    g0538(.A(G283), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n725), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G329), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n353), .A2(new_n379), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n730), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n743), .B1(G326), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n748));
  INV_X1    g0548(.A(G317), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n744), .A2(new_n725), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n740), .A2(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n262), .B1(new_n755), .B2(G294), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n737), .A2(new_n747), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n730), .A2(new_n726), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n729), .B(new_n757), .C1(G322), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n755), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n480), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n736), .A2(G87), .ZN(new_n763));
  INV_X1    g0563(.A(new_n738), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n752), .A2(G68), .B1(new_n764), .B2(G107), .ZN(new_n765));
  INV_X1    g0565(.A(new_n262), .ZN(new_n766));
  INV_X1    g0566(.A(new_n741), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(KEYINPUT32), .A3(G159), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT32), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n741), .B2(new_n337), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n766), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G50), .A2(new_n746), .B1(new_n759), .B2(G58), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n763), .A2(new_n765), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n727), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n762), .B(new_n773), .C1(G77), .C2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n724), .B1(new_n760), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n256), .A2(G45), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n207), .A2(new_n262), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n778), .C1(G45), .C2(new_n238), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n766), .A2(new_n207), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G355), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n779), .B(new_n781), .C1(G116), .C2(new_n208), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n724), .A2(new_n722), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n716), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n723), .A2(new_n776), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n719), .A2(new_n785), .ZN(G396));
  INV_X1    g0586(.A(new_n724), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G143), .A2(new_n759), .B1(new_n752), .B2(G150), .ZN(new_n788));
  INV_X1    g0588(.A(G137), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n788), .B1(new_n789), .B2(new_n745), .C1(new_n337), .C2(new_n727), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT34), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n262), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n790), .ZN(new_n793));
  INV_X1    g0593(.A(G132), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(KEYINPUT34), .B1(new_n794), .B2(new_n741), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n792), .B(new_n795), .C1(G58), .C2(new_n755), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n796), .B1(new_n216), .B2(new_n735), .C1(new_n222), .C2(new_n738), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n766), .B1(new_n727), .B2(new_n434), .C1(new_n739), .C2(new_n751), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n762), .B1(new_n736), .B2(G107), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n490), .B2(new_n745), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n798), .B(new_n800), .C1(G87), .C2(new_n764), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n802), .B2(new_n758), .C1(new_n728), .C2(new_n741), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n787), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n724), .A2(new_n720), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n716), .B(new_n804), .C1(new_n310), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n635), .A2(new_n327), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n326), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n329), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n329), .A2(new_n635), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n806), .B1(new_n721), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT100), .Z(new_n814));
  XNOR2_X1  g0614(.A(new_n667), .B(new_n811), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(new_n707), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n716), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G384));
  INV_X1    g0619(.A(KEYINPUT38), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT16), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n222), .B1(new_n342), .B2(new_n343), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n338), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n346), .A2(new_n823), .A3(new_n281), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n333), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT102), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n824), .A2(KEYINPUT102), .A3(new_n333), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n388), .A2(new_n632), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n362), .A2(new_n369), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n832), .A2(new_n353), .A3(new_n371), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n373), .A2(new_n307), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n632), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n352), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n377), .A2(new_n381), .A3(new_n333), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n837), .A2(new_n827), .A3(new_n828), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n840), .B1(new_n842), .B2(new_n839), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n820), .B1(new_n831), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n830), .B(KEYINPUT38), .C1(new_n843), .C2(new_n841), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(KEYINPUT31), .B(new_n635), .C1(new_n693), .C2(new_n700), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n684), .A2(new_n703), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n425), .A2(new_n635), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n604), .A2(new_n423), .A3(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n425), .B(new_n635), .C1(new_n424), .C2(new_n431), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n811), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n847), .A2(new_n849), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n838), .A2(new_n839), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n838), .A2(new_n840), .A3(new_n839), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n388), .A2(new_n352), .A3(new_n632), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n846), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n864), .A2(new_n849), .A3(KEYINPUT40), .A4(new_n853), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n856), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT104), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n433), .A2(new_n849), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n640), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n682), .A2(new_n433), .A3(new_n668), .A4(new_n670), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT103), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT103), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n671), .A2(new_n873), .A3(new_n433), .A4(new_n682), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n610), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n851), .A2(new_n852), .ZN(new_n876));
  INV_X1    g0676(.A(new_n666), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n634), .B(new_n812), .C1(new_n877), .C2(new_n616), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT101), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n810), .B(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n876), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n847), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  INV_X1    g0684(.A(new_n846), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n885), .B2(new_n862), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n604), .A2(new_n635), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT39), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n607), .A2(new_n632), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n883), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n875), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n870), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n203), .B2(new_n627), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n434), .B1(new_n531), .B2(KEYINPUT35), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n896), .B(new_n235), .C1(KEYINPUT35), .C2(new_n531), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT36), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n238), .A2(new_n334), .A3(new_n310), .A4(new_n335), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n222), .A2(G50), .ZN(new_n900));
  OAI211_X1 g0700(.A(G1), .B(new_n206), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(new_n898), .A3(new_n901), .ZN(G367));
  OR2_X1    g0702(.A1(new_n634), .A2(new_n583), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(new_n664), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  INV_X1    g0706(.A(new_n651), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n646), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n597), .B(new_n542), .C1(new_n535), .C2(new_n634), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n635), .A2(new_n593), .A3(new_n595), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT42), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n911), .B(KEYINPUT105), .Z(new_n914));
  OR2_X1    g0714(.A1(new_n914), .A2(new_n474), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n635), .B1(new_n915), .B2(new_n597), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n906), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n648), .A2(new_n914), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n919), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n656), .B(KEYINPUT41), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n652), .A2(new_n911), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT45), .ZN(new_n924));
  OR3_X1    g0724(.A1(new_n652), .A2(KEYINPUT44), .A3(new_n911), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT44), .B1(new_n652), .B2(new_n911), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n648), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n924), .B2(new_n927), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n646), .A2(new_n907), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n933), .A2(new_n711), .A3(new_n908), .ZN(new_n934));
  INV_X1    g0734(.A(new_n908), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n641), .B1(new_n935), .B2(new_n932), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n683), .A3(new_n707), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT106), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n937), .A2(new_n683), .A3(new_n940), .A4(new_n707), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n931), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n922), .B1(new_n942), .B2(new_n708), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n712), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n921), .A2(new_n944), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n727), .A2(new_n216), .B1(new_n741), .B2(new_n789), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n758), .A2(new_n291), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n761), .A2(new_n222), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n947), .B(new_n948), .C1(G143), .C2(new_n746), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n946), .B1(new_n949), .B2(KEYINPUT109), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n262), .B1(new_n738), .B2(new_n310), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G159), .B2(new_n752), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n950), .B(new_n952), .C1(new_n212), .C2(new_n735), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n949), .A2(KEYINPUT109), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n736), .A2(G116), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT46), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n262), .B1(new_n764), .B2(G97), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT107), .B(G311), .Z(new_n959));
  OAI22_X1  g0759(.A1(new_n745), .A2(new_n959), .B1(new_n758), .B2(new_n490), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n761), .A2(new_n218), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT108), .B(G317), .Z(new_n962));
  AOI211_X1 g0762(.A(new_n960), .B(new_n961), .C1(new_n767), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G294), .B2(new_n752), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n774), .A2(G283), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n955), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT47), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n724), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n904), .A2(new_n722), .ZN(new_n970));
  INV_X1    g0770(.A(new_n778), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n783), .B1(new_n208), .B2(new_n314), .C1(new_n248), .C2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n715), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n945), .A2(new_n973), .ZN(G387));
  INV_X1    g0774(.A(KEYINPUT110), .ZN(new_n975));
  INV_X1    g0775(.A(new_n938), .ZN(new_n976));
  INV_X1    g0776(.A(new_n656), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n938), .A2(KEYINPUT110), .A3(new_n656), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n709), .C2(new_n937), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n245), .A2(new_n464), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n981), .A2(new_n778), .B1(new_n655), .B2(new_n780), .ZN(new_n982));
  INV_X1    g0782(.A(new_n293), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n216), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT50), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n222), .A2(new_n310), .ZN(new_n986));
  NOR4_X1   g0786(.A1(new_n985), .A2(G45), .A3(new_n986), .A4(new_n655), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n982), .A2(new_n987), .B1(G107), .B2(new_n208), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n716), .B1(new_n988), .B2(new_n783), .ZN(new_n989));
  INV_X1    g0789(.A(new_n722), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n989), .B1(new_n647), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n761), .A2(new_n314), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n741), .A2(new_n291), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n992), .A2(new_n766), .A3(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n736), .A2(G77), .B1(G50), .B2(new_n759), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n480), .B2(new_n738), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(G159), .C2(new_n746), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n222), .B2(new_n727), .C1(new_n293), .C2(new_n751), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n759), .A2(new_n962), .B1(new_n774), .B2(G303), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n746), .A2(G322), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n751), .C2(new_n959), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT48), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n739), .B2(new_n761), .C1(new_n802), .C2(new_n735), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT49), .Z(new_n1004));
  AOI21_X1  g0804(.A(new_n262), .B1(new_n767), .B2(G326), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n434), .B2(new_n738), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n998), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n991), .B1(new_n724), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n937), .B2(new_n713), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n980), .A2(new_n1009), .ZN(G393));
  NAND2_X1  g0810(.A1(new_n914), .A2(new_n722), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n745), .A2(new_n749), .B1(new_n758), .B2(new_n728), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT52), .Z(new_n1013));
  AOI22_X1  g0813(.A1(new_n736), .A2(G283), .B1(G116), .B2(new_n755), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n766), .B1(new_n751), .B2(new_n490), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G322), .B2(new_n767), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1014), .B(new_n1016), .C1(new_n218), .C2(new_n738), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1013), .B(new_n1017), .C1(G294), .C2(new_n774), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n745), .A2(new_n291), .B1(new_n758), .B2(new_n337), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT111), .Z(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT51), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n736), .A2(G68), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n751), .A2(new_n216), .B1(new_n738), .B2(new_n577), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n983), .B2(new_n774), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n767), .A2(G143), .B1(new_n755), .B2(G77), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n262), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1021), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n724), .B1(new_n1018), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n253), .A2(new_n778), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n722), .B(new_n724), .C1(G97), .C2(new_n207), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n716), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1011), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n931), .B2(new_n712), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT112), .Z(new_n1034));
  AOI21_X1  g0834(.A(new_n942), .B1(new_n931), .B2(new_n938), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n656), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(G390));
  NOR2_X1   g0837(.A1(new_n868), .A2(new_n640), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n849), .A2(G330), .A3(new_n812), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n876), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n812), .B1(new_n678), .B2(new_n681), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n876), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1043), .A2(G330), .A3(new_n706), .A4(new_n812), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n881), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n849), .A2(G330), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n706), .A2(G330), .A3(new_n812), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1046), .A2(new_n853), .B1(new_n1047), .B2(new_n876), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n880), .B1(new_n667), .B2(new_n812), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n875), .A2(new_n1039), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n886), .A2(new_n888), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n882), .B2(new_n887), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1044), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n876), .B1(new_n1042), .B2(new_n881), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n887), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n864), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1053), .B(new_n1054), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1046), .A2(new_n853), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n634), .B1(new_n616), .B2(new_n679), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT95), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n811), .B1(new_n1064), .B2(new_n680), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1043), .B1(new_n1065), .B2(new_n880), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1057), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1061), .B1(new_n1068), .B2(new_n1053), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1059), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1051), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1056), .B1(new_n1049), .B2(new_n876), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1066), .A2(new_n1067), .B1(new_n1072), .B2(new_n1052), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1058), .B1(new_n1073), .B2(new_n1061), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1074), .A2(new_n875), .A3(new_n1039), .A4(new_n1050), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n656), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1052), .A2(new_n720), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n758), .A2(new_n434), .B1(new_n738), .B2(new_n222), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n763), .A2(new_n766), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT114), .Z(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n310), .B2(new_n761), .C1(new_n802), .C2(new_n741), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1078), .B(new_n1081), .C1(G107), .C2(new_n752), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n480), .B2(new_n727), .C1(new_n739), .C2(new_n745), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n738), .A2(new_n216), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n759), .A2(G132), .B1(new_n755), .B2(G159), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n789), .B2(new_n751), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n766), .B1(new_n767), .B2(G125), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n735), .A2(new_n291), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n1090));
  OAI211_X1 g0890(.A(new_n1087), .B(new_n1088), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1084), .B(new_n1091), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT54), .B(G143), .Z(new_n1093));
  NAND2_X1  g0893(.A1(new_n774), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n746), .A2(G128), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n787), .B1(new_n1083), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n716), .B(new_n1097), .C1(new_n293), .C2(new_n805), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1077), .A2(new_n1098), .B1(new_n1074), .B2(new_n713), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1076), .A2(new_n1099), .ZN(G378));
  INV_X1    g0900(.A(KEYINPUT57), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n856), .A2(G330), .A3(new_n865), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n305), .A2(new_n309), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1106), .A2(new_n1107), .B1(new_n297), .B2(new_n836), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1107), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n297), .A2(new_n836), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n1105), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1102), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1112), .A2(G330), .A3(new_n856), .A4(new_n865), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(KEYINPUT118), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n892), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1114), .A2(KEYINPUT118), .A3(new_n891), .A4(new_n1115), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n871), .A2(KEYINPUT103), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n871), .A2(KEYINPUT103), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n611), .B(new_n1039), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1074), .B2(new_n1050), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1101), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n610), .B(new_n1038), .C1(new_n872), .C2(new_n874), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1050), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1125), .B1(new_n1070), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n891), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1114), .A2(new_n892), .A3(new_n1115), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(KEYINPUT57), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1124), .A2(new_n1131), .A3(new_n656), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n713), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n216), .B1(new_n363), .B2(G41), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n761), .A2(new_n291), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n736), .A2(new_n1093), .B1(G128), .B2(new_n759), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT117), .Z(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n794), .B2(new_n751), .C1(new_n789), .C2(new_n727), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1136), .B(new_n1139), .C1(G125), .C2(new_n746), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT59), .ZN(new_n1141));
  AOI21_X1  g0941(.A(G33), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(G41), .B1(new_n767), .B2(G124), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(new_n337), .C2(new_n738), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1135), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n262), .C1(new_n767), .C2(G283), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n212), .B2(new_n738), .C1(new_n735), .C2(new_n310), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT115), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n751), .A2(new_n480), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n759), .A2(G107), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT116), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1149), .A2(new_n948), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n434), .B2(new_n745), .C1(new_n314), .C2(new_n727), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT58), .Z(new_n1155));
  OAI21_X1  g0955(.A(new_n724), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1112), .A2(new_n720), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n805), .A2(new_n216), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1156), .A2(new_n715), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1134), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1132), .A2(new_n1160), .ZN(G375));
  NAND2_X1  g0961(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n922), .A3(new_n1051), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n724), .A2(G68), .A3(new_n720), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n766), .B1(new_n802), .B2(new_n745), .C1(new_n735), .C2(new_n480), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n738), .A2(new_n310), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n434), .A2(new_n751), .B1(new_n758), .B2(new_n739), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n992), .A4(new_n1167), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n218), .B2(new_n727), .C1(new_n490), .C2(new_n741), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n727), .A2(new_n291), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n262), .B1(new_n738), .B2(new_n212), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n735), .A2(new_n337), .B1(new_n794), .B2(new_n745), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G50), .C2(new_n755), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n752), .A2(new_n1093), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n759), .A2(G137), .B1(new_n767), .B2(G128), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1169), .B1(new_n1170), .B2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n716), .B(new_n1164), .C1(new_n1177), .C2(new_n724), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n876), .A2(new_n720), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT119), .Z(new_n1180));
  AOI22_X1  g0980(.A1(new_n1050), .A2(new_n713), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1163), .A2(new_n1181), .ZN(G381));
  INV_X1    g0982(.A(G378), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1132), .A2(new_n1183), .A3(new_n1160), .ZN(new_n1184));
  INV_X1    g0984(.A(G390), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n973), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n921), .B2(new_n944), .ZN(new_n1187));
  INV_X1    g0987(.A(G396), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n980), .A2(new_n1188), .A3(new_n1009), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1189), .A2(G381), .A3(G384), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1185), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1184), .B1(new_n1192), .B2(KEYINPUT120), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(KEYINPUT120), .B2(new_n1192), .ZN(G407));
  OAI211_X1 g0994(.A(G407), .B(G213), .C1(G343), .C2(new_n1184), .ZN(G409));
  AOI21_X1  g0995(.A(new_n1183), .B1(new_n1132), .B2(new_n1160), .ZN(new_n1196));
  INV_X1    g0996(.A(G213), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(G343), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1127), .A2(new_n922), .A3(new_n1133), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1129), .A2(new_n713), .A3(new_n1130), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT121), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(new_n1159), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1099), .A3(new_n1203), .A4(new_n1076), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n1201), .B2(new_n1159), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1196), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT125), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n818), .A2(KEYINPUT123), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n818), .A2(KEYINPUT123), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT60), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1162), .B2(new_n1051), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1050), .B1(new_n875), .B2(new_n1039), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n656), .B1(new_n1215), .B2(KEYINPUT60), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT122), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n875), .A2(new_n1039), .A3(new_n1050), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT60), .B1(new_n1218), .B2(new_n1215), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n977), .B1(new_n1162), .B2(new_n1213), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT122), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1217), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1181), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1211), .B(new_n1212), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1217), .B2(new_n1222), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(KEYINPUT123), .A3(new_n818), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1198), .A2(G2897), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1225), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1226), .A2(KEYINPUT123), .A3(new_n818), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1212), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1226), .A2(new_n1210), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1228), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1208), .A2(KEYINPUT125), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1209), .A2(new_n1230), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(new_n1208), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1187), .A2(G390), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1189), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1188), .B1(new_n980), .B2(new_n1009), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT126), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G387), .A2(new_n1185), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1189), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1246), .A2(new_n1187), .A3(G390), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1239), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1242), .A2(new_n1187), .A3(new_n1243), .A4(G390), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1238), .A2(KEYINPUT63), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1207), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT124), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1207), .B(new_n1255), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1236), .A2(new_n1250), .A3(new_n1251), .A4(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT62), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1234), .A2(new_n1208), .A3(new_n1230), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1251), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1252), .A2(KEYINPUT62), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1263), .B2(new_n1264), .ZN(G405));
  INV_X1    g1065(.A(new_n1196), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1184), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1184), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1248), .A2(new_n1249), .A3(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1267), .A2(new_n1237), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1237), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(G402));
endmodule


