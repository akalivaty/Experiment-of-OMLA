//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G116), .ZN(new_n210));
  INV_X1    g0010(.A(G270), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n203), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n212), .B(new_n216), .C1(G77), .C2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT67), .Z(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n217), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NOR2_X1   g0025(.A1(new_n223), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND3_X1  g0029(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT66), .Z(new_n231));
  NAND3_X1  g0031(.A1(new_n204), .A2(G50), .A3(new_n205), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n225), .B(new_n229), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n214), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n221), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n211), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT7), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT74), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n253), .A4(new_n254), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n259), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT74), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(G68), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G58), .A2(G68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT75), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G58), .A3(G68), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n204), .A2(new_n265), .A3(new_n267), .A4(new_n205), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n268), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n263), .A2(KEYINPUT16), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT70), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n272), .B2(new_n274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT16), .ZN(new_n279));
  INV_X1    g0079(.A(new_n270), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n203), .B1(new_n257), .B2(new_n259), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n271), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  OAI211_X1 g0090(.A(G223), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(G226), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G87), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  OAI211_X1 g0095(.A(G1), .B(G13), .C1(new_n251), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n287), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n285), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G232), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G200), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n298), .A2(G190), .A3(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n275), .B2(new_n276), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n272), .A2(new_n274), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT70), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(KEYINPUT71), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n253), .A2(G1), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G13), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n306), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT8), .B(G58), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n284), .A2(G20), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(KEYINPUT76), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT76), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n314), .B2(new_n311), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n313), .A2(new_n320), .B1(new_n315), .B2(new_n312), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n283), .A2(new_n303), .A3(new_n304), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT17), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n289), .A2(new_n290), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT7), .B1(new_n325), .B2(new_n253), .ZN(new_n326));
  OAI21_X1  g0126(.A(G68), .B1(new_n326), .B2(new_n261), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n270), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n277), .B1(new_n328), .B2(new_n279), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n321), .B1(new_n329), .B2(new_n271), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n303), .A4(new_n304), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n283), .A2(new_n322), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n294), .A2(new_n297), .ZN(new_n335));
  INV_X1    g0135(.A(new_n287), .ZN(new_n336));
  AND4_X1   g0136(.A1(G179), .A2(new_n335), .A3(new_n301), .A4(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n298), .B2(new_n301), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(KEYINPUT18), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT18), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n337), .A2(new_n339), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n330), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n333), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n252), .A2(new_n254), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n221), .A2(new_n288), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n348), .B(new_n349), .C1(G232), .C2(new_n288), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n297), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n299), .A2(new_n215), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n336), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT13), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n287), .B1(new_n352), .B2(new_n297), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(new_n355), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT73), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(G169), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n359), .B1(new_n358), .B2(new_n355), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n296), .B1(new_n350), .B2(new_n351), .ZN(new_n366));
  NOR4_X1   g0166(.A1(new_n366), .A2(KEYINPUT13), .A3(new_n287), .A4(new_n354), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n362), .B(G169), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n357), .A2(new_n360), .A3(G179), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n306), .A2(new_n310), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n251), .A2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G77), .B1(new_n269), .B2(G50), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n253), .B2(G68), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT11), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G13), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n316), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n203), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT12), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n278), .A2(new_n311), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G68), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n372), .A2(KEYINPUT11), .A3(new_n375), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n378), .A2(new_n382), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n371), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n365), .A2(new_n367), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n386), .B1(G190), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n361), .A2(G200), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n347), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G200), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT68), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n348), .A2(new_n288), .ZN(new_n395));
  INV_X1    g0195(.A(G222), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XOR2_X1   g0197(.A(KEYINPUT69), .B(G223), .Z(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(G1698), .A3(new_n348), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n325), .A2(G77), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n348), .A2(KEYINPUT68), .A3(G222), .A4(new_n288), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n397), .A2(new_n399), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n287), .B1(new_n402), .B2(new_n297), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n300), .A2(G226), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n393), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n312), .A2(G50), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n316), .A2(G50), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n372), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT72), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n373), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n269), .A2(G150), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(new_n206), .C2(new_n253), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n372), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n410), .B1(new_n372), .B2(new_n415), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n407), .B(new_n409), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n405), .B1(new_n419), .B2(KEYINPUT9), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT10), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n403), .A2(G190), .A3(new_n404), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT9), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT71), .B1(new_n308), .B2(new_n309), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n275), .A2(new_n276), .A3(new_n305), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n415), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT72), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n372), .A2(new_n410), .A3(new_n415), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n431), .A2(KEYINPUT9), .A3(new_n407), .A4(new_n409), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n402), .A2(new_n297), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(new_n336), .A3(new_n404), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G200), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n424), .A2(new_n432), .A3(new_n422), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT10), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n425), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n434), .A2(G179), .ZN(new_n439));
  AOI21_X1  g0239(.A(G169), .B1(new_n403), .B2(new_n404), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n439), .A2(new_n419), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n383), .A2(G77), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n380), .A2(new_n207), .ZN(new_n445));
  INV_X1    g0245(.A(new_n269), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n314), .A2(new_n446), .B1(new_n253), .B2(new_n207), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT15), .B(G87), .ZN(new_n448));
  INV_X1    g0248(.A(new_n373), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n278), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n348), .A2(G238), .A3(G1698), .ZN(new_n454));
  INV_X1    g0254(.A(G107), .ZN(new_n455));
  OAI221_X1 g0255(.A(new_n454), .B1(new_n455), .B2(new_n348), .C1(new_n395), .C2(new_n214), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n297), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n300), .A2(G244), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n457), .A2(G190), .A3(new_n336), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n336), .A3(new_n458), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n453), .B(new_n459), .C1(new_n461), .C2(new_n393), .ZN(new_n462));
  INV_X1    g0262(.A(G179), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n457), .A2(new_n463), .A3(new_n336), .A4(new_n458), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n452), .C1(new_n461), .C2(G169), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n392), .A2(new_n443), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n284), .B(G45), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(new_n286), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n470), .A2(new_n296), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G270), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT85), .A2(G303), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT85), .A2(G303), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(new_n252), .A3(new_n254), .A4(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(G264), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n477));
  OAI211_X1 g0277(.A(G257), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n479), .A2(new_n480), .A3(new_n297), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n479), .B2(new_n297), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n471), .B(new_n473), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n253), .C1(G33), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n210), .A2(G20), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n307), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n486), .A2(KEYINPUT20), .A3(new_n307), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n284), .A2(G33), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n312), .A2(G116), .A3(new_n492), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n490), .A2(new_n491), .B1(new_n493), .B2(new_n277), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n380), .A2(new_n210), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n338), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n483), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n483), .A2(G200), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n479), .A2(new_n297), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT86), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n479), .A2(new_n480), .A3(new_n297), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(G190), .A3(new_n471), .A4(new_n473), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n494), .A2(new_n495), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n500), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n502), .A2(new_n503), .B1(G270), .B2(new_n472), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(new_n506), .A3(G179), .A4(new_n471), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n483), .A2(new_n496), .A3(KEYINPUT21), .ZN(new_n511));
  AND4_X1   g0311(.A1(new_n499), .A2(new_n508), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT19), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n253), .B1(new_n351), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  INV_X1    g0315(.A(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n348), .A2(new_n253), .A3(G68), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n514), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n513), .B1(new_n449), .B2(new_n485), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n519), .A2(new_n520), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n278), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n380), .A2(new_n448), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n306), .A2(new_n310), .A3(new_n312), .A4(new_n492), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(new_n516), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n306), .A2(new_n310), .A3(new_n312), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(KEYINPUT84), .A3(G87), .A4(new_n492), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n527), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(G244), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n534));
  OAI211_X1 g0334(.A(G238), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n297), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n284), .A2(G45), .A3(G274), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n284), .A2(G45), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n296), .A2(G250), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  INV_X1    g0344(.A(new_n541), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n537), .B2(new_n297), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n546), .B2(new_n539), .ZN(new_n547));
  OAI21_X1  g0347(.A(G190), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n544), .A3(new_n539), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(G200), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n533), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n463), .B1(new_n543), .B2(new_n547), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n525), .B(new_n526), .C1(new_n448), .C2(new_n529), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n338), .A3(new_n550), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n380), .A2(new_n485), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n529), .B2(new_n485), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  AND2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n515), .ZN(new_n563));
  NAND2_X1  g0363(.A1(KEYINPUT6), .A2(G97), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT77), .B1(new_n564), .B2(G107), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT77), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n566), .A2(new_n455), .A3(KEYINPUT6), .A4(G97), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(G20), .B1(G77), .B2(new_n269), .ZN(new_n569));
  OAI21_X1  g0369(.A(G107), .B1(new_n326), .B2(new_n261), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n277), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT78), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI211_X1 g0373(.A(KEYINPUT78), .B(new_n277), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n560), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n348), .A2(G244), .A3(new_n288), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT79), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n348), .A2(G250), .A3(G1698), .ZN(new_n581));
  INV_X1    g0381(.A(new_n579), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n348), .A2(new_n582), .A3(G244), .A4(new_n288), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n580), .A2(new_n484), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n297), .B1(G257), .B2(new_n472), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n585), .A2(G179), .A3(new_n471), .ZN(new_n586));
  INV_X1    g0386(.A(new_n471), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n472), .A2(G257), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n587), .B(new_n588), .C1(new_n297), .C2(new_n584), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n589), .B2(new_n338), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT81), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n591), .B(new_n560), .C1(new_n573), .C2(new_n574), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n576), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n568), .A2(G20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n269), .A2(G77), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n455), .B1(new_n257), .B2(new_n259), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n278), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT78), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n571), .A2(new_n572), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n559), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT80), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n589), .A2(new_n602), .A3(G190), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n585), .A2(new_n471), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT80), .B1(new_n604), .B2(G200), .ZN(new_n605));
  INV_X1    g0405(.A(G190), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n601), .B(new_n603), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n512), .A2(new_n557), .A3(new_n593), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n348), .A2(G257), .A3(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n348), .A2(G250), .A3(new_n288), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G294), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n297), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT90), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n472), .A2(G264), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(KEYINPUT90), .A3(new_n297), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n471), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G169), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n614), .A2(new_n617), .A3(new_n471), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G179), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n380), .A2(new_n455), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT25), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n529), .B2(new_n455), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n626), .B(KEYINPUT88), .C1(new_n529), .C2(new_n455), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n253), .A2(G107), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT23), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n536), .A2(G20), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT87), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n253), .B(G87), .C1(new_n289), .C2(new_n290), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(KEYINPUT22), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(KEYINPUT22), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n633), .B(new_n635), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT24), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n636), .B(KEYINPUT22), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(KEYINPUT24), .A3(new_n633), .A4(new_n635), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n278), .A3(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n631), .A2(KEYINPUT89), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT89), .B1(new_n631), .B2(new_n644), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n623), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n471), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n614), .A2(new_n617), .A3(new_n471), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n648), .A2(new_n606), .B1(new_n393), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n306), .A2(new_n310), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n651), .A2(G107), .A3(new_n312), .A4(new_n492), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT88), .B1(new_n652), .B2(new_n626), .ZN(new_n653));
  INV_X1    g0453(.A(new_n630), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n644), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n609), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n467), .A2(new_n658), .ZN(G372));
  AND2_X1   g0459(.A1(new_n389), .A2(new_n390), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n387), .B1(new_n660), .B2(new_n465), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n333), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT93), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT18), .B1(new_n334), .B2(new_n340), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n330), .A2(new_n342), .A3(new_n343), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n341), .A2(new_n344), .A3(KEYINPUT93), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n441), .B1(new_n669), .B2(new_n438), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n542), .A2(new_n338), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n553), .A2(new_n554), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n599), .A2(new_n600), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n591), .B1(new_n674), .B2(new_n560), .ZN(new_n675));
  INV_X1    g0475(.A(new_n592), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g0477(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n678));
  NAND4_X1  g0478(.A1(new_n557), .A2(new_n677), .A3(new_n590), .A4(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n542), .A2(G200), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n533), .A2(new_n548), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n672), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n590), .A2(new_n575), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n673), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n593), .A2(new_n608), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n650), .A2(new_n655), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n683), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n620), .A2(new_n622), .B1(new_n631), .B2(new_n644), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n499), .A2(new_n510), .A3(new_n511), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT91), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n623), .A2(new_n655), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT91), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n510), .A2(new_n511), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n693), .A2(new_n694), .A3(new_n499), .A4(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n687), .A2(new_n689), .A3(new_n692), .A4(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n686), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n467), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n670), .B1(new_n698), .B2(new_n699), .ZN(G369));
  NAND3_X1  g0500(.A1(new_n284), .A2(new_n253), .A3(G13), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g0504(.A(KEYINPUT94), .B(G343), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n691), .A2(new_n506), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n508), .A2(new_n499), .A3(new_n510), .A4(new_n511), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n506), .B2(new_n707), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n710), .B2(KEYINPUT95), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(KEYINPUT95), .B2(new_n708), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT89), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n655), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n631), .A2(KEYINPUT89), .A3(new_n644), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n688), .B1(new_n718), .B2(new_n623), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n707), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n623), .A3(new_n707), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n714), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n707), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n691), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n657), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n690), .B2(new_n726), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n729), .ZN(G399));
  INV_X1    g0530(.A(new_n226), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n517), .A2(G116), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(G1), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n232), .B2(new_n733), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT28), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n647), .A2(new_n499), .A3(new_n695), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT96), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n593), .A2(new_n608), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n593), .B2(new_n608), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n738), .B(new_n689), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n683), .A2(new_n684), .A3(new_n680), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n552), .A2(new_n556), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n593), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n678), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n742), .B(new_n672), .C1(new_n743), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n726), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT29), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n707), .B1(new_n686), .B2(new_n697), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n709), .A2(new_n744), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n719), .A2(new_n687), .A3(new_n753), .A4(new_n726), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n509), .A2(new_n585), .A3(G179), .A4(new_n471), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n621), .B1(new_n543), .B2(new_n547), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(G179), .B1(new_n585), .B2(new_n471), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(new_n649), .A3(new_n542), .A4(new_n483), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n483), .A2(new_n463), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n649), .B1(new_n549), .B2(new_n550), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n761), .A2(new_n762), .A3(KEYINPUT30), .A4(new_n585), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n758), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n707), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n764), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n754), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G330), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n749), .A2(new_n752), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n737), .B1(new_n772), .B2(G1), .ZN(G364));
  NAND3_X1  g0573(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n606), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n348), .B1(new_n775), .B2(G326), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(G317), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n463), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n253), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n776), .B(new_n781), .C1(new_n782), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n393), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G179), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G283), .A2(new_n789), .B1(new_n792), .B2(G329), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n253), .A2(new_n606), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n783), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G322), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n794), .A2(new_n787), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n793), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n253), .B1(new_n790), .B2(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n786), .B(new_n800), .C1(G294), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n785), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G77), .ZN(new_n805));
  INV_X1    g0605(.A(new_n799), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G87), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n789), .A2(G107), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n325), .B1(new_n777), .B2(G68), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n805), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OR3_X1    g0611(.A1(new_n791), .A2(KEYINPUT32), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n775), .A2(G50), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n802), .A2(G97), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT32), .B1(new_n791), .B2(new_n811), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n810), .B(new_n816), .C1(G58), .C2(new_n796), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n803), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT100), .Z(new_n819));
  AOI21_X1  g0619(.A(new_n274), .B1(G20), .B2(new_n338), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n253), .A2(G13), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT98), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G45), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n824), .A2(G1), .A3(new_n733), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n232), .A2(G45), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n245), .A2(G45), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n827), .B2(KEYINPUT99), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n731), .A2(new_n348), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(KEYINPUT99), .C2(new_n827), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n731), .A2(new_n325), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G355), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n830), .B(new_n832), .C1(G116), .C2(new_n226), .ZN(new_n833));
  NOR2_X1   g0633(.A1(G13), .A2(G33), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(G20), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n820), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n825), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n836), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n821), .B(new_n838), .C1(new_n712), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n713), .A2(new_n825), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n712), .A2(G330), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(G396));
  NAND2_X1  g0643(.A1(new_n452), .A2(new_n707), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n462), .A2(new_n465), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT102), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n462), .A2(new_n465), .A3(KEYINPUT102), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n750), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n465), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n707), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT103), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n851), .B1(new_n750), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n770), .ZN(new_n857));
  INV_X1    g0657(.A(new_n770), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n858), .B(new_n851), .C1(new_n750), .C2(new_n855), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n857), .A2(new_n825), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n825), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n804), .A2(G159), .B1(G137), .B2(new_n775), .ZN(new_n862));
  INV_X1    g0662(.A(G143), .ZN(new_n863));
  INV_X1    g0663(.A(G150), .ZN(new_n864));
  INV_X1    g0664(.A(new_n777), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n862), .B1(new_n863), .B2(new_n795), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT34), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n348), .B1(new_n791), .B2(new_n868), .C1(new_n220), .C2(new_n799), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(G58), .B2(new_n802), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n867), .B(new_n870), .C1(new_n203), .C2(new_n788), .ZN(new_n871));
  AOI22_X1  g0671(.A1(G107), .A2(new_n806), .B1(new_n804), .B2(G116), .ZN(new_n872));
  INV_X1    g0672(.A(G294), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n872), .B1(new_n873), .B2(new_n795), .C1(new_n782), .C2(new_n791), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n788), .A2(new_n516), .ZN(new_n875));
  INV_X1    g0675(.A(new_n775), .ZN(new_n876));
  INV_X1    g0676(.A(G283), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n814), .B1(new_n876), .B2(new_n798), .C1(new_n877), .C2(new_n865), .ZN(new_n878));
  OR3_X1    g0678(.A1(new_n874), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n871), .B1(new_n348), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n820), .A2(new_n834), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT101), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n880), .A2(new_n820), .B1(new_n207), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n861), .B(new_n884), .C1(new_n854), .C2(new_n835), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n860), .A2(new_n885), .ZN(G384));
  NAND2_X1  g0686(.A1(new_n386), .A2(new_n707), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n387), .A2(new_n391), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n386), .B(new_n707), .C1(new_n660), .C2(new_n371), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(new_n889), .B1(new_n849), .B2(new_n853), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n754), .A2(new_n768), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT104), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n765), .B2(new_n766), .ZN(new_n893));
  AOI211_X1 g0693(.A(KEYINPUT104), .B(KEYINPUT31), .C1(new_n764), .C2(new_n707), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n890), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n334), .A2(new_n340), .ZN(new_n898));
  INV_X1    g0698(.A(new_n704), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n334), .A2(new_n899), .ZN(new_n900));
  AND4_X1   g0700(.A1(new_n897), .A2(new_n898), .A3(new_n900), .A4(new_n323), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n271), .A2(new_n372), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT16), .B1(new_n263), .B2(new_n270), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n904), .A2(new_n321), .B1(new_n340), .B2(new_n899), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n897), .B1(new_n905), .B2(new_n323), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  INV_X1    g0708(.A(new_n903), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n372), .A3(new_n271), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n322), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n899), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n333), .B2(new_n345), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n900), .A2(KEYINPUT93), .A3(new_n323), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n898), .A2(new_n900), .A3(new_n323), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n283), .A2(new_n304), .A3(new_n322), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(new_n303), .B1(new_n334), .B2(new_n899), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n920), .A2(new_n663), .A3(KEYINPUT37), .A4(new_n898), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n666), .A2(new_n667), .B1(new_n324), .B2(new_n332), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n918), .B(new_n921), .C1(new_n922), .C2(new_n900), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n914), .B1(new_n923), .B2(new_n908), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT40), .B1(new_n896), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n888), .A2(new_n889), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n854), .ZN(new_n927));
  INV_X1    g0727(.A(new_n768), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n658), .B2(new_n726), .ZN(new_n929));
  INV_X1    g0729(.A(new_n893), .ZN(new_n930));
  INV_X1    g0730(.A(new_n894), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n927), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n908), .B1(new_n907), .B2(new_n913), .ZN(new_n934));
  INV_X1    g0734(.A(new_n913), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n910), .A2(new_n322), .B1(new_n343), .B2(new_n704), .ZN(new_n936));
  INV_X1    g0736(.A(new_n323), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT37), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n898), .A2(new_n900), .A3(new_n897), .A4(new_n323), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n935), .A2(KEYINPUT38), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT40), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n925), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n754), .B(new_n768), .C1(new_n893), .C2(new_n894), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n467), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(G330), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n465), .A2(new_n707), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n750), .B2(new_n850), .ZN(new_n950));
  INV_X1    g0750(.A(new_n926), .ZN(new_n951));
  INV_X1    g0751(.A(new_n934), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n914), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n387), .A2(new_n707), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n900), .B1(new_n668), .B2(new_n333), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n918), .A2(new_n921), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n908), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT39), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n960), .A3(new_n941), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT39), .B1(new_n952), .B2(new_n914), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n668), .A2(new_n899), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n954), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n948), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n751), .B1(new_n747), .B2(new_n726), .ZN(new_n967));
  INV_X1    g0767(.A(new_n752), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n467), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n670), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n966), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n284), .B2(new_n823), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n210), .B1(new_n568), .B2(KEYINPUT35), .ZN(new_n973));
  INV_X1    g0773(.A(new_n231), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(KEYINPUT35), .C2(new_n568), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT36), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n265), .A2(new_n267), .A3(G77), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n232), .A2(new_n977), .B1(G50), .B2(new_n203), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(G1), .A3(new_n379), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n972), .A2(new_n976), .A3(new_n979), .ZN(G367));
  OR2_X1    g0780(.A1(new_n533), .A2(new_n726), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n672), .A3(new_n682), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT105), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT105), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(new_n672), .C2(new_n981), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(new_n839), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n348), .B1(new_n865), .B2(new_n811), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n789), .A2(G77), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n220), .B2(new_n785), .C1(new_n202), .C2(new_n799), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n802), .A2(G68), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n864), .B2(new_n795), .C1(new_n876), .C2(new_n863), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT109), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n987), .B(new_n989), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(G137), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n993), .B1(new_n992), .B2(new_n991), .C1(new_n994), .C2(new_n791), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT46), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n799), .A2(new_n996), .A3(new_n210), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n799), .B2(new_n210), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n455), .B2(new_n801), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(G311), .C2(new_n775), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n325), .B1(new_n865), .B2(new_n873), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n485), .A2(new_n788), .B1(new_n785), .B2(new_n877), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(G317), .C2(new_n792), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n474), .A2(new_n475), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1000), .B(new_n1003), .C1(new_n1004), .C2(new_n795), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n995), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n825), .B1(new_n1007), .B2(new_n820), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n829), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n837), .B1(new_n226), .B2(new_n448), .C1(new_n241), .C2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n986), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT106), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n740), .A2(new_n741), .B1(new_n601), .B2(new_n726), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n684), .A2(new_n726), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1012), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n728), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT42), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n647), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n593), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n726), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n728), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT42), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT107), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1027), .B(KEYINPUT42), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1033), .A2(KEYINPUT107), .A3(new_n1025), .A4(new_n1024), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1025), .B1(new_n1033), .B2(new_n1024), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n725), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n1019), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1041), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1035), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n732), .B(KEYINPUT41), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT44), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1019), .B2(new_n729), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n729), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1017), .A2(KEYINPUT44), .A3(new_n1049), .A4(new_n1018), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1018), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n729), .B1(new_n1052), .B2(new_n1016), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1019), .A2(KEYINPUT45), .A3(new_n729), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n1040), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1051), .A2(new_n1057), .A3(new_n725), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n723), .A2(new_n727), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1061), .A2(new_n713), .A3(new_n1026), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n713), .B1(new_n1026), .B2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1059), .A2(new_n772), .A3(new_n1060), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1046), .B1(new_n1066), .B2(new_n772), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n824), .A2(G1), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1042), .B(new_n1044), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1069), .A2(KEYINPUT108), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT108), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1035), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1043), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1068), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n771), .B(KEYINPUT97), .Z(new_n1076));
  AND3_X1   g0876(.A1(new_n1051), .A2(new_n1057), .A3(new_n725), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n725), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1076), .B1(new_n1079), .B2(new_n1065), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1075), .B1(new_n1080), .B2(new_n1046), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1071), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1011), .B1(new_n1070), .B2(new_n1082), .ZN(G387));
  INV_X1    g0883(.A(G326), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n325), .B1(new_n791), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1004), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n804), .A2(new_n1086), .B1(G322), .B2(new_n775), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n782), .B2(new_n865), .C1(new_n778), .C2(new_n795), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT48), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n799), .A2(new_n873), .B1(new_n801), .B2(new_n877), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT111), .Z(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT49), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1085), .B(new_n1095), .C1(G116), .C2(new_n789), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n799), .A2(new_n207), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G150), .B2(new_n792), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n220), .B2(new_n795), .C1(new_n203), .C2(new_n785), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n788), .A2(new_n485), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n801), .A2(new_n448), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n775), .B2(G159), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n314), .B2(new_n865), .ZN(new_n1103));
  NOR4_X1   g0903(.A1(new_n1099), .A2(new_n325), .A3(new_n1100), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n820), .B1(new_n1096), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n238), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1009), .B1(new_n1106), .B2(G45), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n734), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n831), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n315), .A2(new_n220), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n734), .B1(new_n203), .B2(new_n207), .C1(new_n1110), .C2(KEYINPUT50), .ZN(new_n1111));
  AOI211_X1 g0911(.A(G45), .B(new_n1111), .C1(KEYINPUT50), .C2(new_n1110), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1109), .A2(new_n1112), .B1(G107), .B2(new_n226), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n825), .B1(new_n1113), .B2(new_n837), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT110), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1105), .B(new_n1115), .C1(new_n724), .C2(new_n839), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n772), .B(new_n1065), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1116), .B1(new_n1075), .B2(new_n1064), .C1(new_n1117), .C2(new_n733), .ZN(G393));
  OAI22_X1  g0918(.A1(new_n1076), .A2(new_n1064), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n732), .A3(new_n1066), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1079), .A2(new_n1068), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n837), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n226), .A2(new_n485), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(new_n248), .C2(new_n829), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G68), .A2(new_n806), .B1(new_n792), .B2(G143), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n314), .B2(new_n785), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G77), .B2(new_n802), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n325), .B(new_n875), .C1(G50), .C2(new_n777), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n876), .A2(new_n864), .B1(new_n795), .B2(new_n811), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT51), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n808), .B1(new_n865), .B2(new_n1004), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n348), .B(new_n1132), .C1(G116), .C2(new_n802), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n876), .A2(new_n778), .B1(new_n795), .B2(new_n782), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT52), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G283), .A2(new_n806), .B1(new_n792), .B2(G322), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n785), .A2(new_n873), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1131), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n825), .B(new_n1124), .C1(new_n1139), .C2(new_n820), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT114), .Z(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1019), .B2(new_n839), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1120), .A2(new_n1121), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(G390));
  INV_X1    g0944(.A(new_n949), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n851), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n955), .B1(new_n1146), .B2(new_n926), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n961), .A2(new_n962), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n747), .A2(new_n726), .A3(new_n850), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n951), .B1(new_n1149), .B2(new_n1145), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n924), .A2(new_n955), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1147), .A2(new_n1148), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(G330), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n896), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT115), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1153), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n858), .A2(new_n854), .A3(new_n926), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT115), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1153), .A2(new_n1161), .A3(new_n1155), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1157), .A2(new_n1160), .A3(new_n1068), .A4(new_n1162), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n788), .A2(new_n203), .B1(new_n791), .B2(new_n873), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT117), .Z(new_n1165));
  OAI22_X1  g0965(.A1(new_n795), .A2(new_n210), .B1(new_n801), .B2(new_n207), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT118), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n325), .B1(new_n785), .B2(new_n485), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n807), .B1(new_n876), .B2(new_n877), .C1(new_n455), .C2(new_n865), .ZN(new_n1169));
  OR4_X1    g0969(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n348), .B1(new_n876), .B2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n865), .A2(new_n994), .B1(new_n801), .B2(new_n811), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(G50), .C2(new_n789), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT54), .B(G143), .Z(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1176), .A2(new_n785), .B1(new_n868), .B2(new_n795), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT53), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n799), .B2(new_n864), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n806), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(G125), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1174), .B(new_n1181), .C1(new_n1182), .C2(new_n791), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1170), .A2(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1184), .A2(new_n820), .B1(new_n314), .B2(new_n883), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n861), .B(new_n1185), .C1(new_n1148), .C2(new_n835), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT116), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n946), .B2(new_n1154), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n945), .A2(new_n467), .A3(KEYINPUT116), .A4(G330), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n969), .A3(new_n670), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n926), .B1(new_n858), .B2(new_n854), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1146), .B1(new_n1192), .B2(new_n1155), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n855), .A2(G330), .A3(new_n945), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n951), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1195), .A2(new_n1159), .A3(new_n1145), .A4(new_n1149), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1191), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n1160), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1157), .A2(new_n1160), .A3(new_n1162), .A4(new_n1197), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n732), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1163), .B(new_n1186), .C1(new_n1199), .C2(new_n1201), .ZN(G378));
  INV_X1    g1002(.A(KEYINPUT121), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT120), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n419), .A2(new_n704), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n443), .A2(KEYINPUT119), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT119), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n438), .A2(new_n1210), .A3(new_n442), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1208), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1210), .B1(new_n438), .B2(new_n442), .ZN(new_n1213));
  AOI211_X1 g1013(.A(KEYINPUT119), .B(new_n441), .C1(new_n425), .C2(new_n437), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n1207), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1206), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1209), .A2(new_n1211), .A3(new_n1208), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1207), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1205), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1204), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n341), .A2(new_n344), .A3(KEYINPUT93), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT93), .B1(new_n341), .B2(new_n344), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n333), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n900), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n898), .A2(new_n920), .B1(new_n915), .B2(KEYINPUT37), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n900), .A2(new_n323), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n330), .A2(new_n343), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1227), .A2(KEYINPUT93), .A3(new_n897), .A4(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT38), .B1(new_n1225), .B2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n945), .B(new_n890), .C1(new_n1231), .C2(new_n914), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1232), .A2(KEYINPUT40), .B1(new_n933), .B2(new_n942), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1220), .B1(new_n1233), .B2(new_n1154), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1217), .A2(new_n1218), .A3(new_n1205), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1205), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1236));
  OAI21_X1  g1036(.A(KEYINPUT120), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n944), .A2(new_n1237), .A3(G330), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n965), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1203), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1234), .A2(new_n965), .A3(new_n1238), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT122), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT122), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1234), .A2(new_n965), .A3(new_n1238), .A4(new_n1244), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1241), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1243), .A2(new_n1245), .B1(new_n1247), .B2(KEYINPUT121), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1191), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1200), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT57), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1247), .B2(new_n1242), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n732), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n865), .A2(new_n868), .B1(new_n876), .B2(new_n1182), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G128), .A2(new_n796), .B1(new_n804), .B2(G137), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n799), .B2(new_n1176), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(G150), .C2(new_n802), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT59), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G41), .B1(new_n792), .B2(G124), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G33), .B1(new_n789), .B2(G159), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n220), .B1(new_n289), .B2(G41), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n990), .B1(new_n876), .B2(new_n210), .C1(new_n485), .C2(new_n865), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(new_n1267), .A2(G41), .A3(new_n348), .A4(new_n1097), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n448), .A2(new_n785), .B1(new_n788), .B2(new_n202), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(G107), .B2(new_n796), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1268), .B(new_n1270), .C1(new_n877), .C2(new_n791), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT58), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1265), .A2(new_n1266), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n825), .B1(new_n1273), .B2(new_n820), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1274), .B1(G50), .B2(new_n882), .C1(new_n1275), .C2(new_n835), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1249), .B2(new_n1068), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1257), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(G375));
  AOI22_X1  g1081(.A1(new_n802), .A2(G50), .B1(new_n1175), .B2(new_n777), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1282), .B(new_n348), .C1(new_n868), .C2(new_n876), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(G137), .A2(new_n796), .B1(new_n806), .B2(G159), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1284), .B1(new_n1171), .B2(new_n791), .C1(new_n864), .C2(new_n785), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1283), .B(new_n1285), .C1(G58), .C2(new_n789), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(G283), .A2(new_n796), .B1(new_n792), .B2(G303), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1287), .B1(new_n485), .B2(new_n799), .C1(new_n455), .C2(new_n785), .ZN(new_n1288));
  OAI221_X1 g1088(.A(new_n988), .B1(new_n876), .B2(new_n873), .C1(new_n210), .C2(new_n865), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1288), .A2(new_n1101), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1286), .B1(new_n325), .B2(new_n1290), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(KEYINPUT123), .Z(new_n1292));
  AOI21_X1  g1092(.A(new_n825), .B1(new_n1292), .B2(new_n820), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n1293), .B1(G68), .B2(new_n882), .C1(new_n926), .C2(new_n835), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1196), .A2(new_n1193), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1296), .B2(new_n1075), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1046), .B1(new_n1296), .B2(new_n1191), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1250), .A2(new_n1295), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(G381));
  OR4_X1    g1101(.A1(G396), .A2(G393), .A3(G390), .A4(G384), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1163), .A2(new_n1186), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1198), .A2(new_n1160), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1299), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1201), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1303), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1280), .A2(new_n1307), .ZN(new_n1308));
  OR4_X1    g1108(.A1(G387), .A2(new_n1302), .A3(new_n1308), .A4(G381), .ZN(G407));
  OAI211_X1 g1109(.A(G407), .B(G213), .C1(new_n705), .C2(new_n1308), .ZN(G409));
  XNOR2_X1  g1110(.A(G393), .B(G396), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1069), .A2(KEYINPUT108), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1074), .A2(new_n1081), .A3(new_n1071), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G390), .B1(new_n1314), .B2(new_n1011), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1011), .ZN(new_n1316));
  AOI211_X1 g1116(.A(new_n1316), .B(new_n1143), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1311), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G387), .A2(new_n1143), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1311), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1314), .A2(new_n1011), .A3(G390), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1318), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n706), .A2(G213), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G378), .B(new_n1278), .C1(new_n1252), .C2(new_n1256), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1241), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1241), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1251), .A2(new_n1045), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1247), .A2(new_n1242), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1068), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(new_n1276), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1307), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1325), .B1(new_n1326), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT60), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1337), .B1(new_n1250), .B2(new_n1295), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(new_n732), .A3(new_n1299), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1191), .A2(new_n1193), .A3(new_n1196), .A4(KEYINPUT60), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1341), .B(KEYINPUT125), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1297), .B1(new_n1340), .B2(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(KEYINPUT126), .B1(new_n1343), .B2(G384), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  INV_X1    g1145(.A(G384), .ZN(new_n1346));
  OR2_X1    g1146(.A1(new_n1341), .A2(KEYINPUT125), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1341), .A2(KEYINPUT125), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1339), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1345), .B(new_n1346), .C1(new_n1349), .C2(new_n1297), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1343), .A2(G384), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1344), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1352), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1336), .A2(KEYINPUT63), .A3(new_n1353), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1323), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT61), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT63), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1326), .A2(new_n1335), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT124), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1326), .A2(KEYINPUT124), .A3(new_n1335), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1360), .A2(new_n1324), .A3(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1325), .A2(G2897), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1352), .B(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1357), .B1(new_n1362), .B2(new_n1364), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1360), .A2(new_n1324), .A3(new_n1353), .A4(new_n1361), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  OAI211_X1 g1167(.A(new_n1355), .B(new_n1356), .C1(new_n1365), .C2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT62), .ZN(new_n1369));
  NOR2_X1   g1169(.A1(new_n1352), .A2(new_n1369), .ZN(new_n1370));
  AND2_X1   g1170(.A1(new_n1336), .A2(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1371), .B1(new_n1366), .B2(new_n1369), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1364), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1356), .B1(new_n1373), .B2(new_n1336), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1323), .B1(new_n1372), .B2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1368), .A2(new_n1375), .ZN(G405));
  NAND2_X1  g1176(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1377), .A2(new_n1253), .ZN(new_n1378));
  INV_X1    g1178(.A(new_n1256), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1180(.A(G378), .B1(new_n1380), .B2(new_n1278), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1326), .ZN(new_n1382));
  NOR2_X1   g1182(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1383));
  XNOR2_X1  g1183(.A(new_n1383), .B(new_n1352), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1384), .A2(KEYINPUT127), .A3(new_n1323), .ZN(new_n1385));
  XNOR2_X1  g1185(.A(new_n1383), .B(new_n1353), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1323), .A2(KEYINPUT127), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT127), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1318), .A2(new_n1322), .A3(new_n1388), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1386), .A2(new_n1387), .A3(new_n1389), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1385), .A2(new_n1390), .ZN(G402));
endmodule


