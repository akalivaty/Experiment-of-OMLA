//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909;
  NAND2_X1  g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT67), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G226gat), .A2(G233gat), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n214), .B(KEYINPUT68), .Z(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  AND2_X1   g016(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT28), .ZN(new_n221));
  AND2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(KEYINPUT26), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT28), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n221), .A2(new_n224), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n222), .A2(new_n230), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n217), .ZN(new_n239));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(KEYINPUT24), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n231), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n231), .A2(new_n237), .A3(new_n241), .A4(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT70), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n229), .A2(new_n244), .A3(new_n249), .A4(new_n246), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n216), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT69), .B(KEYINPUT29), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n216), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n213), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n215), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT29), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n248), .A2(new_n258), .A3(new_n250), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n259), .B2(new_n216), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n255), .B1(new_n260), .B2(new_n213), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n262));
  XNOR2_X1  g061(.A(G8gat), .B(G36gat), .ZN(new_n263));
  INV_X1    g062(.A(G64gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G92gat), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n261), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n262), .B1(new_n261), .B2(new_n266), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT30), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n261), .A2(KEYINPUT30), .A3(new_n266), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT71), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n261), .A2(new_n272), .A3(KEYINPUT30), .A4(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n261), .A2(new_n266), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n269), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT40), .ZN(new_n278));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279));
  AND2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G141gat), .B(G148gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n284), .B1(G155gat), .B2(G162gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G141gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G148gat), .ZN(new_n288));
  INV_X1    g087(.A(G148gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G141gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G155gat), .B(G162gat), .ZN(new_n292));
  INV_X1    g091(.A(G155gat), .ZN(new_n293));
  INV_X1    g092(.A(G162gat), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT2), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n286), .A2(new_n296), .A3(KEYINPUT73), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT73), .B1(new_n286), .B2(new_n296), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT3), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n286), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n286), .A2(new_n296), .A3(KEYINPUT74), .A4(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n306));
  XNOR2_X1  g105(.A(G127gat), .B(G134gat), .ZN(new_n307));
  INV_X1    g106(.A(G113gat), .ZN(new_n308));
  INV_X1    g107(.A(G120gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT65), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G120gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n309), .A2(G113gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n306), .B(new_n307), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n307), .ZN(new_n316));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(KEYINPUT1), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n299), .A2(new_n305), .A3(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n315), .A2(new_n318), .A3(new_n286), .A4(new_n296), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT4), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n286), .A2(new_n296), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n318), .A4(new_n315), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n279), .B1(new_n320), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n297), .A2(new_n298), .ZN(new_n329));
  INV_X1    g128(.A(new_n319), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n279), .ZN(new_n332));
  INV_X1    g131(.A(new_n321), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT39), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n328), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n327), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(new_n335), .A3(new_n332), .ZN(new_n338));
  XOR2_X1   g137(.A(G1gat), .B(G29gat), .Z(new_n339));
  XNOR2_X1  g138(.A(G57gat), .B(G85gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n278), .B1(new_n336), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT81), .B(new_n278), .C1(new_n336), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n321), .A2(new_n332), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n320), .A2(new_n350), .A3(new_n327), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n332), .B1(new_n331), .B2(new_n333), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT5), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n320), .A2(new_n327), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n343), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OR3_X1    g157(.A1(new_n328), .A2(new_n334), .A3(new_n335), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n328), .B2(new_n335), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(KEYINPUT40), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n349), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT82), .B1(new_n277), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT31), .B(G50gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n207), .A2(KEYINPUT78), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n204), .B(new_n367), .C1(new_n205), .C2(new_n206), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n209), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n211), .A2(KEYINPUT78), .A3(new_n207), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n252), .A3(new_n370), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n371), .A2(KEYINPUT79), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT3), .B1(new_n371), .B2(KEYINPUT79), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n324), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n213), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n305), .B2(new_n252), .ZN(new_n378));
  OR3_X1    g177(.A1(new_n374), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n213), .A2(KEYINPUT80), .A3(KEYINPUT29), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT80), .B1(new_n213), .B2(KEYINPUT29), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n329), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n376), .B1(new_n383), .B2(new_n378), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n365), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n384), .A3(new_n365), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  INV_X1    g187(.A(G22gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n390), .ZN(new_n392));
  INV_X1    g191(.A(new_n387), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n385), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n259), .A2(new_n216), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n213), .B1(new_n396), .B2(new_n256), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n248), .A2(new_n250), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n215), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n377), .B1(new_n399), .B2(new_n253), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n266), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT72), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n261), .A2(new_n262), .A3(new_n266), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n405), .A2(new_n275), .A3(new_n271), .A4(new_n273), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n343), .B1(new_n353), .B2(new_n355), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n347), .B2(new_n348), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .A4(new_n361), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT37), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n255), .B(new_n411), .C1(new_n260), .C2(new_n213), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n377), .B1(new_n251), .B2(new_n254), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(KEYINPUT37), .C1(new_n260), .C2(new_n377), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT38), .B(new_n266), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n415), .A2(new_n268), .A3(new_n267), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT76), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n353), .A2(new_n343), .A3(new_n355), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n358), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT76), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n422), .A3(KEYINPUT6), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n418), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n261), .B(new_n411), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT38), .B1(new_n425), .B2(new_n266), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n416), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n363), .A2(new_n395), .A3(new_n410), .A4(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT77), .B1(new_n406), .B2(new_n424), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n267), .A2(new_n268), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n276), .B1(new_n430), .B2(new_n403), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n418), .A2(new_n421), .A3(new_n423), .ZN(new_n433));
  INV_X1    g232(.A(new_n274), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n395), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n247), .A2(new_n330), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n247), .A2(new_n330), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(G227gat), .A3(G233gat), .A4(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  INV_X1    g240(.A(G71gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G99gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT33), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(KEYINPUT32), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(KEYINPUT66), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n440), .A2(KEYINPUT32), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n444), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT66), .B1(new_n440), .B2(new_n447), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n446), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n438), .A2(new_n439), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT34), .ZN(new_n454));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n446), .B(new_n458), .C1(new_n450), .C2(new_n451), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n428), .A2(new_n437), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n431), .A2(new_n466), .A3(new_n433), .A4(new_n434), .ZN(new_n467));
  INV_X1    g266(.A(new_n462), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n395), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT83), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n406), .A2(new_n424), .A3(KEYINPUT35), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n462), .B1(new_n391), .B2(new_n394), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n429), .B2(new_n435), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n470), .B(new_n474), .C1(new_n475), .C2(new_n466), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT97), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT89), .B(G64gat), .ZN(new_n479));
  INV_X1    g278(.A(G57gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT88), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n479), .B(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G71gat), .A2(G78gat), .ZN(new_n483));
  OR2_X1    g282(.A1(G71gat), .A2(G78gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT9), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n480), .A2(new_n264), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n483), .B(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G85gat), .A2(G92gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT7), .ZN(new_n493));
  NAND2_X1  g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494));
  INV_X1    g293(.A(G85gat), .ZN(new_n495));
  INV_X1    g294(.A(G92gat), .ZN(new_n496));
  AOI22_X1  g295(.A1(KEYINPUT8), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(G99gat), .B(G106gat), .Z(new_n499));
  OAI21_X1  g298(.A(KEYINPUT91), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n499), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n493), .A4(new_n497), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n491), .B1(new_n504), .B2(KEYINPUT95), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n498), .A2(new_n499), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n504), .B(new_n506), .C1(new_n491), .C2(KEYINPUT95), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT10), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT10), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n507), .A2(new_n511), .A3(new_n491), .ZN(new_n512));
  INV_X1    g311(.A(G230gat), .ZN(new_n513));
  INV_X1    g312(.A(G233gat), .ZN(new_n514));
  OAI22_X1  g313(.A1(new_n510), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n508), .A2(new_n516), .A3(new_n509), .ZN(new_n517));
  XNOR2_X1  g316(.A(G176gat), .B(G204gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT96), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(G120gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(new_n289), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n515), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n515), .B2(new_n517), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n478), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n515), .A2(new_n517), .ZN(new_n525));
  INV_X1    g324(.A(new_n521), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n515), .A2(new_n517), .A3(new_n521), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT97), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT86), .B(G36gat), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G29gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  INV_X1    g332(.A(G43gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(G50gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n535), .B2(KEYINPUT87), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT14), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n537), .B(KEYINPUT85), .C1(G29gat), .C2(G36gat), .ZN(new_n538));
  OR3_X1    g337(.A1(KEYINPUT85), .A2(G29gat), .A3(G36gat), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT14), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n532), .A2(new_n536), .A3(new_n538), .A4(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n532), .A2(new_n538), .A3(new_n541), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n542), .B(new_n543), .C1(new_n544), .C2(KEYINPUT15), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n542), .A2(new_n543), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(KEYINPUT17), .A3(new_n546), .ZN(new_n550));
  XNOR2_X1  g349(.A(G15gat), .B(G22gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(G1gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(G1gat), .B2(new_n551), .ZN(new_n554));
  INV_X1    g353(.A(G8gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n547), .B(new_n558), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n560), .B(KEYINPUT13), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n557), .A2(KEYINPUT18), .A3(new_n559), .A4(new_n560), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(G169gat), .B(G197gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT12), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n563), .A2(new_n566), .A3(new_n567), .A4(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n530), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n477), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n556), .B1(new_n491), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G183gat), .ZN(new_n584));
  AND2_X1   g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587));
  INV_X1    g386(.A(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n586), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n491), .A2(new_n582), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n591), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT41), .ZN(new_n596));
  INV_X1    g395(.A(G232gat), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n596), .A2(new_n597), .A3(new_n514), .ZN(new_n598));
  INV_X1    g397(.A(new_n507), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n547), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n507), .B1(new_n546), .B2(new_n545), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n598), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n549), .A2(new_n507), .A3(new_n550), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT92), .ZN(new_n607));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608));
  INV_X1    g407(.A(KEYINPUT92), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n549), .A2(new_n609), .A3(new_n507), .A4(new_n550), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n605), .A2(new_n607), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT90), .B(G134gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G162gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n596), .B1(new_n597), .B2(new_n514), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n605), .A2(new_n607), .A3(new_n610), .ZN(new_n618));
  INV_X1    g417(.A(new_n608), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n613), .A2(new_n617), .B1(new_n620), .B2(new_n611), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n620), .A2(KEYINPUT94), .A3(new_n611), .A4(new_n617), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n595), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n581), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n424), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT98), .B(G1gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1324gat));
  NAND2_X1  g428(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n552), .A2(new_n555), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n626), .A2(new_n406), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n626), .ZN(new_n635));
  OAI21_X1  g434(.A(G8gat), .B1(new_n635), .B2(new_n277), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n633), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT99), .ZN(G1325gat));
  AOI21_X1  g438(.A(G15gat), .B1(new_n626), .B2(new_n468), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n626), .A2(G15gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n464), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(G1326gat));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n436), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n389), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n644), .B(new_n646), .ZN(G1327gat));
  INV_X1    g446(.A(new_n624), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n465), .B2(new_n476), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n595), .A2(new_n580), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n651), .A2(G29gat), .A3(new_n433), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT45), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n477), .A2(new_n624), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n649), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n650), .ZN(new_n661));
  OAI21_X1  g460(.A(G29gat), .B1(new_n661), .B2(new_n433), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n653), .A2(new_n662), .ZN(G1328gat));
  NOR3_X1   g462(.A1(new_n651), .A2(new_n531), .A3(new_n277), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT102), .Z(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT46), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT103), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(KEYINPUT46), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n531), .B1(new_n661), .B2(new_n277), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(KEYINPUT103), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .A4(new_n670), .ZN(G1329gat));
  NOR3_X1   g470(.A1(new_n651), .A2(G43gat), .A3(new_n462), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT104), .Z(new_n673));
  OAI21_X1  g472(.A(G43gat), .B1(new_n661), .B2(new_n464), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT47), .Z(G1330gat));
  OR3_X1    g475(.A1(new_n651), .A2(G50gat), .A3(new_n395), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n436), .A3(new_n650), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT106), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G50gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(KEYINPUT106), .ZN(new_n681));
  OAI211_X1 g480(.A(KEYINPUT48), .B(new_n677), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(G50gat), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT48), .B1(new_n683), .B2(new_n677), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(G1331gat));
  NAND4_X1  g487(.A1(new_n477), .A2(new_n625), .A3(new_n579), .A4(new_n530), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT107), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n424), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n406), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT108), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1333gat));
  XOR2_X1   g496(.A(new_n462), .B(KEYINPUT109), .Z(new_n698));
  AOI21_X1  g497(.A(G71gat), .B1(new_n690), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n464), .A2(new_n442), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n690), .B2(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g501(.A1(new_n690), .A2(new_n436), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G78gat), .ZN(G1335gat));
  INV_X1    g503(.A(new_n530), .ZN(new_n705));
  INV_X1    g504(.A(new_n595), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n578), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n477), .A2(new_n624), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT51), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n649), .A2(KEYINPUT51), .A3(new_n707), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n705), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(G85gat), .B1(new_n712), .B2(new_n424), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n656), .A2(new_n530), .A3(new_n659), .A4(new_n707), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(new_n495), .A3(new_n433), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(G1336gat));
  NAND3_X1  g515(.A1(new_n712), .A2(new_n496), .A3(new_n406), .ZN(new_n717));
  OAI21_X1  g516(.A(G92gat), .B1(new_n714), .B2(new_n277), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n705), .A2(G92gat), .A3(new_n277), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT110), .B1(new_n710), .B2(new_n711), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n708), .B2(new_n709), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n721), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n718), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT111), .B1(new_n726), .B2(KEYINPUT52), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n728), .B(new_n719), .C1(new_n725), .C2(new_n718), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n720), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT112), .B(new_n720), .C1(new_n727), .C2(new_n729), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1337gat));
  XOR2_X1   g533(.A(KEYINPUT113), .B(G99gat), .Z(new_n735));
  NAND3_X1  g534(.A1(new_n712), .A2(new_n468), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n714), .A2(new_n464), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n735), .ZN(G1338gat));
  OR2_X1    g537(.A1(new_n714), .A2(new_n395), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G106gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n710), .A2(new_n711), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n705), .A2(G106gat), .A3(new_n395), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT53), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n722), .A2(new_n724), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n742), .B(KEYINPUT114), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n745), .A2(new_n746), .B1(new_n739), .B2(G106gat), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(G1339gat));
  NOR2_X1   g548(.A1(new_n564), .A2(new_n565), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n560), .B1(new_n557), .B2(new_n559), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n573), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n577), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n530), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n508), .A2(new_n509), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n511), .ZN(new_n757));
  INV_X1    g556(.A(new_n512), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(new_n516), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n759), .A2(new_n515), .A3(KEYINPUT54), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n526), .B1(new_n515), .B2(KEYINPUT54), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n755), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n515), .A2(KEYINPUT54), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n515), .A3(KEYINPUT54), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT55), .A4(new_n526), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n762), .A2(new_n578), .A3(new_n528), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n754), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n648), .ZN(new_n768));
  INV_X1    g567(.A(new_n623), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n753), .B1(new_n769), .B2(new_n621), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n762), .A2(new_n528), .A3(new_n765), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT115), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n771), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n773), .A2(new_n624), .A3(new_n774), .A4(new_n753), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n768), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(new_n595), .ZN(new_n777));
  NOR4_X1   g576(.A1(new_n595), .A2(new_n624), .A3(new_n578), .A4(new_n530), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n395), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT116), .B(new_n395), .C1(new_n777), .C2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n406), .A2(new_n433), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n468), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(G113gat), .B1(new_n785), .B2(new_n579), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n779), .A2(new_n462), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n784), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n308), .A3(new_n578), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(G1340gat));
  OAI21_X1  g589(.A(G120gat), .B1(new_n785), .B2(new_n705), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n310), .A2(new_n312), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n792), .A3(new_n530), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT117), .Z(G1341gat));
  AOI21_X1  g594(.A(G127gat), .B1(new_n788), .B2(new_n706), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n785), .A2(new_n595), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g597(.A(G134gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n788), .A2(new_n799), .A3(new_n624), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT56), .Z(new_n801));
  OAI21_X1  g600(.A(G134gat), .B1(new_n785), .B2(new_n648), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1343gat));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n776), .A2(new_n804), .A3(new_n595), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n776), .B2(new_n595), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n778), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT57), .B1(new_n807), .B2(new_n395), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n464), .A2(new_n784), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n778), .B1(new_n776), .B2(new_n595), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n395), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n808), .A2(new_n578), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G141gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n811), .A2(new_n395), .A3(new_n809), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n579), .A2(G141gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT120), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n815), .B2(G141gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n816), .A2(new_n826), .A3(new_n819), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n821), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n816), .B2(new_n819), .ZN(new_n829));
  INV_X1    g628(.A(new_n819), .ZN(new_n830));
  AOI211_X1 g629(.A(KEYINPUT120), .B(new_n830), .C1(new_n815), .C2(G141gat), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n829), .A2(new_n831), .B1(new_n824), .B2(new_n823), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n828), .A2(new_n832), .ZN(G1344gat));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n808), .A2(new_n810), .A3(new_n814), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n834), .B(G148gat), .C1(new_n835), .C2(new_n705), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT57), .B1(new_n811), .B2(new_n395), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n773), .A2(new_n624), .A3(new_n753), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n706), .B1(new_n768), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n813), .B(new_n436), .C1(new_n839), .C2(new_n778), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n705), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n289), .B1(new_n842), .B2(new_n810), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n836), .B1(new_n843), .B2(new_n834), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n817), .A2(new_n289), .A3(new_n530), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1345gat));
  NOR3_X1   g645(.A1(new_n835), .A2(new_n293), .A3(new_n595), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n817), .A2(new_n706), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT121), .Z(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n293), .B2(new_n849), .ZN(G1346gat));
  OR2_X1    g649(.A1(new_n835), .A2(new_n648), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n817), .A2(new_n294), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n851), .A2(G162gat), .B1(new_n624), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g653(.A1(new_n277), .A2(new_n424), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n698), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT123), .Z(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n781), .B2(new_n782), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G169gat), .B1(new_n859), .B2(new_n579), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n787), .A2(new_n855), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n233), .A3(new_n578), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1348gat));
  AOI21_X1  g662(.A(G176gat), .B1(new_n861), .B2(new_n530), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n859), .A2(new_n705), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(G176gat), .ZN(G1349gat));
  AOI21_X1  g665(.A(new_n238), .B1(new_n858), .B2(new_n706), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n218), .A2(new_n219), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n595), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n867), .B1(new_n861), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT60), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n870), .B(new_n872), .ZN(G1350gat));
  AOI211_X1 g672(.A(new_n648), .B(new_n857), .C1(new_n781), .C2(new_n782), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(KEYINPUT125), .A3(new_n217), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n624), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(G190gat), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT126), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT125), .B1(new_n874), .B2(new_n217), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n876), .A3(G190gat), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(KEYINPUT61), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n861), .A2(new_n217), .A3(new_n624), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n886));
  OAI211_X1 g685(.A(KEYINPUT126), .B(new_n886), .C1(new_n875), .C2(new_n878), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(G1351gat));
  INV_X1    g687(.A(new_n841), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n464), .A2(new_n855), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G197gat), .B1(new_n892), .B2(new_n579), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n812), .A2(new_n891), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(G197gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n579), .B2(new_n895), .ZN(G1352gat));
  XOR2_X1   g695(.A(KEYINPUT127), .B(G204gat), .Z(new_n897));
  NOR3_X1   g696(.A1(new_n894), .A2(new_n705), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT62), .ZN(new_n899));
  INV_X1    g698(.A(new_n842), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(new_n890), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1353gat));
  NAND3_X1  g701(.A1(new_n889), .A2(new_n706), .A3(new_n891), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n903), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT63), .B1(new_n903), .B2(G211gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n706), .A2(new_n588), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n904), .A2(new_n905), .B1(new_n894), .B2(new_n906), .ZN(G1354gat));
  OAI21_X1  g706(.A(G218gat), .B1(new_n892), .B2(new_n648), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n894), .A2(G218gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n648), .B2(new_n909), .ZN(G1355gat));
endmodule


