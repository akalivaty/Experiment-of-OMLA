//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT84), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT29), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT74), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  OR2_X1    g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(KEYINPUT2), .ZN(new_n217));
  INV_X1    g016(.A(new_n215), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n211), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n214), .A2(new_n217), .B1(new_n221), .B2(new_n216), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT75), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n212), .B1(new_n210), .B2(new_n211), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n217), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G141gat), .B(G148gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n215), .B(new_n216), .C1(new_n228), .C2(KEYINPUT2), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n227), .A2(KEYINPUT75), .A3(new_n223), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n204), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n235));
  INV_X1    g034(.A(G211gat), .ZN(new_n236));
  INV_X1    g035(.A(G218gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n233), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n233), .B1(new_n238), .B2(new_n234), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n232), .A2(KEYINPUT77), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n204), .B1(new_n239), .B2(new_n240), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n222), .B1(new_n243), .B2(new_n223), .ZN(new_n244));
  INV_X1    g043(.A(G228gat), .ZN(new_n245));
  INV_X1    g044(.A(G233gat), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n223), .A3(new_n229), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT75), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT29), .B1(new_n251), .B2(new_n230), .ZN(new_n252));
  INV_X1    g051(.A(new_n241), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n242), .A2(new_n247), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n252), .A2(new_n253), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(KEYINPUT76), .A3(new_n204), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT3), .B1(new_n243), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n222), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n256), .A2(new_n260), .B1(new_n245), .B2(new_n246), .ZN(new_n261));
  INV_X1    g060(.A(G22gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G78gat), .B(G106gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT31), .ZN(new_n266));
  INV_X1    g065(.A(G50gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n261), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G22gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT78), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n274), .A3(new_n263), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(KEYINPUT78), .ZN(new_n276));
  AND4_X1   g075(.A1(KEYINPUT79), .A2(new_n275), .A3(new_n276), .A4(new_n269), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT78), .B1(new_n271), .B2(G22gat), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n268), .B1(new_n278), .B2(new_n263), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT79), .B1(new_n279), .B2(new_n276), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n273), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n251), .A2(new_n230), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G113gat), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G120gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT1), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G127gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G113gat), .B(G120gat), .ZN(new_n290));
  OAI21_X1  g089(.A(G127gat), .B1(new_n290), .B2(KEYINPUT1), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n291), .A3(G134gat), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n287), .A2(new_n288), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n290), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n227), .A2(new_n229), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n292), .A2(new_n296), .B1(new_n297), .B2(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n222), .A2(new_n296), .A3(new_n292), .ZN(new_n300));
  NAND2_X1  g099(.A1(G225gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n222), .A2(new_n296), .A3(KEYINPUT4), .A4(new_n292), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n299), .A2(new_n303), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT5), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n296), .A2(new_n292), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n297), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n300), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n311), .B2(new_n302), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n302), .A2(KEYINPUT5), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n299), .A2(new_n305), .A3(new_n306), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT0), .B(G57gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G85gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G1gat), .B(G29gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT6), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n313), .A2(new_n315), .A3(new_n320), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n316), .A2(KEYINPUT6), .A3(new_n321), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT64), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT64), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G183gat), .ZN(new_n336));
  INV_X1    g135(.A(G190gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G169gat), .ZN(new_n340));
  INV_X1    g139(.A(G176gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT23), .ZN(new_n342));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n341), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n339), .A2(new_n342), .A3(new_n343), .A4(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n350), .A3(new_n338), .ZN(new_n351));
  AND4_X1   g150(.A1(KEYINPUT25), .A2(new_n351), .A3(new_n342), .A4(new_n346), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n343), .B(KEYINPUT65), .Z(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n344), .A2(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(KEYINPUT26), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n343), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n336), .A2(KEYINPUT27), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT27), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G183gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT66), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n365));
  AOI21_X1  g164(.A(G190gat), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT28), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n363), .A2(new_n368), .A3(G190gat), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n331), .B(new_n359), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n356), .A3(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n347), .A2(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT67), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n361), .A2(G183gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n337), .B1(new_n375), .B2(KEYINPUT66), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n365), .B1(new_n360), .B2(new_n362), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n368), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n363), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(KEYINPUT28), .A3(new_n337), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n378), .A2(new_n380), .B1(G183gat), .B2(G190gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(KEYINPUT67), .A3(new_n359), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n372), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n356), .A2(KEYINPUT29), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n241), .B(new_n371), .C1(new_n383), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n355), .A2(new_n370), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n383), .A2(new_n356), .B1(new_n387), .B2(new_n384), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n386), .B(KEYINPUT72), .C1(new_n388), .C2(new_n241), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n370), .A2(new_n373), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT67), .B1(new_n381), .B2(new_n359), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n355), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n384), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n241), .A4(new_n371), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT73), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G8gat), .ZN(new_n398));
  INV_X1    g197(.A(G36gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n389), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT30), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n389), .B2(new_n395), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI211_X1 g203(.A(KEYINPUT30), .B(new_n400), .C1(new_n389), .C2(new_n395), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n327), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n309), .ZN(new_n409));
  INV_X1    g208(.A(new_n309), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n383), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT32), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT69), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT70), .B(G15gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G43gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n408), .ZN(new_n419));
  AOI211_X1 g218(.A(new_n309), .B(new_n372), .C1(new_n374), .C2(new_n382), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n374), .A2(new_n382), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n410), .B1(new_n421), .B2(new_n355), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n424));
  AOI21_X1  g223(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT69), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n426), .A3(KEYINPUT32), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n414), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n423), .B(KEYINPUT32), .C1(new_n424), .C2(new_n418), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n408), .A3(new_n411), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT34), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n432), .B1(new_n428), .B2(new_n429), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n281), .A2(new_n407), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n202), .A2(KEYINPUT84), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n203), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n203), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n428), .A2(new_n429), .ZN(new_n440));
  INV_X1    g239(.A(new_n432), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n275), .A2(new_n276), .A3(new_n269), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n279), .A2(KEYINPUT79), .A3(new_n276), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n449), .B2(new_n273), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n439), .B1(new_n450), .B2(new_n407), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n325), .A2(new_n326), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n389), .A2(new_n395), .ZN(new_n454));
  INV_X1    g253(.A(new_n400), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT37), .B1(new_n389), .B2(new_n395), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n253), .B(new_n371), .C1(new_n383), .C2(new_n385), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n458), .B(KEYINPUT37), .C1(new_n388), .C2(new_n253), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT38), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n400), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n452), .A2(new_n453), .A3(new_n456), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n325), .A2(new_n456), .A3(new_n326), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n457), .A2(new_n461), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT82), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n389), .A2(KEYINPUT37), .A3(new_n395), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n400), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT83), .ZN(new_n469));
  INV_X1    g268(.A(new_n457), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n471), .A3(new_n400), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n463), .A2(new_n466), .B1(KEYINPUT38), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT39), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n311), .A2(new_n302), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n299), .A2(new_n305), .A3(new_n306), .ZN(new_n477));
  AOI211_X1 g276(.A(new_n475), .B(new_n476), .C1(new_n302), .C2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n282), .A2(new_n298), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n305), .A2(new_n306), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n475), .B(new_n302), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n320), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT80), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n484), .A3(new_n320), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n478), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT81), .B1(new_n486), .B2(KEYINPUT40), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(KEYINPUT40), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n476), .B1(new_n477), .B2(new_n302), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT39), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n481), .A2(new_n484), .A3(new_n320), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n484), .B1(new_n481), .B2(new_n320), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT81), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n487), .A2(new_n322), .A3(new_n488), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n456), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n498));
  INV_X1    g297(.A(new_n405), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n447), .A2(new_n448), .B1(new_n272), .B2(new_n270), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n474), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n449), .A2(new_n406), .A3(new_n273), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT71), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n433), .B2(new_n434), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n444), .A2(new_n505), .A3(KEYINPUT36), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n438), .A2(new_n451), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT85), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT11), .B(G169gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G197gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT86), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT12), .ZN(new_n518));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(KEYINPUT13), .Z(new_n520));
  INV_X1    g319(.A(G43gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G50gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(G50gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n525));
  OR3_X1    g324(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n526), .A2(KEYINPUT87), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n527), .B2(KEYINPUT87), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n522), .B(new_n525), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(KEYINPUT15), .A3(new_n522), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT88), .B(G50gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n523), .B1(new_n533), .B2(new_n521), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n532), .B(new_n529), .C1(new_n534), .C2(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n526), .A2(new_n527), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n531), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT16), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(G1gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(G1gat), .B2(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G8gat), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n541), .B(new_n544), .C1(G1gat), .C2(new_n539), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n538), .A2(new_n546), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n520), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n538), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n531), .B(KEYINPUT17), .C1(new_n535), .C2(new_n537), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n553), .A2(new_n543), .A3(new_n545), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n546), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(KEYINPUT18), .A3(new_n519), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n538), .B(new_n546), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT89), .A3(new_n520), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n551), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n519), .A3(new_n556), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n518), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT91), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(KEYINPUT90), .A3(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n564), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n518), .B1(new_n569), .B2(KEYINPUT90), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT12), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n517), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n564), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n560), .B1(KEYINPUT90), .B2(new_n569), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT91), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n565), .B1(new_n571), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT98), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n584), .B2(new_n585), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n590), .A2(new_n591), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n582), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n590), .A2(new_n591), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT96), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G57gat), .B(G64gat), .Z(new_n599));
  INV_X1    g398(.A(KEYINPUT9), .ZN(new_n600));
  INV_X1    g399(.A(G71gat), .ZN(new_n601));
  INV_X1    g400(.A(G78gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G71gat), .B(G78gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n605), .A3(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(KEYINPUT92), .A3(new_n608), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n598), .A2(new_n613), .A3(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n592), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n607), .A2(KEYINPUT92), .A3(new_n608), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT92), .B1(new_n607), .B2(new_n608), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n609), .A2(new_n596), .A3(new_n592), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT10), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n581), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n609), .A2(new_n596), .A3(new_n592), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n613), .B2(new_n615), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n580), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n341), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(G204gat), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n625), .B(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n578), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n473), .A2(KEYINPUT38), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n325), .A2(new_n456), .A3(new_n326), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n453), .B1(new_n634), .B2(new_n462), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT82), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n497), .A2(new_n500), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n281), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT85), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n640), .B(new_n641), .C1(new_n451), .C2(new_n438), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n512), .A2(new_n631), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n546), .B1(new_n613), .B2(KEYINPUT21), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n336), .ZN(new_n645));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G127gat), .B(G155gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n236), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n647), .B(new_n649), .Z(new_n650));
  OR2_X1    g449(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n647), .B(new_n649), .ZN(new_n655));
  INV_X1    g454(.A(new_n653), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G134gat), .B(G162gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT95), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G232gat), .A2(G233gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT93), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n598), .A2(new_n538), .B1(KEYINPUT41), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n553), .A2(new_n597), .A3(new_n595), .A4(new_n554), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n666), .B2(new_n667), .ZN(new_n670));
  OAI22_X1  g469(.A1(new_n669), .A2(new_n670), .B1(KEYINPUT41), .B2(new_n665), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT97), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n665), .A2(KEYINPUT41), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G190gat), .B(G218gat), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT94), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n671), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n671), .B2(new_n676), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n662), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n671), .A2(new_n676), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n678), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n671), .A2(new_n676), .A3(new_n679), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n661), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n659), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n643), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n452), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G1gat), .ZN(G1324gat));
  INV_X1    g492(.A(new_n500), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT99), .B(G8gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT16), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n691), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  OR3_X1    g496(.A1(new_n697), .A2(KEYINPUT100), .A3(KEYINPUT42), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n699));
  OAI21_X1  g498(.A(G8gat), .B1(new_n690), .B2(new_n500), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT100), .B1(new_n697), .B2(KEYINPUT42), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n701), .ZN(G1325gat));
  AOI21_X1  g501(.A(G15gat), .B1(new_n691), .B2(new_n435), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n508), .A2(new_n509), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(G15gat), .B2(new_n706), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n690), .A2(new_n281), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n658), .A2(new_n630), .A3(new_n578), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n512), .A2(new_n642), .A3(new_n688), .A4(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G29gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n452), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n712), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n512), .A2(new_n688), .A3(new_n642), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT44), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n503), .A2(KEYINPUT101), .A3(new_n510), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n438), .A2(new_n451), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n640), .A2(KEYINPUT101), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n687), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n682), .A2(new_n686), .A3(KEYINPUT103), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n730));
  NAND3_X1  g529(.A1(new_n725), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n719), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n715), .B1(new_n732), .B2(new_n452), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n711), .B1(new_n718), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n716), .B(KEYINPUT45), .ZN(new_n735));
  INV_X1    g534(.A(new_n733), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(G1328gat));
  INV_X1    g537(.A(new_n732), .ZN(new_n739));
  OAI21_X1  g538(.A(G36gat), .B1(new_n739), .B2(new_n500), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n713), .A2(G36gat), .A3(new_n500), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1329gat));
  AOI21_X1  g542(.A(new_n521), .B1(new_n732), .B2(new_n704), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n713), .A2(G43gat), .A3(new_n444), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n745), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n746), .B(KEYINPUT47), .C1(new_n744), .C2(new_n749), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1330gat));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n281), .B(new_n719), .C1(new_n721), .C2(new_n731), .ZN(new_n755));
  INV_X1    g554(.A(new_n533), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n714), .A2(KEYINPUT106), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n713), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n758), .A2(new_n756), .A3(new_n502), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n755), .B2(new_n756), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n757), .A2(new_n762), .A3(KEYINPUT48), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  OAI221_X1 g563(.A(new_n761), .B1(new_n754), .B2(new_n764), .C1(new_n755), .C2(new_n756), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n763), .A2(new_n765), .ZN(G1331gat));
  AND4_X1   g565(.A1(new_n689), .A2(new_n725), .A3(new_n630), .A4(new_n578), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n452), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n694), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT49), .B(G64gat), .Z(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(G1333gat));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n601), .A3(new_n435), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n767), .A2(new_n704), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n601), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g576(.A1(new_n767), .A2(new_n502), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g578(.A1(new_n721), .A2(new_n731), .ZN(new_n780));
  INV_X1    g579(.A(new_n630), .ZN(new_n781));
  INV_X1    g580(.A(new_n565), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n568), .A2(new_n570), .A3(new_n566), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT91), .B1(new_n575), .B2(new_n576), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n658), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n787), .A2(new_n584), .A3(new_n327), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n658), .A2(new_n785), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n725), .A2(new_n688), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n688), .A4(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n452), .A3(new_n630), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n788), .B1(new_n584), .B2(new_n795), .ZN(G1336gat));
  OAI21_X1  g595(.A(G92gat), .B1(new_n787), .B2(new_n500), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n790), .A2(new_n799), .A3(KEYINPUT51), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT51), .B1(new_n790), .B2(new_n799), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n500), .A2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n800), .A2(new_n801), .A3(new_n781), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n794), .A2(new_n630), .A3(new_n802), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n797), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n787), .B2(new_n705), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n444), .A2(G99gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n630), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1338gat));
  XOR2_X1   g612(.A(KEYINPUT109), .B(G106gat), .Z(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n787), .B2(new_n281), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n281), .A2(G106gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n630), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n800), .A2(new_n801), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT53), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n794), .A2(new_n630), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT110), .ZN(new_n822));
  XNOR2_X1  g621(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n794), .A2(new_n824), .A3(new_n630), .A4(new_n817), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n822), .A2(new_n815), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n826), .ZN(G1339gat));
  AND4_X1   g626(.A1(new_n658), .A2(new_n687), .A3(new_n781), .A4(new_n578), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n598), .A2(new_n613), .A3(KEYINPUT10), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n580), .B(new_n829), .C1(new_n623), .C2(KEYINPUT10), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n621), .A2(new_n830), .A3(KEYINPUT54), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n621), .A2(new_n830), .A3(new_n833), .A4(KEYINPUT54), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n628), .B1(new_n621), .B2(KEYINPUT54), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n625), .A2(new_n629), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n837), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n516), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n558), .A2(new_n520), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT113), .Z(new_n847));
  AND2_X1   g646(.A1(new_n555), .A2(new_n556), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(new_n519), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n571), .A2(new_n577), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n844), .A2(new_n727), .A3(new_n728), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n845), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n630), .B(new_n853), .C1(new_n783), .C2(new_n784), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n854), .B(KEYINPUT114), .C1(new_n843), .C2(new_n578), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n727), .A2(new_n728), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT55), .B1(new_n835), .B2(new_n837), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n839), .B(new_n836), .C1(new_n832), .C2(new_n834), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n785), .A2(new_n841), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT114), .B1(new_n861), .B2(new_n854), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n852), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n828), .B1(new_n863), .B2(new_n659), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT115), .B1(new_n864), .B2(new_n502), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n854), .B1(new_n843), .B2(new_n578), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n856), .A3(new_n855), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n658), .B1(new_n870), .B2(new_n852), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n866), .B(new_n281), .C1(new_n871), .C2(new_n828), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n865), .A2(new_n435), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n694), .A2(new_n327), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n578), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n864), .A2(new_n502), .A3(new_n444), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n874), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n285), .A3(new_n785), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n879), .ZN(G1340gat));
  OAI21_X1  g679(.A(G120gat), .B1(new_n875), .B2(new_n781), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n283), .A3(new_n630), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1341gat));
  NOR3_X1   g682(.A1(new_n875), .A2(new_n288), .A3(new_n659), .ZN(new_n884));
  AOI21_X1  g683(.A(G127gat), .B1(new_n878), .B2(new_n658), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(G1342gat));
  NAND3_X1  g685(.A1(new_n878), .A2(new_n293), .A3(new_n688), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT56), .Z(new_n888));
  OAI21_X1  g687(.A(G134gat), .B1(new_n875), .B2(new_n687), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1343gat));
  NAND2_X1  g689(.A1(new_n863), .A2(new_n659), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n658), .A2(new_n687), .A3(new_n781), .A4(new_n578), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n281), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n705), .A2(new_n874), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(G141gat), .A3(new_n578), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n867), .A2(new_n687), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n658), .B1(new_n898), .B2(new_n852), .ZN(new_n899));
  OAI211_X1 g698(.A(KEYINPUT57), .B(new_n502), .C1(new_n899), .C2(new_n828), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n851), .A2(new_n860), .A3(new_n841), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n729), .A2(new_n903), .B1(new_n687), .B2(new_n867), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n892), .B1(new_n904), .B2(new_n658), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n905), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n502), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n902), .B(new_n906), .C1(new_n893), .C2(KEYINPUT57), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n907), .A2(KEYINPUT117), .A3(new_n895), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT117), .B1(new_n907), .B2(new_n895), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n785), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n897), .B1(new_n910), .B2(G141gat), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n907), .A2(new_n895), .ZN(new_n913));
  OAI21_X1  g712(.A(G141gat), .B1(new_n913), .B2(new_n578), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n912), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n897), .B(KEYINPUT118), .ZN(new_n916));
  OAI22_X1  g715(.A1(new_n911), .A2(new_n912), .B1(new_n915), .B2(new_n916), .ZN(G1344gat));
  NAND2_X1  g716(.A1(new_n903), .A2(new_n688), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n658), .B1(new_n898), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n502), .B1(new_n919), .B2(new_n828), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT119), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI211_X1 g721(.A(KEYINPUT57), .B(new_n502), .C1(new_n871), .C2(new_n828), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n893), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n926), .A2(KEYINPUT59), .A3(new_n630), .A4(new_n895), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n907), .A2(KEYINPUT117), .A3(new_n895), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n781), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n931), .B2(KEYINPUT59), .ZN(new_n932));
  INV_X1    g731(.A(new_n896), .ZN(new_n933));
  AOI21_X1  g732(.A(G148gat), .B1(new_n933), .B2(new_n630), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n932), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n934), .ZN(G1345gat));
  NOR2_X1   g734(.A1(new_n896), .A2(new_n659), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT120), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n658), .B1(new_n908), .B2(new_n909), .ZN(new_n938));
  MUX2_X1   g737(.A(new_n937), .B(new_n938), .S(G155gat), .Z(G1346gat));
  OAI21_X1  g738(.A(new_n729), .B1(new_n908), .B2(new_n909), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n942), .B(new_n729), .C1(new_n908), .C2(new_n909), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(G162gat), .A3(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n896), .A2(G162gat), .A3(new_n687), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT121), .Z(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1347gat));
  NOR2_X1   g746(.A1(new_n500), .A2(new_n452), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n877), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n340), .A3(new_n785), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n865), .A2(new_n872), .A3(new_n435), .A4(new_n948), .ZN(new_n951));
  OAI21_X1  g750(.A(G169gat), .B1(new_n951), .B2(new_n578), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT123), .Z(G1348gat));
  AOI21_X1  g753(.A(G176gat), .B1(new_n949), .B2(new_n630), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n951), .A2(new_n341), .A3(new_n781), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(G1349gat));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n873), .A2(new_n958), .A3(new_n658), .A4(new_n948), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT124), .B1(new_n951), .B2(new_n659), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(G183gat), .A3(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT60), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n949), .A2(new_n658), .A3(new_n379), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n963), .B1(new_n961), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(G1350gat));
  OAI21_X1  g766(.A(G190gat), .B1(new_n951), .B2(new_n687), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT61), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n337), .A3(new_n729), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1351gat));
  NAND2_X1  g770(.A1(new_n705), .A2(new_n948), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n926), .A2(new_n785), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G197gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n893), .A2(new_n973), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n976), .A2(G197gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n975), .B1(new_n578), .B2(new_n977), .ZN(G1352gat));
  NOR3_X1   g777(.A1(new_n976), .A2(G204gat), .A3(new_n781), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT62), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n926), .A2(new_n630), .A3(new_n973), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G204gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1353gat));
  INV_X1    g782(.A(new_n976), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n984), .A2(new_n236), .A3(new_n658), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n924), .A2(new_n925), .A3(new_n658), .A4(new_n973), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n991), .B(new_n985), .C1(new_n987), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1354gat));
  NAND3_X1  g792(.A1(new_n926), .A2(new_n688), .A3(new_n973), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(G218gat), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n984), .A2(new_n237), .A3(new_n729), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(KEYINPUT127), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n995), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1000), .ZN(G1355gat));
endmodule


