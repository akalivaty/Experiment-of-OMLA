

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n530), .A2(G2104), .ZN(n888) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(n527), .Z(n879) );
  NOR2_X1 U555 ( .A1(n535), .A2(n534), .ZN(G160) );
  AND2_X1 U556 ( .A1(n521), .A2(n812), .ZN(n520) );
  AND2_X1 U557 ( .A1(n795), .A2(n794), .ZN(n521) );
  OR2_X1 U558 ( .A1(n770), .A2(n769), .ZN(n522) );
  AND2_X1 U559 ( .A1(n767), .A2(n766), .ZN(n523) );
  NOR2_X1 U560 ( .A1(n731), .A2(n945), .ZN(n692) );
  NOR2_X1 U561 ( .A1(n967), .A2(n695), .ZN(n701) );
  AND2_X1 U562 ( .A1(n738), .A2(n736), .ZN(n725) );
  NOR2_X1 U563 ( .A1(n726), .A2(n725), .ZN(n727) );
  INV_X1 U564 ( .A(KEYINPUT99), .ZN(n762) );
  XNOR2_X1 U565 ( .A(n763), .B(n762), .ZN(n765) );
  NAND2_X1 U566 ( .A1(G160), .A2(G40), .ZN(n773) );
  NOR2_X1 U567 ( .A1(G651), .A2(n631), .ZN(n649) );
  NOR2_X1 U568 ( .A1(G543), .A2(G651), .ZN(n655) );
  XNOR2_X1 U569 ( .A(n542), .B(KEYINPUT87), .ZN(n772) );
  INV_X1 U570 ( .A(n772), .ZN(G164) );
  INV_X1 U571 ( .A(G2105), .ZN(n530) );
  NAND2_X1 U572 ( .A1(G101), .A2(n888), .ZN(n526) );
  XNOR2_X1 U573 ( .A(KEYINPUT23), .B(KEYINPUT66), .ZN(n524) );
  XNOR2_X1 U574 ( .A(n524), .B(KEYINPUT65), .ZN(n525) );
  XNOR2_X1 U575 ( .A(n526), .B(n525), .ZN(n529) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n879), .A2(G137), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n535) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U580 ( .A1(n881), .A2(G113), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n530), .A2(G2104), .ZN(n531) );
  XNOR2_X1 U582 ( .A(n531), .B(KEYINPUT64), .ZN(n883) );
  NAND2_X1 U583 ( .A1(G125), .A2(n883), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n534) );
  AND2_X1 U585 ( .A1(n879), .A2(G138), .ZN(n541) );
  NAND2_X1 U586 ( .A1(G126), .A2(n883), .ZN(n539) );
  NAND2_X1 U587 ( .A1(G114), .A2(n881), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G102), .A2(n888), .ZN(n536) );
  AND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n542) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G651), .ZN(n546) );
  NOR2_X1 U594 ( .A1(G543), .A2(n546), .ZN(n543) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n543), .Z(n648) );
  NAND2_X1 U596 ( .A1(G65), .A2(n648), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G91), .A2(n655), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n550) );
  XOR2_X1 U599 ( .A(G543), .B(KEYINPUT0), .Z(n631) );
  NAND2_X1 U600 ( .A1(G53), .A2(n649), .ZN(n548) );
  NOR2_X1 U601 ( .A1(n631), .A2(n546), .ZN(n646) );
  NAND2_X1 U602 ( .A1(G78), .A2(n646), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n705) );
  INV_X1 U605 ( .A(n705), .ZN(G299) );
  INV_X1 U606 ( .A(G132), .ZN(G219) );
  INV_X1 U607 ( .A(G82), .ZN(G220) );
  NAND2_X1 U608 ( .A1(G64), .A2(n648), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G52), .A2(n649), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G77), .A2(n646), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G90), .A2(n655), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U615 ( .A1(n557), .A2(n556), .ZN(G171) );
  NAND2_X1 U616 ( .A1(G63), .A2(n648), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G51), .A2(n649), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(KEYINPUT6), .B(n560), .ZN(n568) );
  NAND2_X1 U620 ( .A1(n646), .A2(G76), .ZN(n561) );
  XNOR2_X1 U621 ( .A(KEYINPUT74), .B(n561), .ZN(n565) );
  XOR2_X1 U622 ( .A(KEYINPUT73), .B(KEYINPUT4), .Z(n563) );
  NAND2_X1 U623 ( .A1(G89), .A2(n655), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U626 ( .A(n566), .B(KEYINPUT5), .Z(n567) );
  NOR2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U628 ( .A(KEYINPUT75), .B(n569), .Z(n570) );
  XOR2_X1 U629 ( .A(KEYINPUT7), .B(n570), .Z(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U632 ( .A(n571), .B(KEYINPUT70), .ZN(n572) );
  XNOR2_X1 U633 ( .A(KEYINPUT10), .B(n572), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n822) );
  NAND2_X1 U635 ( .A1(n822), .A2(G567), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n648), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n574), .Z(n581) );
  NAND2_X1 U639 ( .A1(G81), .A2(n655), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT71), .B(n575), .Z(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G68), .A2(n646), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n579), .Z(n580) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n649), .A2(G43), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n967) );
  INV_X1 U648 ( .A(G860), .ZN(n613) );
  OR2_X1 U649 ( .A1(n967), .A2(n613), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U652 ( .A1(G92), .A2(n655), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G66), .A2(n648), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G79), .A2(n646), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n649), .A2(G54), .ZN(n586) );
  XOR2_X1 U657 ( .A(KEYINPUT72), .B(n586), .Z(n587) );
  NOR2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT15), .ZN(n976) );
  OR2_X1 U661 ( .A1(n976), .A2(G868), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(G284) );
  INV_X1 U663 ( .A(G868), .ZN(n594) );
  NOR2_X1 U664 ( .A1(G286), .A2(n594), .ZN(n596) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U666 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n613), .A2(G559), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n597), .A2(n976), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U670 ( .A1(G868), .A2(n967), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G868), .A2(n976), .ZN(n599) );
  NOR2_X1 U672 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U673 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U674 ( .A1(G123), .A2(n883), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G135), .A2(n879), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U678 ( .A(KEYINPUT76), .B(n605), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G111), .A2(n881), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G99), .A2(n888), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n925) );
  XNOR2_X1 U683 ( .A(G2096), .B(n925), .ZN(n611) );
  INV_X1 U684 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U686 ( .A1(G559), .A2(n976), .ZN(n612) );
  XOR2_X1 U687 ( .A(n967), .B(n612), .Z(n666) );
  NAND2_X1 U688 ( .A1(n613), .A2(n666), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G67), .A2(n648), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G55), .A2(n649), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U692 ( .A(KEYINPUT78), .B(n616), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G80), .A2(n646), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G93), .A2(n655), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U696 ( .A(KEYINPUT77), .B(n619), .Z(n620) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n668) );
  XOR2_X1 U698 ( .A(n622), .B(n668), .Z(G145) );
  NAND2_X1 U699 ( .A1(G86), .A2(n655), .ZN(n629) );
  NAND2_X1 U700 ( .A1(G61), .A2(n648), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G48), .A2(n649), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n646), .A2(G73), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n630), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G87), .A2(n631), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n648), .A2(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G49), .A2(n649), .ZN(n635) );
  XOR2_X1 U713 ( .A(KEYINPUT79), .B(n635), .Z(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G60), .A2(n648), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G47), .A2(n649), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U718 ( .A(KEYINPUT68), .B(n640), .ZN(n643) );
  NAND2_X1 U719 ( .A1(G72), .A2(n646), .ZN(n641) );
  XNOR2_X1 U720 ( .A(KEYINPUT67), .B(n641), .ZN(n642) );
  NOR2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n655), .A2(G85), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U724 ( .A1(G75), .A2(n646), .ZN(n647) );
  XOR2_X1 U725 ( .A(KEYINPUT82), .B(n647), .Z(n654) );
  NAND2_X1 U726 ( .A1(G62), .A2(n648), .ZN(n651) );
  NAND2_X1 U727 ( .A1(G50), .A2(n649), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U729 ( .A(KEYINPUT81), .B(n652), .Z(n653) );
  NOR2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n655), .A2(G88), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(G303) );
  INV_X1 U733 ( .A(G303), .ZN(G166) );
  XOR2_X1 U734 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n658) );
  XNOR2_X1 U735 ( .A(G288), .B(n658), .ZN(n659) );
  XOR2_X1 U736 ( .A(n659), .B(KEYINPUT84), .Z(n661) );
  XNOR2_X1 U737 ( .A(n705), .B(KEYINPUT83), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n668), .B(n662), .ZN(n664) );
  XNOR2_X1 U740 ( .A(G290), .B(G166), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U742 ( .A(G305), .B(n665), .Z(n908) );
  XNOR2_X1 U743 ( .A(n666), .B(n908), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n667), .A2(G868), .ZN(n670) );
  OR2_X1 U745 ( .A1(G868), .A2(n668), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U751 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U754 ( .A1(G108), .A2(G120), .ZN(n675) );
  NOR2_X1 U755 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G69), .A2(n676), .ZN(n827) );
  NAND2_X1 U757 ( .A1(G567), .A2(n827), .ZN(n681) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U760 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(G96), .A2(n679), .ZN(n828) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n828), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U764 ( .A(KEYINPUT86), .B(n682), .Z(G319) );
  INV_X1 U765 ( .A(G319), .ZN(n684) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U767 ( .A1(n684), .A2(n683), .ZN(n826) );
  NAND2_X1 U768 ( .A1(n826), .A2(G36), .ZN(G176) );
  INV_X1 U769 ( .A(n773), .ZN(n685) );
  INV_X1 U770 ( .A(G1384), .ZN(n771) );
  AND2_X1 U771 ( .A1(n685), .A2(n771), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n686), .A2(n772), .ZN(n731) );
  NAND2_X1 U773 ( .A1(G8), .A2(n731), .ZN(n770) );
  NOR2_X1 U774 ( .A1(G1966), .A2(n770), .ZN(n726) );
  INV_X1 U775 ( .A(n731), .ZN(n712) );
  NAND2_X1 U776 ( .A1(n712), .A2(G2072), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT27), .ZN(n689) );
  INV_X1 U778 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U779 ( .A1(n998), .A2(n712), .ZN(n688) );
  NOR2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n704) );
  NOR2_X1 U781 ( .A1(n705), .A2(n704), .ZN(n690) );
  XOR2_X1 U782 ( .A(n690), .B(KEYINPUT28), .Z(n709) );
  INV_X1 U783 ( .A(G1996), .ZN(n945) );
  INV_X1 U784 ( .A(KEYINPUT26), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n692), .B(n691), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n731), .A2(G1341), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n701), .A2(n976), .ZN(n699) );
  NOR2_X1 U789 ( .A1(n712), .A2(G1348), .ZN(n697) );
  NOR2_X1 U790 ( .A1(G2067), .A2(n731), .ZN(n696) );
  NOR2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U793 ( .A(n700), .B(KEYINPUT93), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n976), .A2(n701), .ZN(n702) );
  OR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n711) );
  XOR2_X1 U799 ( .A(KEYINPUT94), .B(KEYINPUT29), .Z(n710) );
  XNOR2_X1 U800 ( .A(n711), .B(n710), .ZN(n716) );
  NAND2_X1 U801 ( .A1(G1961), .A2(n731), .ZN(n714) );
  XOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .Z(n947) );
  NAND2_X1 U803 ( .A1(n712), .A2(n947), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n717) );
  OR2_X1 U805 ( .A1(G301), .A2(n717), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n738) );
  NAND2_X1 U807 ( .A1(G301), .A2(n717), .ZN(n718) );
  XNOR2_X1 U808 ( .A(n718), .B(KEYINPUT95), .ZN(n723) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n731), .ZN(n728) );
  NOR2_X1 U810 ( .A1(n728), .A2(n726), .ZN(n719) );
  NAND2_X1 U811 ( .A1(G8), .A2(n719), .ZN(n720) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n720), .ZN(n721) );
  NOR2_X1 U813 ( .A1(n721), .A2(G168), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U815 ( .A(KEYINPUT31), .B(n724), .Z(n736) );
  XNOR2_X1 U816 ( .A(n727), .B(KEYINPUT96), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n728), .A2(G8), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n746) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n731), .ZN(n732) );
  XNOR2_X1 U820 ( .A(KEYINPUT97), .B(n732), .ZN(n735) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n770), .ZN(n733) );
  NOR2_X1 U822 ( .A1(G166), .A2(n733), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n739) );
  AND2_X1 U824 ( .A1(n736), .A2(n739), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n742) );
  INV_X1 U826 ( .A(n739), .ZN(n740) );
  OR2_X1 U827 ( .A1(n740), .A2(G286), .ZN(n741) );
  AND2_X1 U828 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U829 ( .A1(n743), .A2(G8), .ZN(n744) );
  XNOR2_X1 U830 ( .A(n744), .B(KEYINPUT32), .ZN(n745) );
  NAND2_X1 U831 ( .A1(n746), .A2(n745), .ZN(n753) );
  NOR2_X1 U832 ( .A1(G2090), .A2(G303), .ZN(n747) );
  NAND2_X1 U833 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n753), .A2(n748), .ZN(n749) );
  NAND2_X1 U835 ( .A1(n749), .A2(n770), .ZN(n767) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n970) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n970), .A2(n750), .ZN(n751) );
  XNOR2_X1 U839 ( .A(n751), .B(KEYINPUT98), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n757) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U842 ( .A(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n974), .A2(n754), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n755), .A2(n770), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n761) );
  INV_X1 U846 ( .A(n770), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n970), .A2(n758), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n759), .A2(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n763) );
  XOR2_X1 U850 ( .A(G305), .B(G1981), .Z(n764) );
  XNOR2_X1 U851 ( .A(KEYINPUT100), .B(n764), .ZN(n983) );
  NAND2_X1 U852 ( .A1(n765), .A2(n983), .ZN(n766) );
  NOR2_X1 U853 ( .A1(G305), .A2(G1981), .ZN(n768) );
  XOR2_X1 U854 ( .A(n768), .B(KEYINPUT24), .Z(n769) );
  NAND2_X1 U855 ( .A1(n523), .A2(n522), .ZN(n806) );
  XNOR2_X1 U856 ( .A(G1986), .B(G290), .ZN(n969) );
  AND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n774) );
  NOR2_X1 U858 ( .A1(n774), .A2(n773), .ZN(n817) );
  NAND2_X1 U859 ( .A1(n969), .A2(n817), .ZN(n775) );
  XNOR2_X1 U860 ( .A(n775), .B(KEYINPUT88), .ZN(n795) );
  NAND2_X1 U861 ( .A1(G107), .A2(n881), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G95), .A2(n888), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U864 ( .A1(n883), .A2(G119), .ZN(n778) );
  XOR2_X1 U865 ( .A(KEYINPUT90), .B(n778), .Z(n779) );
  NOR2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n879), .A2(G131), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n877) );
  NAND2_X1 U869 ( .A1(G1991), .A2(n877), .ZN(n783) );
  XOR2_X1 U870 ( .A(KEYINPUT91), .B(n783), .Z(n793) );
  NAND2_X1 U871 ( .A1(G105), .A2(n888), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT38), .ZN(n791) );
  NAND2_X1 U873 ( .A1(n879), .A2(G141), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G129), .A2(n883), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n881), .A2(G117), .ZN(n787) );
  XOR2_X1 U877 ( .A(KEYINPUT92), .B(n787), .Z(n788) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n896) );
  NAND2_X1 U880 ( .A1(G1996), .A2(n896), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n924) );
  NAND2_X1 U882 ( .A1(n924), .A2(n817), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n881), .A2(G116), .ZN(n797) );
  NAND2_X1 U884 ( .A1(G128), .A2(n883), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(KEYINPUT35), .ZN(n803) );
  NAND2_X1 U887 ( .A1(G140), .A2(n879), .ZN(n800) );
  NAND2_X1 U888 ( .A1(G104), .A2(n888), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U890 ( .A(KEYINPUT34), .B(n801), .Z(n802) );
  NAND2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(KEYINPUT36), .ZN(n900) );
  XOR2_X1 U893 ( .A(G2067), .B(KEYINPUT37), .Z(n814) );
  NAND2_X1 U894 ( .A1(n900), .A2(n814), .ZN(n805) );
  XNOR2_X1 U895 ( .A(n805), .B(KEYINPUT89), .ZN(n929) );
  NAND2_X1 U896 ( .A1(n817), .A2(n929), .ZN(n812) );
  NAND2_X1 U897 ( .A1(n806), .A2(n520), .ZN(n820) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n896), .ZN(n920) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U900 ( .A1(G1991), .A2(n877), .ZN(n923) );
  NOR2_X1 U901 ( .A1(n807), .A2(n923), .ZN(n808) );
  NOR2_X1 U902 ( .A1(n924), .A2(n808), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n920), .A2(n809), .ZN(n811) );
  XOR2_X1 U904 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n810) );
  XNOR2_X1 U905 ( .A(n811), .B(n810), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n816) );
  NOR2_X1 U907 ( .A1(n814), .A2(n900), .ZN(n815) );
  XOR2_X1 U908 ( .A(KEYINPUT102), .B(n815), .Z(n936) );
  NAND2_X1 U909 ( .A1(n816), .A2(n936), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U912 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n822), .ZN(G217) );
  NAND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n823) );
  XNOR2_X1 U915 ( .A(KEYINPUT107), .B(n823), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(G661), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G108), .ZN(G238) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XOR2_X1 U926 ( .A(G2443), .B(G2451), .Z(n830) );
  XNOR2_X1 U927 ( .A(KEYINPUT104), .B(G2427), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U929 ( .A(n831), .B(G2430), .Z(n833) );
  XNOR2_X1 U930 ( .A(G1341), .B(G1348), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U932 ( .A(G2438), .B(G2435), .Z(n835) );
  XNOR2_X1 U933 ( .A(KEYINPUT105), .B(G2454), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U935 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2446), .B(KEYINPUT103), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  NAND2_X1 U938 ( .A1(G14), .A2(n840), .ZN(n841) );
  XOR2_X1 U939 ( .A(KEYINPUT106), .B(n841), .Z(G401) );
  XOR2_X1 U940 ( .A(G2096), .B(KEYINPUT108), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2090), .B(KEYINPUT43), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n844), .B(KEYINPUT42), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U946 ( .A(G2678), .B(G2100), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2084), .B(G2078), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n852) );
  XNOR2_X1 U951 ( .A(G1961), .B(G1956), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U956 ( .A(G2474), .B(G1981), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1966), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G112), .A2(n881), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G100), .A2(n888), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U963 ( .A1(n883), .A2(G124), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n862), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G136), .A2(n879), .ZN(n863) );
  XOR2_X1 U966 ( .A(KEYINPUT109), .B(n863), .Z(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U968 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G118), .A2(n881), .ZN(n876) );
  XNOR2_X1 U970 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G142), .A2(n879), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G106), .A2(n888), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n871), .B(n870), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G130), .A2(n883), .ZN(n872) );
  XOR2_X1 U976 ( .A(KEYINPUT110), .B(n872), .Z(n873) );
  NOR2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n905) );
  XOR2_X1 U980 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n894) );
  NAND2_X1 U981 ( .A1(n879), .A2(G139), .ZN(n880) );
  XNOR2_X1 U982 ( .A(KEYINPUT113), .B(n880), .ZN(n892) );
  NAND2_X1 U983 ( .A1(n881), .A2(G115), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n882), .B(KEYINPUT114), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G127), .A2(n883), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U987 ( .A(KEYINPUT115), .B(n886), .Z(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(KEYINPUT47), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G103), .A2(n888), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  NOR2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n932) );
  XNOR2_X1 U992 ( .A(n932), .B(KEYINPUT116), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U994 ( .A(KEYINPUT117), .B(n895), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n896), .B(KEYINPUT46), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(n899), .B(G162), .Z(n902) );
  XNOR2_X1 U998 ( .A(G164), .B(n900), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(G160), .B(n903), .Z(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n906), .B(n925), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(n967), .B(n908), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(G171), .B(n976), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n911), .B(G286), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n913) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n914), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G401), .A2(n915), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n916), .B(KEYINPUT118), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n921), .Z(n931) );
  XOR2_X1 U1020 ( .A(G2084), .B(G160), .Z(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n939) );
  XOR2_X1 U1026 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1031 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n940), .ZN(n941) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n963), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n942), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n958) );
  XNOR2_X1 U1037 ( .A(G1991), .B(G25), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(G32), .B(n945), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G27), .B(n947), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT120), .B(n948), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1046 ( .A(KEYINPUT119), .B(G2067), .Z(n953) );
  XNOR2_X1 U1047 ( .A(G26), .B(n953), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1055 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n966), .ZN(n1023) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1059 ( .A(G1341), .B(n967), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n990) );
  XNOR2_X1 U1061 ( .A(G303), .B(G1971), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(n970), .B(KEYINPUT122), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(n975), .B(KEYINPUT123), .ZN(n982) );
  XNOR2_X1 U1066 ( .A(n976), .B(G1348), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G171), .B(G1961), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G299), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n988) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(n985), .B(KEYINPUT121), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(n986), .B(KEYINPUT57), .ZN(n987) );
  NOR2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n1021) );
  INV_X1 U1079 ( .A(G16), .ZN(n1019) );
  XOR2_X1 U1080 ( .A(G1961), .B(G5), .Z(n1004) );
  XNOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n993), .B(G4), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(KEYINPUT124), .B(n998), .Z(n999) );
  XNOR2_X1 U1088 ( .A(G20), .B(n999), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(n1002), .B(KEYINPUT60), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G21), .B(G1966), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1015) );
  XOR2_X1 U1094 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n1013) );
  XNOR2_X1 U1095 ( .A(G1986), .B(G24), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G1976), .B(KEYINPUT125), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(G23), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(n1016), .B(KEYINPUT61), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT127), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

