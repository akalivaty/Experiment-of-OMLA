//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  OR2_X1    g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT26), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  OAI22_X1  g004(.A1(new_n202), .A2(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT26), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT28), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(new_n205), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT27), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n213), .A2(new_n219), .A3(KEYINPUT67), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n204), .A2(KEYINPUT27), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(G183gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(new_n205), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT28), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n210), .B1(new_n220), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n207), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n202), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n208), .B2(KEYINPUT23), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n202), .A2(KEYINPUT64), .A3(new_n230), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n205), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237));
  OAI21_X1  g036(.A(G190gat), .B1(new_n237), .B2(new_n204), .ZN(new_n238));
  NOR2_X1   g037(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n207), .B1(KEYINPUT23), .B2(new_n208), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT64), .B1(new_n202), .B2(new_n230), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n208), .A2(new_n232), .A3(KEYINPUT23), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n242), .B(new_n243), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n235), .A2(new_n241), .B1(new_n246), .B2(KEYINPUT25), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NOR4_X1   g048(.A1(new_n248), .A2(new_n242), .A3(new_n240), .A4(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n228), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(G127gat), .A2(G134gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(G127gat), .A2(G134gat), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G113gat), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT70), .ZN(new_n259));
  OR3_X1    g058(.A1(new_n257), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n254), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(G127gat), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G127gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G127gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n268), .A3(G134gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n256), .A2(new_n258), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n264), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n261), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n264), .A2(new_n269), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n254), .A2(new_n259), .A3(new_n260), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n251), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n246), .A2(KEYINPUT25), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n234), .A2(new_n233), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n241), .A2(new_n283), .A3(new_n243), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n235), .A2(KEYINPUT65), .A3(KEYINPUT25), .A4(new_n241), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n287), .A2(new_n273), .A3(new_n279), .A4(new_n228), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G227gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G71gat), .B(G99gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT33), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n288), .A3(new_n290), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(KEYINPUT34), .Z(new_n302));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n292), .A2(new_n303), .A3(new_n297), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n290), .B1(new_n281), .B2(new_n288), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT72), .B1(new_n305), .B2(KEYINPUT33), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n296), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n300), .B(new_n302), .C1(new_n307), .C2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n302), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n304), .B2(new_n306), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(new_n299), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G78gat), .B(G106gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT83), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G22gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT31), .B(G50gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  INV_X1    g121(.A(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G218gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT73), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  AND2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT77), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G155gat), .ZN(new_n337));
  INV_X1    g136(.A(G162gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(KEYINPUT78), .A3(KEYINPUT2), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G141gat), .B(G148gat), .Z(new_n345));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n334), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n341), .A2(new_n350), .A3(KEYINPUT2), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G141gat), .B(G148gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n350), .B1(new_n341), .B2(KEYINPUT2), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n341), .ZN(new_n356));
  OAI221_X1 g155(.A(new_n333), .B1(new_n344), .B2(new_n349), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n330), .A2(new_n332), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n344), .A2(new_n349), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n353), .A2(new_n354), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n356), .B1(new_n361), .B2(new_n351), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n328), .A2(new_n358), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n333), .ZN(new_n365));
  OAI211_X1 g164(.A(G228gat), .B(G233gat), .C1(new_n359), .C2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n328), .B1(new_n357), .B2(new_n358), .ZN(new_n367));
  AND2_X1   g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368));
  OR3_X1    g167(.A1(new_n367), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n320), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n369), .A3(new_n320), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n318), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  INV_X1    g173(.A(new_n318), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n374), .A2(new_n375), .A3(new_n370), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n315), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n251), .B2(new_n358), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n287), .B2(new_n228), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n382), .A2(new_n328), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n330), .A2(new_n332), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT67), .B1(new_n213), .B2(new_n219), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n225), .A2(new_n221), .A3(new_n226), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n285), .A2(new_n286), .B1(new_n388), .B2(new_n210), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n380), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n251), .A2(new_n381), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n379), .B1(new_n384), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n385), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(new_n382), .B2(new_n383), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n329), .A3(new_n391), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT74), .ZN(new_n397));
  XOR2_X1   g196(.A(G8gat), .B(G36gat), .Z(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n400), .B(KEYINPUT75), .Z(new_n401));
  NAND3_X1  g200(.A1(new_n393), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n384), .B2(new_n392), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT30), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n395), .A2(new_n396), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT30), .A3(new_n400), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT0), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n411), .B(new_n412), .Z(new_n413));
  OAI21_X1  g212(.A(KEYINPUT3), .B1(new_n360), .B2(new_n362), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n276), .A2(new_n278), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n357), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n417));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n363), .A2(new_n273), .A3(new_n420), .A4(new_n279), .ZN(new_n421));
  OAI22_X1  g220(.A1(new_n355), .A2(new_n356), .B1(new_n344), .B2(new_n349), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT4), .B1(new_n422), .B2(new_n415), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT80), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT80), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n419), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n421), .A2(new_n426), .A3(new_n423), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n426), .B1(new_n421), .B2(new_n423), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT81), .A3(new_n419), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n422), .B(new_n415), .ZN(new_n436));
  INV_X1    g235(.A(new_n418), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n417), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n363), .A2(new_n273), .A3(new_n279), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT4), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n363), .A2(new_n420), .A3(new_n276), .A4(new_n278), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n440), .A2(KEYINPUT79), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n418), .B(new_n416), .C1(new_n440), .C2(KEYINPUT79), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n413), .B1(new_n435), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT6), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT81), .B1(new_n433), .B2(new_n419), .ZN(new_n448));
  AND4_X1   g247(.A1(KEYINPUT81), .A2(new_n419), .A3(new_n425), .A4(new_n427), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n413), .B(new_n444), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n450), .A2(KEYINPUT82), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT82), .B1(new_n450), .B2(new_n451), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n452), .A2(new_n453), .A3(new_n445), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n378), .B(new_n409), .C1(new_n447), .C2(new_n454), .ZN(new_n455));
  NOR4_X1   g254(.A1(new_n315), .A2(new_n377), .A3(KEYINPUT35), .A4(new_n408), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT85), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n450), .A2(new_n451), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(new_n445), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n460));
  INV_X1    g259(.A(new_n413), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n462), .A2(KEYINPUT85), .A3(new_n451), .A4(new_n450), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n446), .A3(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n455), .A2(KEYINPUT35), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n393), .A2(KEYINPUT37), .A3(new_n397), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT37), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n400), .B1(new_n406), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n384), .B2(new_n392), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n401), .A2(new_n467), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n329), .B1(new_n390), .B2(new_n391), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n390), .A2(new_n391), .A3(new_n385), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT37), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n403), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n377), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n425), .A2(new_n416), .A3(new_n427), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n437), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n436), .A2(new_n437), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT39), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n487), .A3(new_n437), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n486), .A2(KEYINPUT40), .A3(new_n413), .A4(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT84), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT40), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n413), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n485), .A2(KEYINPUT39), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n437), .B2(new_n483), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n491), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n408), .A2(new_n462), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n482), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n466), .B1(new_n481), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n408), .A2(new_n462), .A3(new_n495), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n492), .A2(new_n494), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT84), .A3(KEYINPUT40), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n489), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n377), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n479), .A2(new_n446), .A3(new_n459), .A4(new_n463), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT86), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n311), .A2(new_n314), .A3(KEYINPUT36), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT36), .B1(new_n311), .B2(new_n314), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n409), .B1(new_n454), .B2(new_n447), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n377), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n465), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(G1gat), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  OAI221_X1 g317(.A(new_n517), .B1(KEYINPUT89), .B2(new_n518), .C1(G1gat), .C2(new_n515), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT87), .ZN(new_n523));
  NOR3_X1   g322(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n526), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n524), .B(KEYINPUT88), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n532), .A2(new_n523), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n534), .A2(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(KEYINPUT17), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n521), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n537), .A2(new_n538), .B1(new_n521), .B2(new_n534), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT90), .B1(new_n540), .B2(new_n521), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT91), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT18), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n539), .A2(new_n541), .A3(KEYINPUT18), .A4(new_n543), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n521), .B(new_n534), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n543), .B(KEYINPUT13), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G197gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT11), .B(G169gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT12), .Z(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n546), .A2(new_n558), .A3(new_n547), .A4(new_n550), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n514), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G57gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(G64gat), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT92), .B(G57gat), .Z(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(G64gat), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n565), .B1(KEYINPUT9), .B2(new_n566), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n521), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n579), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n576), .A2(new_n577), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT93), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT94), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G183gat), .B(G211gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n589), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n588), .B(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n591), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n584), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n591), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n592), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n599), .A3(new_n583), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT95), .B(G92gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  INV_X1    g405(.A(G99gat), .ZN(new_n607));
  INV_X1    g406(.A(G106gat), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT8), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT96), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n617), .A2(new_n534), .B1(KEYINPUT41), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n616), .B(KEYINPUT97), .Z(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n620), .B2(new_n540), .ZN(new_n621));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n601), .A2(new_n629), .A3(KEYINPUT98), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT98), .B1(new_n601), .B2(new_n629), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT99), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n613), .B1(new_n610), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n611), .A2(KEYINPUT99), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n615), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n636), .A3(new_n634), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n576), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n576), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n616), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n639), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n633), .A2(new_n634), .B1(new_n615), .B2(new_n636), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n643), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT10), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n616), .A2(new_n650), .A3(new_n576), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n641), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n641), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n650), .B1(new_n640), .B2(new_n643), .ZN(new_n656));
  INV_X1    g455(.A(new_n651), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT101), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n644), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  OR3_X1    g463(.A1(new_n660), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n660), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n664), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n658), .A2(new_n668), .A3(new_n644), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n630), .A2(new_n631), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n562), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n562), .A2(KEYINPUT103), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n454), .A2(new_n447), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  AND3_X1   g480(.A1(new_n677), .A2(new_n408), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n518), .B1(new_n677), .B2(new_n408), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n682), .ZN(G1325gat));
  INV_X1    g484(.A(new_n677), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n686), .A2(G15gat), .A3(new_n315), .ZN(new_n687));
  INV_X1    g486(.A(new_n511), .ZN(new_n688));
  OAI21_X1  g487(.A(G15gat), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(G1326gat));
  NOR3_X1   g489(.A1(new_n686), .A2(KEYINPUT104), .A3(new_n482), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n692), .B1(new_n677), .B2(new_n377), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n691), .B2(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1327gat));
  AOI21_X1  g497(.A(new_n669), .B1(new_n665), .B2(new_n666), .ZN(new_n699));
  INV_X1    g498(.A(new_n601), .ZN(new_n700));
  INV_X1    g499(.A(new_n629), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT105), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n562), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n678), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n704), .A2(G29gat), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT45), .Z(new_n707));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n514), .B2(new_n629), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n505), .A2(KEYINPUT86), .A3(new_n506), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT86), .B1(new_n505), .B2(new_n506), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n513), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT106), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n513), .B(new_n713), .C1(new_n709), .C2(new_n710), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n465), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n629), .B(KEYINPUT107), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT44), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n708), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n671), .A2(new_n561), .A3(new_n601), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n705), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n707), .A2(new_n721), .ZN(G1328gat));
  NOR3_X1   g521(.A1(new_n704), .A2(G36gat), .A3(new_n409), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT46), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n720), .B2(new_n409), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  OAI21_X1  g525(.A(G43gat), .B1(new_n720), .B2(new_n688), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT47), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n315), .A2(G43gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n704), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n729), .B(new_n731), .ZN(G1330gat));
  OAI21_X1  g531(.A(G50gat), .B1(new_n720), .B2(new_n482), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n482), .A2(G50gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT48), .Z(G1331gat));
  NOR2_X1   g538(.A1(new_n630), .A2(new_n631), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n561), .A3(new_n671), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n715), .A2(KEYINPUT110), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT110), .B1(new_n715), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n705), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(new_n573), .ZN(G1332gat));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n408), .A3(new_n743), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n744), .B2(new_n688), .ZN(new_n751));
  INV_X1    g550(.A(new_n315), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n563), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n751), .B(KEYINPUT50), .C1(new_n744), .C2(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1334gat));
  NOR2_X1   g557(.A1(new_n744), .A2(new_n482), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(new_n564), .ZN(G1335gat));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n699), .A2(new_n601), .A3(new_n560), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n718), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n718), .B2(new_n762), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n705), .ZN(new_n767));
  INV_X1    g566(.A(new_n715), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n601), .A2(new_n560), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n701), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT51), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n715), .A2(new_n773), .A3(new_n770), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n671), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n603), .A3(new_n678), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n767), .A2(new_n777), .ZN(G1336gat));
  AOI21_X1  g577(.A(new_n602), .B1(new_n765), .B2(new_n408), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n699), .A2(G92gat), .A3(new_n409), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT112), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n772), .B2(new_n774), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n784), .B(new_n781), .C1(new_n772), .C2(new_n774), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT52), .B1(new_n779), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n780), .B1(new_n772), .B2(new_n774), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n718), .A2(new_n762), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n409), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n788), .B(new_n789), .C1(new_n791), .C2(new_n602), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(new_n792), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n766), .B2(new_n688), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n607), .A3(new_n752), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1338gat));
  OAI21_X1  g595(.A(G106gat), .B1(new_n790), .B2(new_n482), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n377), .A2(new_n608), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n797), .B(new_n798), .C1(new_n775), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n775), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n765), .A2(new_n377), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(G106gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n803), .B2(new_n798), .ZN(G1339gat));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n629), .B(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n654), .A2(new_n659), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n668), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(KEYINPUT114), .A3(new_n668), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n658), .A2(new_n807), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n656), .A2(new_n655), .A3(new_n657), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n669), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n808), .A2(KEYINPUT114), .A3(new_n668), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT114), .B1(new_n808), .B2(new_n668), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n814), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n823), .A3(new_n560), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n543), .B1(new_n539), .B2(new_n541), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n548), .A2(new_n549), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n555), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n559), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n671), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n806), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n818), .A2(new_n823), .A3(new_n828), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n716), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n700), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n740), .A2(new_n561), .A3(new_n699), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n678), .A2(new_n409), .A3(new_n378), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n561), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(new_n257), .ZN(G1340gat));
  NOR2_X1   g638(.A1(new_n837), .A2(new_n699), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(new_n255), .ZN(G1341gat));
  INV_X1    g640(.A(new_n837), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n601), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n266), .A2(new_n268), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(G1342gat));
  AND2_X1   g644(.A1(new_n262), .A2(new_n263), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n701), .A2(new_n846), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n837), .A2(KEYINPUT56), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G134gat), .B1(new_n837), .B2(new_n629), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT56), .B1(new_n837), .B2(new_n847), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT115), .ZN(G1343gat));
  NOR3_X1   g651(.A1(new_n705), .A2(new_n408), .A3(new_n511), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT116), .ZN(new_n854));
  INV_X1    g653(.A(G141gat), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n561), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n835), .B2(new_n377), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  XNOR2_X1  g657(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n822), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n818), .A2(new_n860), .A3(new_n560), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n701), .B1(new_n861), .B2(new_n829), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n700), .B1(new_n862), .B2(new_n832), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n858), .B(new_n482), .C1(new_n863), .C2(new_n834), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n854), .B(new_n856), .C1(new_n857), .C2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n835), .A2(new_n377), .A3(new_n853), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n855), .B1(new_n866), .B2(new_n561), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(KEYINPUT58), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(KEYINPUT118), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(KEYINPUT118), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n865), .A2(new_n867), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI211_X1 g673(.A(KEYINPUT119), .B(KEYINPUT58), .C1(new_n865), .C2(new_n867), .ZN(new_n875));
  OAI22_X1  g674(.A1(new_n869), .A2(new_n870), .B1(new_n874), .B2(new_n875), .ZN(G1344gat));
  OR2_X1    g675(.A1(new_n857), .A2(new_n864), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n854), .A2(new_n671), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(KEYINPUT59), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT59), .B1(new_n866), .B2(new_n699), .ZN(new_n880));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n877), .A2(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n818), .A2(new_n823), .A3(new_n701), .A4(new_n828), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT121), .B1(new_n862), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(new_n560), .A3(new_n670), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n888), .A2(new_n860), .B1(new_n671), .B2(new_n828), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n886), .B(new_n883), .C1(new_n889), .C2(new_n701), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n885), .A2(new_n890), .A3(new_n700), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n834), .B(KEYINPUT120), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n377), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n858), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n482), .A2(new_n858), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n835), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n878), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n882), .B1(new_n899), .B2(new_n900), .ZN(G1345gat));
  NAND2_X1  g700(.A1(new_n877), .A2(new_n854), .ZN(new_n902));
  OAI21_X1  g701(.A(G155gat), .B1(new_n902), .B2(new_n700), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n601), .A2(new_n337), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n866), .B2(new_n904), .ZN(G1346gat));
  OAI21_X1  g704(.A(new_n338), .B1(new_n866), .B2(new_n629), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n806), .A2(G162gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT122), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n910), .B(new_n906), .C1(new_n902), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n678), .A2(new_n409), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n378), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n835), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n560), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(G169gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(G1348gat));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n671), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(G176gat), .ZN(G1349gat));
  NOR3_X1   g721(.A1(new_n915), .A2(new_n212), .A3(new_n700), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n916), .A2(new_n601), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n204), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g725(.A(new_n205), .B1(new_n916), .B2(new_n701), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT124), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(KEYINPUT124), .ZN(new_n929));
  XOR2_X1   g728(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n205), .A3(new_n806), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n927), .B(new_n933), .ZN(new_n934));
  OR2_X1    g733(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n931), .B(new_n932), .C1(new_n934), .C2(new_n935), .ZN(G1351gat));
  NOR3_X1   g735(.A1(new_n511), .A2(new_n482), .A3(new_n409), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n705), .B1(new_n937), .B2(KEYINPUT126), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n938), .B1(KEYINPUT126), .B2(new_n937), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n835), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n560), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n913), .A2(new_n688), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n942), .B1(new_n895), .B2(new_n898), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n560), .A2(G197gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(G204gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(new_n946), .A3(new_n671), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT62), .Z(new_n948));
  AND2_X1   g747(.A1(new_n943), .A2(new_n671), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n946), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n940), .A2(new_n323), .A3(new_n601), .ZN(new_n951));
  INV_X1    g750(.A(new_n942), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT57), .B1(new_n893), .B2(new_n377), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n601), .B(new_n952), .C1(new_n953), .C2(new_n897), .ZN(new_n954));
  OAI21_X1  g753(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n954), .B2(new_n956), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  NAND3_X1  g759(.A1(new_n940), .A2(new_n324), .A3(new_n806), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n943), .A2(new_n701), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n324), .ZN(G1355gat));
endmodule


