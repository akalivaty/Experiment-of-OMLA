

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U553 ( .A1(n715), .A2(n714), .ZN(n716) );
  BUF_X2 U554 ( .A(n657), .Z(n696) );
  NOR2_X2 U555 ( .A1(n592), .A2(n547), .ZN(n794) );
  NOR2_X1 U556 ( .A1(n968), .A2(n662), .ZN(n664) );
  INV_X1 U557 ( .A(KEYINPUT64), .ZN(n663) );
  XNOR2_X1 U558 ( .A(KEYINPUT66), .B(n521), .ZN(n523) );
  XOR2_X1 U559 ( .A(KEYINPUT95), .B(n691), .Z(n519) );
  OR2_X1 U560 ( .A1(n725), .A2(n734), .ZN(n520) );
  INV_X1 U561 ( .A(G8), .ZN(n687) );
  AND2_X1 U562 ( .A1(n980), .A2(n520), .ZN(n726) );
  INV_X1 U563 ( .A(KEYINPUT97), .ZN(n739) );
  NOR2_X1 U564 ( .A1(G2105), .A2(n528), .ZN(n533) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n635) );
  INV_X1 U566 ( .A(G2104), .ZN(n528) );
  XOR2_X1 U567 ( .A(G651), .B(KEYINPUT68), .Z(n547) );
  NOR2_X1 U568 ( .A1(n592), .A2(G651), .ZN(n798) );
  XNOR2_X1 U569 ( .A(n644), .B(KEYINPUT15), .ZN(n971) );
  NOR2_X1 U570 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U571 ( .A1(n656), .A2(n655), .ZN(n968) );
  NAND2_X1 U572 ( .A1(G101), .A2(n533), .ZN(n521) );
  INV_X1 U573 ( .A(KEYINPUT23), .ZN(n522) );
  XNOR2_X1 U574 ( .A(n523), .B(n522), .ZN(n526) );
  NAND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XNOR2_X1 U576 ( .A(n524), .B(KEYINPUT67), .ZN(n880) );
  NAND2_X1 U577 ( .A1(G113), .A2(n880), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X2 U580 ( .A(KEYINPUT17), .B(n527), .Z(n884) );
  NAND2_X1 U581 ( .A1(G137), .A2(n884), .ZN(n530) );
  AND2_X1 U582 ( .A1(n528), .A2(G2105), .ZN(n881) );
  NAND2_X1 U583 ( .A1(G125), .A2(n881), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X2 U585 ( .A1(n532), .A2(n531), .ZN(G160) );
  NAND2_X1 U586 ( .A1(G138), .A2(n884), .ZN(n536) );
  INV_X1 U587 ( .A(n533), .ZN(n534) );
  INV_X1 U588 ( .A(n534), .ZN(n885) );
  NAND2_X1 U589 ( .A1(G102), .A2(n885), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G114), .A2(n880), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G126), .A2(n881), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U594 ( .A1(n540), .A2(n539), .ZN(G164) );
  XOR2_X1 U595 ( .A(KEYINPUT0), .B(G543), .Z(n592) );
  NAND2_X1 U596 ( .A1(n798), .A2(G47), .ZN(n544) );
  XNOR2_X1 U597 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n542) );
  NOR2_X1 U598 ( .A1(G543), .A2(n547), .ZN(n541) );
  XNOR2_X2 U599 ( .A(n542), .B(n541), .ZN(n797) );
  NAND2_X1 U600 ( .A1(n797), .A2(G60), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U602 ( .A(KEYINPUT70), .B(n545), .Z(n551) );
  NOR2_X1 U603 ( .A1(G543), .A2(G651), .ZN(n546) );
  XOR2_X2 U604 ( .A(KEYINPUT65), .B(n546), .Z(n793) );
  NAND2_X1 U605 ( .A1(G85), .A2(n793), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G72), .A2(n794), .ZN(n548) );
  AND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(G290) );
  NAND2_X1 U609 ( .A1(G65), .A2(n797), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G53), .A2(n798), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U612 ( .A(KEYINPUT74), .B(n554), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G91), .A2(n793), .ZN(n555) );
  XNOR2_X1 U614 ( .A(KEYINPUT73), .B(n555), .ZN(n556) );
  NOR2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n794), .A2(G78), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(G299) );
  NAND2_X1 U618 ( .A1(G64), .A2(n797), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G52), .A2(n798), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n568) );
  XNOR2_X1 U621 ( .A(KEYINPUT9), .B(KEYINPUT72), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n793), .A2(G90), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n794), .A2(G77), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT71), .B(n562), .Z(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U626 ( .A(n566), .B(n565), .Z(n567) );
  NOR2_X1 U627 ( .A1(n568), .A2(n567), .ZN(G171) );
  NAND2_X1 U628 ( .A1(n793), .A2(G89), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n569), .B(KEYINPUT4), .ZN(n571) );
  NAND2_X1 U630 ( .A1(G76), .A2(n794), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U632 ( .A(n572), .B(KEYINPUT5), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G63), .A2(n797), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G51), .A2(n798), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT6), .B(n575), .Z(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U638 ( .A(n578), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U639 ( .A1(G62), .A2(n797), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G88), .A2(n793), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G50), .A2(n798), .ZN(n581) );
  XNOR2_X1 U643 ( .A(KEYINPUT83), .B(n581), .ZN(n582) );
  NOR2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n794), .A2(G75), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(G303) );
  XNOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .ZN(n586) );
  XNOR2_X1 U648 ( .A(n586), .B(KEYINPUT77), .ZN(G286) );
  NAND2_X1 U649 ( .A1(G651), .A2(G74), .ZN(n587) );
  XNOR2_X1 U650 ( .A(n587), .B(KEYINPUT80), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G49), .A2(n798), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U653 ( .A(KEYINPUT81), .B(n590), .Z(n591) );
  NOR2_X1 U654 ( .A1(n797), .A2(n591), .ZN(n594) );
  NAND2_X1 U655 ( .A1(n592), .A2(G87), .ZN(n593) );
  NAND2_X1 U656 ( .A1(n594), .A2(n593), .ZN(G288) );
  NAND2_X1 U657 ( .A1(G86), .A2(n793), .ZN(n601) );
  NAND2_X1 U658 ( .A1(G61), .A2(n797), .ZN(n596) );
  NAND2_X1 U659 ( .A1(G48), .A2(n798), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U661 ( .A1(n794), .A2(G73), .ZN(n597) );
  XOR2_X1 U662 ( .A(KEYINPUT2), .B(n597), .Z(n598) );
  NOR2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U664 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U665 ( .A(n602), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U666 ( .A1(G160), .A2(G40), .ZN(n634) );
  NOR2_X1 U667 ( .A1(n635), .A2(n634), .ZN(n754) );
  XNOR2_X1 U668 ( .A(G2067), .B(KEYINPUT37), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n603), .B(KEYINPUT88), .ZN(n744) );
  NAND2_X1 U670 ( .A1(G140), .A2(n884), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G104), .A2(n885), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U673 ( .A(KEYINPUT34), .B(n606), .ZN(n611) );
  NAND2_X1 U674 ( .A1(G116), .A2(n880), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G128), .A2(n881), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U677 ( .A(KEYINPUT35), .B(n609), .Z(n610) );
  NOR2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U679 ( .A(KEYINPUT36), .B(n612), .ZN(n899) );
  NOR2_X1 U680 ( .A1(n744), .A2(n899), .ZN(n930) );
  NAND2_X1 U681 ( .A1(n754), .A2(n930), .ZN(n750) );
  XNOR2_X1 U682 ( .A(G1986), .B(G290), .ZN(n970) );
  NAND2_X1 U683 ( .A1(n754), .A2(n970), .ZN(n613) );
  XNOR2_X1 U684 ( .A(KEYINPUT87), .B(n613), .ZN(n632) );
  NAND2_X1 U685 ( .A1(G131), .A2(n884), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G107), .A2(n880), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U688 ( .A1(G119), .A2(n881), .ZN(n616) );
  XNOR2_X1 U689 ( .A(KEYINPUT89), .B(n616), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n885), .A2(G95), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n866) );
  NAND2_X1 U693 ( .A1(G1991), .A2(n866), .ZN(n629) );
  NAND2_X1 U694 ( .A1(G141), .A2(n884), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G117), .A2(n880), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n885), .A2(G105), .ZN(n623) );
  XOR2_X1 U698 ( .A(KEYINPUT38), .B(n623), .Z(n624) );
  NOR2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n881), .A2(G129), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n867) );
  NAND2_X1 U702 ( .A1(G1996), .A2(n867), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n916) );
  NAND2_X1 U704 ( .A1(n916), .A2(n754), .ZN(n630) );
  XOR2_X1 U705 ( .A(n630), .B(KEYINPUT90), .Z(n631) );
  NOR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  AND2_X1 U707 ( .A1(n750), .A2(n633), .ZN(n742) );
  INV_X1 U708 ( .A(n634), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n657) );
  NAND2_X1 U710 ( .A1(G8), .A2(n657), .ZN(n734) );
  NAND2_X1 U711 ( .A1(G92), .A2(n793), .ZN(n643) );
  NAND2_X1 U712 ( .A1(G66), .A2(n797), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G54), .A2(n798), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n794), .A2(G79), .ZN(n639) );
  XOR2_X1 U716 ( .A(KEYINPUT76), .B(n639), .Z(n640) );
  NOR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  INV_X1 U719 ( .A(n971), .ZN(n780) );
  NAND2_X1 U720 ( .A1(G1348), .A2(n696), .ZN(n646) );
  INV_X1 U721 ( .A(n657), .ZN(n682) );
  NAND2_X1 U722 ( .A1(G2067), .A2(n682), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT93), .B(n647), .Z(n667) );
  OR2_X2 U725 ( .A1(n780), .A2(n667), .ZN(n666) );
  NAND2_X1 U726 ( .A1(G56), .A2(n797), .ZN(n648) );
  XOR2_X1 U727 ( .A(KEYINPUT14), .B(n648), .Z(n654) );
  NAND2_X1 U728 ( .A1(n793), .A2(G81), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(KEYINPUT12), .ZN(n651) );
  NAND2_X1 U730 ( .A1(G68), .A2(n794), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U732 ( .A(KEYINPUT13), .B(n652), .Z(n653) );
  NAND2_X1 U733 ( .A1(n798), .A2(G43), .ZN(n655) );
  INV_X1 U734 ( .A(G1996), .ZN(n945) );
  NOR2_X1 U735 ( .A1(n657), .A2(n945), .ZN(n659) );
  INV_X1 U736 ( .A(KEYINPUT26), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n659), .B(n658), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n696), .A2(G1341), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n666), .A2(n665), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n780), .A2(n667), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n670), .B(KEYINPUT94), .ZN(n675) );
  NAND2_X1 U745 ( .A1(n682), .A2(G2072), .ZN(n671) );
  XNOR2_X1 U746 ( .A(n671), .B(KEYINPUT27), .ZN(n673) );
  INV_X1 U747 ( .A(G1956), .ZN(n990) );
  NOR2_X1 U748 ( .A1(n990), .A2(n682), .ZN(n672) );
  NOR2_X1 U749 ( .A1(n673), .A2(n672), .ZN(n676) );
  INV_X1 U750 ( .A(G299), .ZN(n807) );
  NAND2_X1 U751 ( .A1(n676), .A2(n807), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U753 ( .A1(n676), .A2(n807), .ZN(n677) );
  XOR2_X1 U754 ( .A(n677), .B(KEYINPUT28), .Z(n678) );
  NAND2_X1 U755 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U756 ( .A(KEYINPUT29), .B(n680), .Z(n686) );
  OR2_X1 U757 ( .A1(n682), .A2(G1961), .ZN(n684) );
  XNOR2_X1 U758 ( .A(G2078), .B(KEYINPUT25), .ZN(n681) );
  XNOR2_X1 U759 ( .A(n681), .B(KEYINPUT92), .ZN(n948) );
  NAND2_X1 U760 ( .A1(n682), .A2(n948), .ZN(n683) );
  NAND2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n692), .A2(G171), .ZN(n685) );
  NAND2_X1 U763 ( .A1(n686), .A2(n685), .ZN(n709) );
  NOR2_X1 U764 ( .A1(G1966), .A2(n734), .ZN(n712) );
  INV_X1 U765 ( .A(n712), .ZN(n689) );
  NOR2_X1 U766 ( .A1(n696), .A2(G2084), .ZN(n710) );
  NOR2_X1 U767 ( .A1(n710), .A2(n687), .ZN(n688) );
  NAND2_X1 U768 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U769 ( .A(KEYINPUT30), .B(n690), .ZN(n691) );
  NOR2_X1 U770 ( .A1(G168), .A2(n519), .ZN(n694) );
  NOR2_X1 U771 ( .A1(G171), .A2(n692), .ZN(n693) );
  NOR2_X1 U772 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U773 ( .A(KEYINPUT31), .B(n695), .Z(n708) );
  NOR2_X1 U774 ( .A1(G1971), .A2(n734), .ZN(n698) );
  NOR2_X1 U775 ( .A1(G2090), .A2(n696), .ZN(n697) );
  NOR2_X1 U776 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U777 ( .A1(n699), .A2(G303), .ZN(n700) );
  OR2_X1 U778 ( .A1(n687), .A2(n700), .ZN(n702) );
  AND2_X1 U779 ( .A1(n708), .A2(n702), .ZN(n701) );
  NAND2_X1 U780 ( .A1(n709), .A2(n701), .ZN(n706) );
  INV_X1 U781 ( .A(n702), .ZN(n704) );
  AND2_X1 U782 ( .A1(G286), .A2(G8), .ZN(n703) );
  OR2_X1 U783 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U784 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U785 ( .A(n707), .B(KEYINPUT32), .ZN(n717) );
  AND2_X1 U786 ( .A1(n709), .A2(n708), .ZN(n715) );
  NAND2_X1 U787 ( .A1(G8), .A2(n710), .ZN(n711) );
  XNOR2_X1 U788 ( .A(KEYINPUT91), .B(n711), .ZN(n713) );
  OR2_X1 U789 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U790 ( .A1(n717), .A2(n716), .ZN(n728) );
  NOR2_X1 U791 ( .A1(G1976), .A2(G288), .ZN(n724) );
  NOR2_X1 U792 ( .A1(G1971), .A2(G303), .ZN(n718) );
  NOR2_X1 U793 ( .A1(n724), .A2(n718), .ZN(n975) );
  NAND2_X1 U794 ( .A1(n728), .A2(n975), .ZN(n719) );
  NAND2_X1 U795 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NAND2_X1 U796 ( .A1(n719), .A2(n974), .ZN(n720) );
  XNOR2_X1 U797 ( .A(KEYINPUT96), .B(n720), .ZN(n721) );
  NOR2_X1 U798 ( .A1(n734), .A2(n721), .ZN(n722) );
  NOR2_X1 U799 ( .A1(n722), .A2(KEYINPUT33), .ZN(n723) );
  INV_X1 U800 ( .A(n723), .ZN(n727) );
  XOR2_X1 U801 ( .A(G1981), .B(G305), .Z(n980) );
  NAND2_X1 U802 ( .A1(n724), .A2(KEYINPUT33), .ZN(n725) );
  NAND2_X1 U803 ( .A1(n727), .A2(n726), .ZN(n738) );
  NOR2_X1 U804 ( .A1(G2090), .A2(G303), .ZN(n729) );
  NAND2_X1 U805 ( .A1(G8), .A2(n729), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n728), .A2(n730), .ZN(n731) );
  AND2_X1 U807 ( .A1(n731), .A2(n734), .ZN(n736) );
  NOR2_X1 U808 ( .A1(G1981), .A2(G305), .ZN(n732) );
  XOR2_X1 U809 ( .A(n732), .B(KEYINPUT24), .Z(n733) );
  NOR2_X1 U810 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U813 ( .A(n740), .B(n739), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U815 ( .A(n743), .B(KEYINPUT98), .ZN(n757) );
  NAND2_X1 U816 ( .A1(n744), .A2(n899), .ZN(n917) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n867), .ZN(n920) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n866), .ZN(n927) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n927), .A2(n745), .ZN(n746) );
  XOR2_X1 U821 ( .A(KEYINPUT99), .B(n746), .Z(n747) );
  NOR2_X1 U822 ( .A1(n916), .A2(n747), .ZN(n748) );
  NOR2_X1 U823 ( .A1(n920), .A2(n748), .ZN(n749) );
  XNOR2_X1 U824 ( .A(n749), .B(KEYINPUT39), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n917), .A2(n752), .ZN(n753) );
  XNOR2_X1 U827 ( .A(KEYINPUT100), .B(n753), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U829 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U830 ( .A(n758), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U831 ( .A(G2435), .B(G2454), .Z(n760) );
  XNOR2_X1 U832 ( .A(G2430), .B(G2438), .ZN(n759) );
  XNOR2_X1 U833 ( .A(n760), .B(n759), .ZN(n767) );
  XOR2_X1 U834 ( .A(G2446), .B(KEYINPUT101), .Z(n762) );
  XNOR2_X1 U835 ( .A(G2451), .B(G2443), .ZN(n761) );
  XNOR2_X1 U836 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U837 ( .A(n763), .B(G2427), .Z(n765) );
  XNOR2_X1 U838 ( .A(G1341), .B(G1348), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n765), .B(n764), .ZN(n766) );
  XNOR2_X1 U840 ( .A(n767), .B(n766), .ZN(n768) );
  AND2_X1 U841 ( .A1(n768), .A2(G14), .ZN(G401) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U843 ( .A1(G135), .A2(n884), .ZN(n770) );
  NAND2_X1 U844 ( .A1(G111), .A2(n880), .ZN(n769) );
  NAND2_X1 U845 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U846 ( .A1(n881), .A2(G123), .ZN(n771) );
  XOR2_X1 U847 ( .A(KEYINPUT18), .B(n771), .Z(n772) );
  NOR2_X1 U848 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U849 ( .A1(n885), .A2(G99), .ZN(n774) );
  NAND2_X1 U850 ( .A1(n775), .A2(n774), .ZN(n928) );
  XNOR2_X1 U851 ( .A(G2096), .B(n928), .ZN(n776) );
  OR2_X1 U852 ( .A1(G2100), .A2(n776), .ZN(G156) );
  INV_X1 U853 ( .A(G132), .ZN(G219) );
  INV_X1 U854 ( .A(G82), .ZN(G220) );
  INV_X1 U855 ( .A(G120), .ZN(G236) );
  NAND2_X1 U856 ( .A1(G7), .A2(G661), .ZN(n777) );
  XNOR2_X1 U857 ( .A(n777), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U858 ( .A(G223), .ZN(n832) );
  NAND2_X1 U859 ( .A1(n832), .A2(G567), .ZN(n778) );
  XNOR2_X1 U860 ( .A(n778), .B(KEYINPUT75), .ZN(n779) );
  XNOR2_X1 U861 ( .A(KEYINPUT11), .B(n779), .ZN(G234) );
  INV_X1 U862 ( .A(G860), .ZN(n785) );
  OR2_X1 U863 ( .A1(n968), .A2(n785), .ZN(G153) );
  INV_X1 U864 ( .A(G171), .ZN(G301) );
  NAND2_X1 U865 ( .A1(G868), .A2(G301), .ZN(n782) );
  INV_X1 U866 ( .A(G868), .ZN(n815) );
  NAND2_X1 U867 ( .A1(n780), .A2(n815), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(G284) );
  NOR2_X1 U869 ( .A1(G286), .A2(n815), .ZN(n784) );
  NOR2_X1 U870 ( .A1(G868), .A2(G299), .ZN(n783) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(G297) );
  NAND2_X1 U872 ( .A1(n785), .A2(G559), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n786), .A2(n971), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U875 ( .A1(n971), .A2(G868), .ZN(n788) );
  NOR2_X1 U876 ( .A1(G559), .A2(n788), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n789), .B(KEYINPUT78), .ZN(n791) );
  NOR2_X1 U878 ( .A1(n968), .A2(G868), .ZN(n790) );
  NOR2_X1 U879 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U880 ( .A1(G559), .A2(n971), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n792), .B(n968), .ZN(n811) );
  NOR2_X1 U882 ( .A1(n811), .A2(G860), .ZN(n804) );
  NAND2_X1 U883 ( .A1(G93), .A2(n793), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G80), .A2(n794), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n803) );
  NAND2_X1 U886 ( .A1(G67), .A2(n797), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U889 ( .A(KEYINPUT79), .B(n801), .Z(n802) );
  OR2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n814) );
  XOR2_X1 U891 ( .A(n804), .B(n814), .Z(G145) );
  INV_X1 U892 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U893 ( .A(G305), .B(n814), .ZN(n805) );
  XNOR2_X1 U894 ( .A(G288), .B(n805), .ZN(n806) );
  XOR2_X1 U895 ( .A(n806), .B(KEYINPUT19), .Z(n809) );
  XNOR2_X1 U896 ( .A(n807), .B(G166), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n809), .B(n808), .ZN(n810) );
  XNOR2_X1 U898 ( .A(n810), .B(G290), .ZN(n903) );
  XNOR2_X1 U899 ( .A(KEYINPUT84), .B(n811), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n903), .B(n812), .ZN(n813) );
  NAND2_X1 U901 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U902 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U903 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U904 ( .A1(G2078), .A2(G2084), .ZN(n818) );
  XOR2_X1 U905 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U906 ( .A1(G2090), .A2(n819), .ZN(n820) );
  XNOR2_X1 U907 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U908 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XOR2_X1 U909 ( .A(KEYINPUT85), .B(G44), .Z(n822) );
  XNOR2_X1 U910 ( .A(KEYINPUT3), .B(n822), .ZN(G218) );
  NAND2_X1 U911 ( .A1(G69), .A2(G57), .ZN(n823) );
  NOR2_X1 U912 ( .A1(G236), .A2(n823), .ZN(n824) );
  XNOR2_X1 U913 ( .A(KEYINPUT86), .B(n824), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n825), .A2(G108), .ZN(n836) );
  NAND2_X1 U915 ( .A1(G567), .A2(n836), .ZN(n830) );
  NOR2_X1 U916 ( .A1(G220), .A2(G219), .ZN(n826) );
  XOR2_X1 U917 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U918 ( .A1(G218), .A2(n827), .ZN(n828) );
  NAND2_X1 U919 ( .A1(G96), .A2(n828), .ZN(n837) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n837), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n830), .A2(n829), .ZN(n838) );
  NAND2_X1 U922 ( .A1(G483), .A2(G661), .ZN(n831) );
  NOR2_X1 U923 ( .A1(n838), .A2(n831), .ZN(n835) );
  NAND2_X1 U924 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U927 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G188) );
  XOR2_X1 U930 ( .A(G69), .B(KEYINPUT102), .Z(G235) );
  INV_X1 U932 ( .A(G108), .ZN(G238) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G57), .ZN(G237) );
  NOR2_X1 U935 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U937 ( .A(KEYINPUT103), .B(n838), .ZN(G319) );
  XOR2_X1 U938 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n840) );
  XNOR2_X1 U939 ( .A(G2678), .B(KEYINPUT105), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U941 ( .A(KEYINPUT104), .B(G2090), .Z(n842) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U945 ( .A(G2096), .B(G2100), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U947 ( .A(G2078), .B(G2084), .Z(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1976), .B(G1981), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1971), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n851), .B(G2474), .Z(n853) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1956), .Z(n855) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1961), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U959 ( .A1(n885), .A2(G100), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G136), .A2(n884), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G112), .A2(n880), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n881), .A2(G124), .ZN(n860) );
  XOR2_X1 U964 ( .A(KEYINPUT44), .B(n860), .Z(n861) );
  NOR2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U967 ( .A(KEYINPUT106), .B(n865), .Z(G162) );
  XOR2_X1 U968 ( .A(n867), .B(n866), .Z(n868) );
  XNOR2_X1 U969 ( .A(n928), .B(n868), .ZN(n869) );
  XNOR2_X1 U970 ( .A(G162), .B(n869), .ZN(n879) );
  NAND2_X1 U971 ( .A1(G139), .A2(n884), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G103), .A2(n885), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G115), .A2(n880), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G127), .A2(n881), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT110), .B(n875), .ZN(n876) );
  NOR2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n935) );
  XNOR2_X1 U980 ( .A(G164), .B(n935), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n901) );
  XOR2_X1 U982 ( .A(KEYINPUT111), .B(KEYINPUT109), .Z(n894) );
  NAND2_X1 U983 ( .A1(G118), .A2(n880), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G130), .A2(n881), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G142), .A2(n884), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G106), .A2(n885), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U989 ( .A(KEYINPUT107), .B(n888), .ZN(n889) );
  XNOR2_X1 U990 ( .A(KEYINPUT45), .B(n889), .ZN(n890) );
  NOR2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n892), .B(KEYINPUT46), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U994 ( .A(n895), .B(KEYINPUT108), .Z(n897) );
  XNOR2_X1 U995 ( .A(G160), .B(KEYINPUT48), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U1000 ( .A(n903), .B(G286), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G171), .B(n971), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n906), .B(n968), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n912), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(KEYINPUT114), .B(n913), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(n916), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n925) );
  XOR2_X1 U1017 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n923) );
  XOR2_X1 U1018 ( .A(G2090), .B(KEYINPUT116), .Z(n919) );
  XNOR2_X1 U1019 ( .A(G162), .B(n919), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n934) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1027 ( .A(KEYINPUT115), .B(n932), .Z(n933) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1029 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n1021) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n1021), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n943), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1038 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n957) );
  XNOR2_X1 U1039 ( .A(KEYINPUT119), .B(G2072), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n944), .B(G33), .ZN(n952) );
  XOR2_X1 U1041 ( .A(G2067), .B(G26), .Z(n947) );
  XNOR2_X1 U1042 ( .A(n945), .B(G32), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1044 ( .A(n948), .B(G27), .Z(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1047 ( .A(G1991), .B(G25), .Z(n953) );
  NAND2_X1 U1048 ( .A1(G28), .A2(n953), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n957), .B(n956), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(G2084), .B(G34), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n958), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G2090), .B(G35), .Z(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT118), .B(n961), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n1022) );
  NOR2_X1 U1057 ( .A1(G29), .A2(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n1022), .A2(n964), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n965), .ZN(n1026) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n989) );
  XNOR2_X1 U1061 ( .A(G301), .B(G1961), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(G299), .B(G1956), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n987) );
  XNOR2_X1 U1064 ( .A(G1341), .B(n968), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n979) );
  XNOR2_X1 U1066 ( .A(n971), .B(G1348), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(G1971), .A2(G303), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n985) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(n982), .B(KEYINPUT57), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n983), .B(KEYINPUT121), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n1019) );
  INV_X1 U1079 ( .A(G16), .ZN(n1017) );
  XNOR2_X1 U1080 ( .A(KEYINPUT126), .B(KEYINPUT125), .ZN(n1003) );
  XNOR2_X1 U1081 ( .A(n990), .B(G20), .ZN(n1000) );
  XOR2_X1 U1082 ( .A(KEYINPUT124), .B(G4), .Z(n992) );
  XNOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n992), .B(n991), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G1341), .B(G19), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(KEYINPUT122), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(G6), .B(G1981), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(n996), .B(KEYINPUT123), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT60), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1003), .B(n1002), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G21), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(G1961), .B(G5), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1986), .B(G24), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1101 ( .A(G1976), .B(G23), .Z(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(n1020), .B(KEYINPUT127), .ZN(n1024) );
  OR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

