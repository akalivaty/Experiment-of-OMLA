//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G68), .B2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n202), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n205), .A2(new_n224), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n221), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G58), .A2(G232), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n210), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n210), .A2(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n212), .B(new_n231), .C1(new_n214), .C2(new_n218), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT0), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n234), .A2(new_n209), .A3(new_n235), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n229), .A2(new_n233), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n220), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n202), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  OAI21_X1  g0053(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  OAI211_X1 g0059(.A(G1), .B(G13), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n254), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G238), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G97), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI211_X1 g0067(.A(G232), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(G226), .B1(new_n266), .B2(new_n267), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT70), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n258), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT65), .B(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .A4(G226), .ZN(new_n281));
  AOI211_X1 g0081(.A(new_n265), .B(new_n269), .C1(new_n274), .C2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n257), .B(new_n263), .C1(new_n282), .C2(new_n260), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT72), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n274), .A2(new_n281), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(new_n264), .A3(new_n268), .ZN(new_n288));
  INV_X1    g0088(.A(new_n260), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n284), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n290), .A2(new_n257), .A3(new_n291), .A4(new_n263), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n285), .A2(new_n286), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n283), .A2(KEYINPUT72), .A3(new_n284), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G169), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT14), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT13), .B1(new_n283), .B2(KEYINPUT73), .ZN(new_n298));
  OAI211_X1 g0098(.A(G179), .B(new_n292), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT14), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n293), .A2(new_n300), .A3(G169), .A4(new_n294), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n296), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n235), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n209), .A2(G33), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT66), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n307), .A2(new_n205), .B1(new_n209), .B2(G68), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G20), .A2(G33), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n202), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n304), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(new_n312), .B(KEYINPUT11), .Z(new_n313));
  AOI21_X1  g0113(.A(new_n304), .B1(new_n208), .B2(G20), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G68), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n230), .A2(new_n209), .A3(G1), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n316), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT12), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n313), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n302), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n293), .A2(G200), .A3(new_n294), .ZN(new_n325));
  OAI211_X1 g0125(.A(G190), .B(new_n292), .C1(new_n297), .C2(new_n298), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(new_n322), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n256), .B1(new_n262), .B2(G244), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT69), .ZN(new_n329));
  AND2_X1   g0129(.A1(G238), .A2(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n266), .A2(new_n267), .ZN(new_n331));
  AOI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(G232), .C2(new_n279), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n289), .B1(new_n278), .B2(G107), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n329), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G20), .A2(G77), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT8), .B(G58), .ZN(new_n337));
  XOR2_X1   g0137(.A(KEYINPUT15), .B(G87), .Z(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n336), .B1(new_n337), .B2(new_n310), .C1(new_n307), .C2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(new_n304), .B1(new_n205), .B2(new_n318), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n314), .A2(G77), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n335), .B(new_n344), .C1(new_n345), .C2(new_n334), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n324), .A2(new_n327), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n309), .A2(G150), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n348), .B1(new_n307), .B2(new_n337), .C1(new_n204), .C2(new_n209), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n304), .B1(new_n202), .B2(new_n318), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT67), .ZN(new_n352));
  INV_X1    g0152(.A(new_n304), .ZN(new_n353));
  INV_X1    g0153(.A(new_n318), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(KEYINPUT67), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G223), .ZN(new_n358));
  INV_X1    g0158(.A(G1698), .ZN(new_n359));
  INV_X1    g0159(.A(G222), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n278), .B1(new_n358), .B2(new_n359), .C1(new_n273), .C2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n289), .C1(G77), .C2(new_n278), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n257), .C1(new_n222), .C2(new_n261), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n357), .B(new_n365), .C1(G179), .C2(new_n363), .ZN(new_n366));
  XOR2_X1   g0166(.A(new_n366), .B(KEYINPUT68), .Z(new_n367));
  OR2_X1    g0167(.A1(new_n334), .A2(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n334), .A2(new_n364), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n367), .B1(new_n343), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(G200), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT9), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n372), .B1(new_n345), .B2(new_n363), .C1(new_n357), .C2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n373), .B2(new_n357), .ZN(new_n375));
  XOR2_X1   g0175(.A(new_n375), .B(KEYINPUT10), .Z(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n379), .A2(new_n380), .A3(new_n258), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n267), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n279), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n256), .B1(new_n384), .B2(new_n289), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n262), .A2(G232), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT76), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n378), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n273), .A2(new_n358), .B1(new_n222), .B2(new_n359), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT74), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n275), .ZN(new_n391));
  NAND2_X1  g0191(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(G33), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n276), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n386), .B(new_n257), .C1(new_n395), .C2(new_n260), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n377), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n396), .A2(G190), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n337), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n318), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n315), .B2(new_n403), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n248), .A2(new_n316), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n406), .B2(new_n201), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n309), .A2(G159), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n393), .A2(new_n209), .A3(new_n276), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n316), .B1(new_n410), .B2(KEYINPUT7), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n393), .A2(new_n412), .A3(new_n209), .A4(new_n276), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n409), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n353), .B1(new_n414), .B2(KEYINPUT16), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n258), .B1(new_n379), .B2(new_n380), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n418), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n277), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n412), .B1(new_n278), .B2(G20), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n316), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n417), .B1(new_n421), .B2(new_n409), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n405), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n402), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n396), .A2(new_n397), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n384), .A2(new_n289), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n426), .A2(KEYINPUT76), .A3(new_n257), .A4(new_n386), .ZN(new_n427));
  AOI21_X1  g0227(.A(G200), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(KEYINPUT77), .B(new_n423), .C1(new_n428), .C2(new_n400), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n396), .A2(G179), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n425), .A2(new_n427), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n364), .ZN(new_n434));
  INV_X1    g0234(.A(new_n423), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n434), .A2(KEYINPUT18), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT18), .B1(new_n434), .B2(new_n435), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n424), .B(new_n431), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n347), .A2(new_n371), .A3(new_n376), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT21), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT78), .ZN(new_n444));
  OAI21_X1  g0244(.A(G274), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT5), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(KEYINPUT78), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n208), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n449));
  OR3_X1    g0249(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n260), .B(G270), .C1(new_n449), .C2(new_n447), .ZN(new_n451));
  INV_X1    g0251(.A(G303), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n278), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G264), .A2(G1698), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n273), .B2(new_n214), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n455), .B2(new_n394), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n450), .B(new_n451), .C1(new_n456), .C2(new_n260), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n208), .A2(G33), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n354), .A2(G116), .A3(new_n353), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n318), .A2(new_n219), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n303), .A2(new_n235), .B1(G20), .B2(new_n219), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(new_n209), .C1(G33), .C2(new_n213), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT20), .B1(new_n462), .B2(new_n464), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n460), .B(new_n461), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G169), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n442), .B1(new_n458), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n458), .A2(G179), .A3(new_n467), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n457), .A2(KEYINPUT21), .A3(G169), .A4(new_n467), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n467), .B1(new_n457), .B2(G200), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(KEYINPUT84), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT84), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n475), .B(new_n467), .C1(new_n457), .C2(G200), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n458), .A2(G190), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n211), .A2(G20), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT22), .B1(new_n278), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n480), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n393), .B2(new_n276), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n481), .B1(new_n483), .B2(KEYINPUT22), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n209), .A2(G107), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT23), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n258), .A2(new_n219), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n209), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n490), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n484), .A2(new_n492), .A3(new_n486), .A4(new_n488), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n304), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n354), .A2(new_n353), .A3(new_n459), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G107), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n318), .A2(new_n217), .ZN(new_n497));
  XOR2_X1   g0297(.A(new_n497), .B(KEYINPUT25), .Z(new_n498));
  AND3_X1   g0298(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  INV_X1    g0300(.A(G294), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n258), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(G250), .B1(new_n271), .B2(new_n272), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G257), .A2(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(new_n394), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n500), .B1(new_n506), .B2(new_n260), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n503), .A2(new_n504), .B1(new_n393), .B2(new_n276), .ZN(new_n508));
  OAI211_X1 g0308(.A(KEYINPUT86), .B(new_n289), .C1(new_n508), .C2(new_n502), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n260), .B(G264), .C1(new_n449), .C2(new_n447), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n507), .A2(new_n450), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT88), .B1(new_n511), .B2(G190), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n509), .A2(new_n450), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT88), .ZN(new_n514));
  INV_X1    g0314(.A(new_n510), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n289), .B1(new_n508), .B2(new_n502), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n500), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(new_n514), .A3(new_n517), .A4(new_n345), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n510), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT87), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT87), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n516), .A2(new_n522), .A3(new_n510), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(G200), .B1(new_n524), .B2(new_n450), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n499), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n527));
  INV_X1    g0327(.A(G179), .ZN(new_n528));
  INV_X1    g0328(.A(new_n450), .ZN(new_n529));
  AOI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n521), .C2(new_n523), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n364), .B1(new_n513), .B2(new_n517), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n479), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(G238), .B(new_n279), .C1(new_n381), .C2(new_n267), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n224), .B1(new_n393), .B2(new_n276), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n487), .B1(new_n536), .B2(G1698), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT80), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n394), .A2(new_n538), .A3(G238), .A4(new_n279), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n289), .ZN(new_n541));
  INV_X1    g0341(.A(G45), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n212), .B1(new_n542), .B2(G1), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n208), .A2(new_n255), .A3(G45), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n260), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT81), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n541), .A2(KEYINPUT81), .A3(new_n546), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n364), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT81), .B1(new_n541), .B2(new_n546), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n548), .B(new_n545), .C1(new_n540), .C2(new_n289), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n528), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n307), .B2(new_n213), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n209), .B1(new_n264), .B2(new_n555), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT82), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n211), .A2(new_n213), .A3(new_n217), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n394), .A2(new_n209), .A3(G68), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n556), .A2(new_n562), .A3(KEYINPUT83), .A4(new_n563), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n304), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n495), .A2(new_n338), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n339), .A2(new_n318), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n551), .A2(new_n554), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n549), .A2(G200), .A3(new_n550), .ZN(new_n573));
  OAI21_X1  g0373(.A(G190), .B1(new_n552), .B2(new_n553), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n495), .A2(G87), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n568), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(KEYINPUT4), .B(G244), .C1(new_n271), .C2(new_n272), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G250), .A2(G1698), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n331), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(new_n279), .C1(new_n381), .C2(new_n267), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n260), .B1(new_n584), .B2(new_n463), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n260), .B(G257), .C1(new_n449), .C2(new_n447), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n450), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n364), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n318), .A2(new_n213), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n495), .A2(G97), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n217), .B1(new_n419), .B2(new_n420), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n310), .A2(new_n205), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT6), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n213), .A2(new_n217), .ZN(new_n594));
  NOR2_X1   g0394(.A1(G97), .A2(G107), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n209), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n591), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n589), .B(new_n590), .C1(new_n599), .C2(new_n353), .ZN(new_n600));
  INV_X1    g0400(.A(new_n587), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT4), .B1(new_n536), .B2(new_n279), .ZN(new_n602));
  INV_X1    g0402(.A(new_n463), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n602), .A2(new_n603), .A3(new_n581), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n528), .B(new_n601), .C1(new_n604), .C2(new_n260), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n588), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT79), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n588), .A2(new_n600), .A3(new_n605), .A4(KEYINPUT79), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n585), .A2(new_n587), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G190), .ZN(new_n612));
  INV_X1    g0412(.A(new_n600), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n601), .B1(new_n604), .B2(new_n260), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n533), .A2(new_n578), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n441), .A2(new_n618), .ZN(G372));
  INV_X1    g0419(.A(new_n367), .ZN(new_n620));
  INV_X1    g0420(.A(new_n437), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT18), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n327), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n370), .A2(new_n343), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n324), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n429), .B(KEYINPUT17), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n376), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n620), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n547), .A2(G200), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT89), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT89), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n547), .A2(new_n635), .A3(G200), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n574), .A2(new_n634), .A3(new_n576), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n547), .A2(new_n364), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n554), .A2(new_n571), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n612), .A2(new_n615), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n608), .A2(new_n609), .B1(new_n641), .B2(new_n613), .ZN(new_n642));
  INV_X1    g0442(.A(new_n472), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n532), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n640), .A2(new_n642), .A3(new_n526), .A4(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(new_n606), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n637), .A2(new_n646), .A3(new_n639), .A4(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT26), .B1(new_n578), .B2(new_n610), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n645), .A2(new_n639), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n441), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n632), .A2(new_n651), .ZN(G369));
  NOR2_X1   g0452(.A1(new_n230), .A2(G20), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OR3_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .A3(G1), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT27), .B1(new_n654), .B2(G1), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n526), .B(new_n532), .C1(new_n499), .C2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n532), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n643), .A2(new_n659), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n659), .A2(new_n467), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n479), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n643), .B2(new_n665), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT90), .B(G330), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n663), .A2(new_n526), .A3(new_n532), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n532), .B2(new_n659), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT91), .Z(G399));
  NOR2_X1   g0475(.A1(new_n231), .A2(G41), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT92), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n560), .A2(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n234), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n279), .A2(G257), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n682), .A2(new_n454), .B1(new_n276), .B2(new_n393), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n289), .B1(new_n683), .B2(new_n453), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(G179), .A3(new_n450), .A4(new_n451), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n521), .B2(new_n523), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n611), .B(new_n686), .C1(new_n552), .C2(new_n553), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n614), .A2(new_n528), .A3(new_n457), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n529), .B1(new_n521), .B2(new_n523), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n688), .A2(new_n687), .B1(new_n692), .B2(new_n547), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n689), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n547), .ZN(new_n696));
  INV_X1    g0496(.A(new_n687), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(KEYINPUT30), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT93), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n618), .B2(new_n660), .ZN(new_n703));
  INV_X1    g0503(.A(new_n689), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n660), .B1(new_n704), .B2(new_n693), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n701), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n668), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n637), .A2(new_n639), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT26), .B1(new_n709), .B2(new_n606), .ZN(new_n710));
  INV_X1    g0510(.A(new_n610), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n646), .A3(new_n572), .A4(new_n577), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n644), .A2(new_n610), .A3(new_n616), .A4(new_n526), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n639), .B1(new_n714), .B2(new_n709), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n660), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n650), .A2(new_n718), .A3(new_n660), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n708), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n681), .B1(new_n721), .B2(G1), .ZN(G364));
  AOI21_X1  g0522(.A(new_n208), .B1(new_n653), .B2(G45), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n677), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n670), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n668), .B2(new_n667), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n235), .B1(G20), .B2(new_n364), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n209), .A2(G179), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G190), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G159), .ZN(new_n734));
  XOR2_X1   g0534(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n209), .A2(new_n528), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT95), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT95), .B1(new_n209), .B2(new_n528), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n345), .A2(G200), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n345), .A2(new_n377), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n730), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n736), .B1(new_n248), .B2(new_n742), .C1(new_n211), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n734), .A2(new_n735), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n741), .A2(new_n528), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n213), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n377), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n730), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n278), .B1(new_n752), .B2(new_n217), .ZN(new_n753));
  OR3_X1    g0553(.A1(new_n746), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n737), .A2(new_n743), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n745), .B(new_n754), .C1(G50), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n737), .A2(new_n751), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n739), .A2(new_n731), .A3(new_n740), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n757), .B1(new_n316), .B2(new_n758), .C1(new_n205), .C2(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G326), .A2(new_n756), .B1(new_n748), .B2(G294), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n759), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT97), .ZN(new_n764));
  INV_X1    g0564(.A(new_n758), .ZN(new_n765));
  INV_X1    g0565(.A(G317), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT33), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n766), .A2(KEYINPUT33), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n752), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G283), .ZN(new_n771));
  INV_X1    g0571(.A(G329), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n331), .B1(new_n732), .B2(new_n772), .C1(new_n452), .C2(new_n744), .ZN(new_n773));
  INV_X1    g0573(.A(new_n742), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(G322), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n764), .A2(new_n769), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n729), .B1(new_n760), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n230), .A2(new_n258), .A3(KEYINPUT94), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT94), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G13), .B2(G33), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n728), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n249), .A2(G45), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n394), .A2(new_n231), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n234), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n787), .B1(new_n542), .B2(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n785), .A2(new_n789), .B1(new_n219), .B2(new_n231), .ZN(new_n790));
  INV_X1    g0590(.A(new_n231), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G355), .A3(new_n278), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n724), .B(new_n777), .C1(new_n784), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n783), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n667), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n727), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  NAND2_X1  g0598(.A1(new_n650), .A2(new_n660), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n346), .B1(new_n344), .B2(new_n660), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n626), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n370), .A2(new_n343), .A3(new_n660), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n799), .B(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(new_n707), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n724), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n774), .A2(G143), .B1(G150), .B2(new_n765), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n755), .C1(new_n809), .C2(new_n759), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  NOR2_X1   g0611(.A1(new_n752), .A2(new_n316), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n733), .A2(G132), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n811), .A2(new_n382), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n814), .B1(new_n202), .B2(new_n744), .C1(new_n248), .C2(new_n749), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n752), .A2(new_n211), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT98), .B(G283), .Z(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n758), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n750), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n744), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G107), .A2(new_n821), .B1(new_n733), .B2(G311), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n278), .B1(new_n756), .B2(G303), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n219), .B2(new_n759), .C1(new_n501), .C2(new_n742), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n815), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n724), .B1(new_n826), .B2(new_n728), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n781), .A2(new_n728), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n827), .B1(G77), .B2(new_n829), .C1(new_n782), .C2(new_n803), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n806), .A2(new_n830), .ZN(G384));
  AND2_X1   g0631(.A1(new_n596), .A2(new_n597), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT35), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n209), .B(new_n235), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n834), .B(G116), .C1(new_n833), .C2(new_n832), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT36), .ZN(new_n836));
  OAI21_X1  g0636(.A(G77), .B1(new_n248), .B2(new_n316), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n234), .B1(G50), .B2(new_n316), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(G1), .A3(new_n230), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT99), .ZN(new_n841));
  INV_X1    g0641(.A(new_n657), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT101), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n411), .A2(new_n413), .ZN(new_n844));
  INV_X1    g0644(.A(new_n409), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n844), .A2(KEYINPUT16), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n304), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT100), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT100), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n416), .B1(new_n414), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n843), .B1(new_n852), .B2(new_n405), .ZN(new_n853));
  INV_X1    g0653(.A(new_n405), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n849), .A2(new_n851), .ZN(new_n855));
  OAI211_X1 g0655(.A(KEYINPUT101), .B(new_n854), .C1(new_n855), .C2(new_n847), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n438), .A2(new_n842), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  AOI21_X1  g0659(.A(G169), .B1(new_n425), .B2(new_n427), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n657), .B1(new_n860), .B2(new_n432), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n853), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n402), .A2(new_n423), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n435), .B1(new_n434), .B2(new_n842), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n865), .A2(new_n863), .A3(new_n859), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n858), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n866), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n862), .A2(new_n863), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n859), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n438), .A2(new_n842), .A3(new_n857), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT103), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n323), .A2(new_n659), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n324), .A2(new_n327), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n302), .A2(new_n323), .A3(new_n659), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n479), .A2(new_n526), .A3(new_n532), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n572), .A2(new_n577), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(new_n642), .A4(new_n660), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n705), .B1(new_n883), .B2(KEYINPUT31), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n705), .A2(KEYINPUT31), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n880), .B(new_n803), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n875), .B1(new_n876), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n703), .B2(new_n705), .ZN(new_n889));
  OR2_X1    g0689(.A1(KEYINPUT103), .A2(KEYINPUT40), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n889), .A2(new_n803), .A3(new_n880), .A4(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n873), .B(KEYINPUT38), .C1(new_n866), .C2(new_n864), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n435), .A2(new_n842), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n628), .B2(new_n623), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n859), .B1(new_n865), .B2(new_n863), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n866), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n868), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n889), .A2(new_n803), .A3(new_n898), .A4(new_n880), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n888), .A2(new_n891), .B1(KEYINPUT40), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n884), .A2(new_n886), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(new_n440), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n900), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n668), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n892), .A2(new_n897), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT102), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT39), .B1(new_n869), .B2(new_n874), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT102), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n892), .A2(new_n897), .A3(new_n909), .A4(new_n905), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n302), .A2(new_n323), .A3(new_n660), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n880), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n650), .A2(new_n660), .A3(new_n803), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(new_n802), .ZN(new_n917));
  INV_X1    g0717(.A(new_n875), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n917), .A2(new_n918), .B1(new_n624), .B2(new_n657), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n720), .A2(new_n441), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n632), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n904), .B(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n653), .A2(new_n208), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n841), .B1(new_n924), .B2(new_n925), .ZN(G367));
  OAI21_X1  g0726(.A(new_n642), .B1(new_n613), .B2(new_n660), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n647), .A2(new_n659), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(new_n672), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n610), .B1(new_n929), .B2(new_n532), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n660), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n931), .A2(KEYINPUT104), .A3(new_n933), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n936), .B(new_n937), .C1(KEYINPUT42), .C2(new_n930), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n576), .A2(new_n660), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n939), .A2(new_n554), .A3(new_n571), .A4(new_n638), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n709), .B2(new_n939), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n929), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n671), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n938), .A2(new_n945), .A3(new_n942), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n947), .A2(new_n950), .A3(new_n948), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n929), .A2(new_n673), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT105), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT45), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT105), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n954), .B(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n929), .A2(new_n673), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT44), .Z(new_n962));
  NAND3_X1  g0762(.A1(new_n956), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n664), .A2(new_n672), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT106), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n670), .B1(new_n964), .B2(KEYINPUT106), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n671), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n708), .B(new_n720), .C1(new_n963), .C2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n677), .B(KEYINPUT41), .Z(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n723), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n952), .A2(new_n953), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n759), .A2(new_n818), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n382), .B1(new_n213), .B2(new_n752), .C1(new_n766), .C2(new_n732), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n821), .A2(G116), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT46), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT107), .Z(new_n979));
  AOI22_X1  g0779(.A1(new_n774), .A2(G303), .B1(G107), .B2(new_n748), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G311), .A2(new_n756), .B1(new_n765), .B2(G294), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n975), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n973), .B(new_n982), .C1(new_n977), .C2(new_n976), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT109), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n752), .A2(new_n205), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n759), .A2(new_n202), .B1(new_n248), .B2(new_n744), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G150), .C2(new_n774), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n756), .A2(G143), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G68), .A2(new_n748), .B1(new_n765), .B2(G159), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n331), .B1(new_n733), .B2(G137), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n728), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n941), .A2(new_n795), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n784), .B1(new_n791), .B2(new_n339), .C1(new_n244), .C2(new_n787), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n994), .A2(new_n725), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n972), .A2(new_n997), .ZN(G387));
  NAND2_X1  g0798(.A1(new_n721), .A2(new_n967), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n677), .B(KEYINPUT111), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n721), .B2(new_n967), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n723), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n967), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n662), .A2(new_n795), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n403), .A2(new_n202), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n316), .A2(new_n205), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n678), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1008), .A2(G45), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n786), .B1(new_n241), .B2(new_n542), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n791), .A3(new_n278), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n791), .A2(G107), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n784), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n749), .A2(new_n339), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G159), .A2(new_n756), .B1(new_n821), .B2(G77), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n202), .B2(new_n742), .C1(new_n337), .C2(new_n758), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n759), .A2(new_n316), .ZN(new_n1020));
  INV_X1    g0820(.A(G150), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n732), .A2(new_n1021), .ZN(new_n1022));
  OR4_X1    g0822(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n382), .B(new_n1023), .C1(G97), .C2(new_n770), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n774), .A2(G317), .B1(G311), .B2(new_n765), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n756), .A2(G322), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n452), .C2(new_n759), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n501), .B2(new_n744), .C1(new_n749), .C2(new_n818), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT49), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n382), .B1(new_n219), .B2(new_n752), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G326), .B2(new_n733), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1024), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n725), .B(new_n1016), .C1(new_n1033), .C2(new_n729), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT110), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1006), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1035), .B2(new_n1034), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1003), .A2(new_n1005), .A3(new_n1037), .ZN(G393));
  NAND2_X1  g0838(.A1(new_n1000), .A2(new_n963), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(KEYINPUT115), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n963), .A2(new_n671), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n671), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n956), .A2(new_n960), .A3(new_n1042), .A4(new_n962), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1040), .B1(new_n1045), .B2(new_n1000), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1000), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1001), .B1(new_n1047), .B2(KEYINPUT115), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1004), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n252), .A2(new_n786), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n784), .B1(new_n213), .B2(new_n791), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G116), .A2(new_n748), .B1(new_n765), .B2(G303), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n501), .B2(new_n759), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT112), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G107), .B2(new_n770), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n733), .A2(G322), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n742), .A2(new_n762), .B1(new_n766), .B2(new_n755), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n278), .B1(new_n821), .B2(new_n817), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n742), .A2(new_n809), .B1(new_n1021), .B2(new_n755), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT51), .Z(new_n1063));
  NOR2_X1   g0863(.A1(new_n759), .A2(new_n337), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n202), .A2(new_n758), .B1(new_n744), .B2(new_n316), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n733), .A2(G143), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n748), .A2(G77), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1066), .A2(new_n394), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1061), .B1(new_n1069), .B2(new_n816), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT113), .Z(new_n1071));
  OAI221_X1 g0871(.A(new_n725), .B1(new_n1051), .B2(new_n1052), .C1(new_n1071), .C2(new_n729), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT114), .Z(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n795), .B2(new_n944), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1049), .A2(new_n1050), .A3(new_n1074), .ZN(G390));
  INV_X1    g0875(.A(G330), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n901), .A2(new_n440), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n440), .B1(new_n717), .B2(new_n719), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n1078), .A3(new_n631), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n706), .A2(new_n668), .A3(new_n803), .A4(new_n880), .ZN(new_n1080));
  OAI211_X1 g0880(.A(G330), .B(new_n803), .C1(new_n884), .C2(new_n886), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n915), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n660), .B(new_n801), .C1(new_n713), .C2(new_n715), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1083), .A2(new_n802), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n702), .B(new_n660), .C1(new_n695), .C2(new_n699), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n668), .B(new_n803), .C1(new_n884), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n915), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n889), .A2(G330), .A3(new_n803), .A4(new_n880), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1088), .A2(new_n1089), .B1(new_n802), .B2(new_n916), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1079), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n898), .B(new_n912), .C1(new_n1084), .C2(new_n915), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n916), .A2(new_n802), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n913), .B1(new_n1093), .B2(new_n880), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1094), .B2(new_n911), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1089), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1080), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1092), .B(new_n1097), .C1(new_n1094), .C2(new_n911), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1091), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT116), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1001), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n902), .A2(G330), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n921), .A3(new_n632), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1093), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1089), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1093), .A2(new_n880), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n912), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1108), .B1(new_n1112), .B2(new_n1092), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1098), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1091), .A2(new_n1096), .A3(new_n1116), .A4(new_n1098), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1100), .A2(new_n1101), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1004), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n774), .A2(G132), .B1(G128), .B2(new_n756), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT117), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n749), .A2(new_n809), .B1(new_n758), .B2(new_n808), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G125), .B2(new_n733), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n278), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n744), .A2(new_n1021), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1125), .B(new_n1127), .C1(new_n759), .C2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n752), .A2(new_n202), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n774), .A2(G116), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n812), .B1(G77), .B2(new_n748), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G87), .A2(new_n821), .B1(new_n733), .B2(G294), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n331), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(G283), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n759), .A2(new_n213), .B1(new_n1136), .B2(new_n755), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G107), .B2(new_n765), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT118), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1130), .A2(new_n1131), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT119), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n724), .B1(new_n1141), .B2(new_n728), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n403), .B2(new_n829), .C1(new_n911), .C2(new_n782), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1119), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1118), .A2(new_n1145), .ZN(G378));
  OAI22_X1  g0946(.A1(new_n749), .A2(new_n316), .B1(new_n742), .B2(new_n217), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n759), .A2(new_n339), .B1(new_n248), .B2(new_n752), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n205), .B2(new_n744), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G97), .B2(new_n765), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n219), .B2(new_n755), .C1(new_n1136), .C2(new_n732), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1152), .A2(G41), .A3(new_n394), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT58), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n202), .B1(new_n381), .B2(G41), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n759), .A2(new_n808), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G150), .A2(new_n748), .B1(new_n765), .B2(G132), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n756), .A2(G125), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1158), .C1(new_n1159), .C2(new_n742), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1156), .B(new_n1160), .C1(new_n821), .C2(new_n1128), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT59), .ZN(new_n1162));
  AOI21_X1  g0962(.A(G33), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(G41), .B1(new_n733), .B2(G124), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n809), .C2(new_n752), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1155), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n728), .B1(new_n1154), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n724), .B1(new_n202), .B2(new_n828), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n376), .A2(new_n366), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n357), .A2(new_n842), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1172));
  XOR2_X1   g0972(.A(new_n1171), .B(new_n1172), .Z(new_n1173));
  XOR2_X1   g0973(.A(new_n1170), .B(new_n1173), .Z(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1168), .B(new_n1169), .C1(new_n1175), .C2(new_n782), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT120), .Z(new_n1177));
  INV_X1    g0977(.A(new_n920), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n887), .A2(new_n876), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n891), .A2(new_n1179), .A3(new_n918), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n899), .A2(KEYINPUT40), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1175), .B1(new_n1182), .B2(G330), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1076), .B(new_n1174), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1178), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1174), .B1(new_n900), .B2(new_n1076), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(G330), .A3(new_n1175), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n920), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1091), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1185), .B(new_n1188), .C1(new_n1189), .C2(new_n1103), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT57), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1001), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1177), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1186), .A2(new_n1187), .A3(KEYINPUT121), .A4(new_n920), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1101), .A2(new_n1191), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1115), .B2(new_n1079), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1199), .B2(new_n1004), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1193), .A2(new_n1200), .ZN(G375));
  NOR2_X1   g1001(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(new_n723), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n985), .B1(G97), .B2(new_n821), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n501), .B2(new_n755), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n759), .A2(new_n217), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n758), .A2(new_n219), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1205), .A2(new_n1017), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n278), .B1(new_n733), .B2(G303), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n1136), .C2(new_n742), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT122), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n749), .A2(new_n202), .B1(new_n759), .B2(new_n1021), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT123), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n394), .B1(new_n742), .B2(new_n808), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n752), .A2(new_n248), .B1(new_n732), .B2(new_n1159), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n765), .A2(new_n1128), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n821), .A2(G159), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G132), .B2(new_n756), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n728), .B1(new_n1211), .B2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n725), .C1(G68), .C2(new_n829), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n915), .B2(new_n781), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1203), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1202), .A2(new_n1103), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n969), .A3(new_n1091), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(G381));
  NOR3_X1   g1027(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT124), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1046), .A2(new_n1048), .B1(new_n1004), .B2(new_n1045), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1230), .A2(new_n997), .A3(new_n972), .A4(new_n1074), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1189), .B1(KEYINPUT116), .B2(new_n1099), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1117), .A2(new_n1101), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1144), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1193), .A2(new_n1234), .A3(new_n1200), .ZN(new_n1235));
  OR4_X1    g1035(.A1(G381), .A2(new_n1229), .A3(new_n1231), .A4(new_n1235), .ZN(G407));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G343), .C2(new_n1235), .ZN(G409));
  XNOR2_X1  g1037(.A(G393), .B(G396), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G390), .A2(G387), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT126), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1231), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1240), .B1(new_n1239), .B2(new_n1231), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1238), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1238), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G343), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1193), .A2(G378), .A3(new_n1200), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1185), .A2(new_n1004), .A3(new_n1188), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n969), .B1(new_n1189), .B2(new_n1103), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1176), .B(new_n1251), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1234), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1249), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(new_n1225), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT60), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1101), .B1(new_n1225), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1224), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n806), .A3(new_n830), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G384), .B(new_n1224), .C1(new_n1258), .C2(new_n1260), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1250), .A2(new_n1255), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT125), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1249), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1250), .A2(new_n1255), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1249), .A2(G2897), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1264), .B(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1265), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1269), .A2(new_n1270), .A3(new_n1277), .A4(new_n1272), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1247), .B(new_n1267), .C1(new_n1276), .C2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1243), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1241), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1245), .B1(new_n1282), .B2(new_n1238), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1264), .A2(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1256), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1278), .B2(new_n1284), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1277), .B(new_n1274), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(new_n1256), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1283), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1280), .A2(new_n1291), .ZN(G405));
  NAND2_X1  g1092(.A1(G375), .A2(G378), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1293), .B(new_n1235), .C1(new_n1294), .C2(new_n1277), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1264), .A2(KEYINPUT127), .ZN(new_n1296));
  OR2_X1    g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1247), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1283), .A2(new_n1298), .A3(new_n1297), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(G402));
endmodule


