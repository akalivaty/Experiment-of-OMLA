

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791;

  BUF_X1 U370 ( .A(n744), .Z(n347) );
  AND2_X1 U371 ( .A1(n403), .A2(KEYINPUT44), .ZN(n475) );
  XNOR2_X1 U372 ( .A(n510), .B(n369), .ZN(n672) );
  INV_X2 U373 ( .A(G953), .ZN(n776) );
  XNOR2_X2 U374 ( .A(n565), .B(KEYINPUT33), .ZN(n722) );
  XNOR2_X2 U375 ( .A(KEYINPUT72), .B(KEYINPUT19), .ZN(n492) );
  INV_X2 U376 ( .A(G125), .ZN(n460) );
  XNOR2_X2 U377 ( .A(n460), .B(G146), .ZN(n388) );
  XNOR2_X2 U378 ( .A(G113), .B(KEYINPUT67), .ZN(n404) );
  XNOR2_X2 U379 ( .A(n652), .B(KEYINPUT57), .ZN(n653) );
  XNOR2_X2 U380 ( .A(n347), .B(n745), .ZN(n746) );
  XNOR2_X2 U381 ( .A(n353), .B(n738), .ZN(n740) );
  XNOR2_X2 U382 ( .A(n558), .B(KEYINPUT103), .ZN(n352) );
  AND2_X2 U383 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X2 U384 ( .A(n351), .B(G472), .ZN(n559) );
  XNOR2_X1 U385 ( .A(n448), .B(KEYINPUT40), .ZN(n662) );
  NOR2_X2 U386 ( .A1(n673), .A2(n672), .ZN(n637) );
  XNOR2_X2 U387 ( .A(n391), .B(n534), .ZN(n563) );
  NOR2_X2 U388 ( .A1(n350), .A2(n590), .ZN(n565) );
  NOR2_X1 U389 ( .A1(G237), .A2(G953), .ZN(n506) );
  INV_X1 U390 ( .A(n583), .ZN(n590) );
  INV_X1 U391 ( .A(n564), .ZN(n612) );
  AND2_X1 U392 ( .A1(n420), .A2(n449), .ZN(n348) );
  AND2_X1 U393 ( .A1(n414), .A2(n385), .ZN(n413) );
  NAND2_X1 U394 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U395 ( .A1(n662), .A2(n788), .ZN(n440) );
  AND2_X1 U396 ( .A1(n791), .A2(n477), .ZN(n471) );
  NAND2_X1 U397 ( .A1(n638), .A2(n627), .ZN(n448) );
  AND2_X1 U398 ( .A1(n617), .A2(n357), .ZN(n661) );
  OR2_X1 U399 ( .A1(n560), .A2(n394), .ZN(n561) );
  AND2_X1 U400 ( .A1(n623), .A2(n624), .ZN(n625) );
  XNOR2_X1 U401 ( .A(n427), .B(n516), .ZN(n751) );
  NOR2_X1 U402 ( .A1(n423), .A2(G953), .ZN(n422) );
  XNOR2_X1 U403 ( .A(KEYINPUT17), .B(KEYINPUT73), .ZN(n480) );
  XOR2_X1 U404 ( .A(KEYINPUT83), .B(KEYINPUT46), .Z(n628) );
  AND2_X2 U405 ( .A1(n348), .A2(n349), .ZN(n725) );
  NAND2_X1 U406 ( .A1(n455), .A2(n452), .ZN(n349) );
  NAND2_X1 U407 ( .A1(n563), .A2(n701), .ZN(n350) );
  BUF_X1 U408 ( .A(n583), .Z(n394) );
  NOR2_X1 U409 ( .A1(n664), .A2(G902), .ZN(n351) );
  BUF_X1 U410 ( .A(n739), .Z(n353) );
  XNOR2_X1 U411 ( .A(n558), .B(KEYINPUT103), .ZN(n403) );
  XNOR2_X2 U412 ( .A(n567), .B(KEYINPUT35), .ZN(n786) );
  AND2_X1 U413 ( .A1(n580), .A2(n473), .ZN(n472) );
  OR2_X1 U414 ( .A1(n574), .A2(n672), .ZN(n370) );
  INV_X1 U415 ( .A(n370), .ZN(n390) );
  XNOR2_X1 U416 ( .A(n398), .B(G104), .ZN(n502) );
  INV_X1 U417 ( .A(G122), .ZN(n398) );
  XNOR2_X1 U418 ( .A(n401), .B(n400), .ZN(n553) );
  XNOR2_X1 U419 ( .A(n404), .B(n402), .ZN(n401) );
  XNOR2_X1 U420 ( .A(n424), .B(n422), .ZN(n539) );
  XNOR2_X1 U421 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n424) );
  INV_X1 U422 ( .A(G234), .ZN(n423) );
  XNOR2_X1 U423 ( .A(n661), .B(n365), .ZN(n364) );
  INV_X1 U424 ( .A(KEYINPUT78), .ZN(n365) );
  NAND2_X1 U425 ( .A1(n609), .A2(n608), .ZN(n366) );
  NAND2_X1 U426 ( .A1(n607), .A2(n596), .ZN(n608) );
  XNOR2_X1 U427 ( .A(n575), .B(KEYINPUT100), .ZN(n694) );
  NOR2_X1 U428 ( .A1(n627), .A2(n637), .ZN(n575) );
  NOR2_X1 U429 ( .A1(n454), .A2(n453), .ZN(n451) );
  INV_X1 U430 ( .A(n790), .ZN(n450) );
  NOR2_X1 U431 ( .A1(n785), .A2(KEYINPUT82), .ZN(n452) );
  NAND2_X1 U432 ( .A1(n413), .A2(n415), .ZN(n420) );
  AND2_X1 U433 ( .A1(n418), .A2(KEYINPUT82), .ZN(n414) );
  XNOR2_X1 U434 ( .A(n374), .B(KEYINPUT10), .ZN(n538) );
  NAND2_X1 U435 ( .A1(n371), .A2(n372), .ZN(n696) );
  OR2_X1 U436 ( .A1(n751), .A2(G902), .ZN(n518) );
  XNOR2_X1 U437 ( .A(n397), .B(n553), .ZN(n396) );
  XOR2_X1 U438 ( .A(KEYINPUT91), .B(G128), .Z(n536) );
  XNOR2_X1 U439 ( .A(G119), .B(G110), .ZN(n535) );
  XNOR2_X1 U440 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n540) );
  XNOR2_X1 U441 ( .A(n538), .B(n468), .ZN(n773) );
  INV_X1 U442 ( .A(n537), .ZN(n468) );
  XNOR2_X1 U443 ( .A(G116), .B(G122), .ZN(n517) );
  INV_X1 U444 ( .A(KEYINPUT99), .ZN(n511) );
  XNOR2_X1 U445 ( .A(G107), .B(G134), .ZN(n513) );
  XNOR2_X1 U446 ( .A(n442), .B(n441), .ZN(n721) );
  INV_X1 U447 ( .A(KEYINPUT41), .ZN(n441) );
  NAND2_X1 U448 ( .A1(n699), .A2(n632), .ZN(n442) );
  NAND2_X1 U449 ( .A1(n360), .A2(n630), .ZN(n367) );
  NAND2_X1 U450 ( .A1(n426), .A2(n425), .ZN(n607) );
  INV_X1 U451 ( .A(KEYINPUT76), .ZN(n425) );
  NAND2_X1 U452 ( .A1(n694), .A2(KEYINPUT47), .ZN(n426) );
  NAND2_X1 U453 ( .A1(n361), .A2(n367), .ZN(n629) );
  NOR2_X1 U454 ( .A1(n363), .A2(n362), .ZN(n361) );
  NAND2_X1 U455 ( .A1(n366), .A2(n364), .ZN(n363) );
  INV_X1 U456 ( .A(KEYINPUT48), .ZN(n419) );
  XNOR2_X1 U457 ( .A(G902), .B(KEYINPUT88), .ZN(n488) );
  XNOR2_X1 U458 ( .A(G134), .B(G131), .ZN(n525) );
  XOR2_X1 U459 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n541) );
  XNOR2_X1 U460 ( .A(n502), .B(n355), .ZN(n444) );
  XNOR2_X1 U461 ( .A(G143), .B(G140), .ZN(n503) );
  XOR2_X1 U462 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n504) );
  XNOR2_X1 U463 ( .A(G140), .B(G137), .ZN(n537) );
  XNOR2_X1 U464 ( .A(G101), .B(G104), .ZN(n529) );
  INV_X1 U465 ( .A(n729), .ZN(n649) );
  NAND2_X1 U466 ( .A1(G237), .A2(G234), .ZN(n493) );
  NOR2_X1 U467 ( .A1(n451), .A2(n450), .ZN(n449) );
  INV_X1 U468 ( .A(G237), .ZN(n489) );
  AND2_X1 U469 ( .A1(n624), .A2(n696), .ZN(n699) );
  INV_X1 U470 ( .A(KEYINPUT0), .ZN(n446) );
  NAND2_X1 U471 ( .A1(G469), .A2(n408), .ZN(n407) );
  BUF_X1 U472 ( .A(n725), .Z(n775) );
  XNOR2_X1 U473 ( .A(n487), .B(n396), .ZN(n739) );
  NAND2_X1 U474 ( .A1(n434), .A2(n435), .ZN(n432) );
  XNOR2_X1 U475 ( .A(n509), .B(G475), .ZN(n369) );
  INV_X1 U476 ( .A(KEYINPUT124), .ZN(n395) );
  XNOR2_X1 U477 ( .A(n469), .B(n467), .ZN(n756) );
  INV_X1 U478 ( .A(n773), .ZN(n467) );
  XNOR2_X1 U479 ( .A(n544), .B(n545), .ZN(n469) );
  XNOR2_X1 U480 ( .A(n512), .B(n428), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n517), .B(n511), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n657), .B(n656), .ZN(n759) );
  NOR2_X1 U483 ( .A1(n721), .A2(n621), .ZN(n447) );
  NOR2_X1 U484 ( .A1(n711), .A2(n445), .ZN(n573) );
  INV_X1 U485 ( .A(KEYINPUT97), .ZN(n461) );
  INV_X1 U486 ( .A(n367), .ZN(n691) );
  XNOR2_X1 U487 ( .A(n661), .B(n368), .ZN(G45) );
  INV_X1 U488 ( .A(G143), .ZN(n368) );
  INV_X1 U489 ( .A(G110), .ZN(n405) );
  AND2_X1 U490 ( .A1(n433), .A2(n620), .ZN(n354) );
  INV_X1 U491 ( .A(n632), .ZN(n457) );
  XOR2_X1 U492 ( .A(G113), .B(G131), .Z(n355) );
  XOR2_X1 U493 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n356) );
  AND2_X1 U494 ( .A1(n620), .A2(n619), .ZN(n357) );
  INV_X1 U495 ( .A(G902), .ZN(n408) );
  AND2_X1 U496 ( .A1(n466), .A2(n589), .ZN(n358) );
  XNOR2_X1 U497 ( .A(KEYINPUT84), .B(KEYINPUT36), .ZN(n359) );
  INV_X1 U498 ( .A(KEYINPUT101), .ZN(n389) );
  INV_X1 U499 ( .A(KEYINPUT34), .ZN(n435) );
  INV_X1 U500 ( .A(KEYINPUT82), .ZN(n453) );
  INV_X1 U501 ( .A(KEYINPUT44), .ZN(n477) );
  XNOR2_X1 U502 ( .A(n594), .B(n359), .ZN(n360) );
  AND2_X1 U503 ( .A1(n604), .A2(n683), .ZN(n362) );
  NAND2_X1 U504 ( .A1(n390), .A2(n389), .ZN(n371) );
  NAND2_X1 U505 ( .A1(n370), .A2(KEYINPUT101), .ZN(n372) );
  XNOR2_X1 U506 ( .A(n592), .B(n492), .ZN(n373) );
  XNOR2_X1 U507 ( .A(n592), .B(n492), .ZN(n412) );
  XNOR2_X1 U508 ( .A(G146), .B(G125), .ZN(n374) );
  BUF_X1 U509 ( .A(n646), .Z(n764) );
  BUF_X1 U510 ( .A(n352), .Z(n375) );
  BUF_X1 U511 ( .A(n393), .Z(n376) );
  NAND2_X1 U512 ( .A1(n373), .A2(n501), .ZN(n377) );
  NAND2_X1 U513 ( .A1(n412), .A2(n501), .ZN(n458) );
  BUF_X1 U514 ( .A(n396), .Z(n378) );
  BUF_X1 U515 ( .A(n577), .Z(n379) );
  BUF_X1 U516 ( .A(n515), .Z(n380) );
  BUF_X1 U517 ( .A(n722), .Z(n381) );
  NAND2_X2 U518 ( .A1(n386), .A2(n632), .ZN(n592) );
  BUF_X1 U519 ( .A(n553), .Z(n382) );
  INV_X1 U520 ( .A(n705), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n470), .B(n555), .ZN(n664) );
  XNOR2_X1 U522 ( .A(n470), .B(n532), .ZN(n651) );
  AND2_X1 U523 ( .A1(n385), .A2(n418), .ZN(n384) );
  BUF_X1 U524 ( .A(n786), .Z(n383) );
  NOR2_X1 U525 ( .A1(n629), .A2(n419), .ZN(n416) );
  NAND2_X1 U526 ( .A1(n722), .A2(KEYINPUT34), .ZN(n430) );
  INV_X1 U527 ( .A(n386), .ZN(n618) );
  BUF_X1 U528 ( .A(n563), .Z(n630) );
  NAND2_X1 U529 ( .A1(n439), .A2(n419), .ZN(n385) );
  INV_X1 U530 ( .A(n599), .ZN(n708) );
  NAND2_X1 U531 ( .A1(n409), .A2(n406), .ZN(n601) );
  XNOR2_X2 U532 ( .A(n490), .B(n387), .ZN(n386) );
  AND2_X1 U533 ( .A1(n491), .A2(G210), .ZN(n387) );
  NOR2_X2 U534 ( .A1(n599), .A2(n457), .ZN(n456) );
  BUF_X2 U535 ( .A(n559), .Z(n599) );
  XNOR2_X1 U536 ( .A(n456), .B(KEYINPUT30), .ZN(n623) );
  NAND2_X1 U537 ( .A1(n625), .A2(n626), .ZN(n421) );
  NAND2_X2 U538 ( .A1(n409), .A2(n406), .ZN(n391) );
  AND2_X2 U539 ( .A1(n673), .A2(n672), .ZN(n627) );
  XOR2_X1 U540 ( .A(KEYINPUT62), .B(n664), .Z(n665) );
  XNOR2_X1 U541 ( .A(n377), .B(n446), .ZN(n392) );
  XNOR2_X1 U542 ( .A(n458), .B(n446), .ZN(n568) );
  AND2_X2 U543 ( .A1(n650), .A2(n649), .ZN(n393) );
  XNOR2_X2 U544 ( .A(n645), .B(KEYINPUT64), .ZN(n650) );
  XNOR2_X1 U545 ( .A(n559), .B(KEYINPUT6), .ZN(n583) );
  XNOR2_X1 U546 ( .A(n378), .B(n395), .ZN(n763) );
  XNOR2_X1 U547 ( .A(n399), .B(n502), .ZN(n397) );
  XNOR2_X1 U548 ( .A(n527), .B(KEYINPUT16), .ZN(n399) );
  XNOR2_X2 U549 ( .A(G110), .B(G107), .ZN(n527) );
  XNOR2_X1 U550 ( .A(G101), .B(G116), .ZN(n400) );
  XNOR2_X2 U551 ( .A(KEYINPUT3), .B(G119), .ZN(n402) );
  XNOR2_X1 U552 ( .A(n388), .B(n480), .ZN(n483) );
  NOR2_X1 U553 ( .A1(n476), .A2(n352), .ZN(n437) );
  XNOR2_X1 U554 ( .A(n375), .B(n405), .ZN(G12) );
  OR2_X1 U555 ( .A1(n651), .A2(n407), .ZN(n406) );
  NAND2_X1 U556 ( .A1(n533), .A2(G902), .ZN(n410) );
  NAND2_X1 U557 ( .A1(n651), .A2(n533), .ZN(n411) );
  AND2_X1 U558 ( .A1(n373), .A2(n603), .ZN(n683) );
  NAND2_X1 U559 ( .A1(n384), .A2(n415), .ZN(n455) );
  INV_X1 U560 ( .A(n439), .ZN(n417) );
  NAND2_X1 U561 ( .A1(n629), .A2(n419), .ZN(n418) );
  XNOR2_X1 U562 ( .A(n526), .B(n486), .ZN(n487) );
  XNOR2_X2 U563 ( .A(n421), .B(KEYINPUT39), .ZN(n638) );
  INV_X1 U564 ( .A(n785), .ZN(n454) );
  NAND2_X1 U565 ( .A1(n474), .A2(n472), .ZN(n436) );
  XNOR2_X1 U566 ( .A(n436), .B(KEYINPUT45), .ZN(n646) );
  NOR2_X2 U567 ( .A1(n431), .A2(n429), .ZN(n567) );
  NAND2_X1 U568 ( .A1(n430), .A2(n354), .ZN(n429) );
  NOR2_X1 U569 ( .A1(n722), .A2(n432), .ZN(n431) );
  NAND2_X1 U570 ( .A1(n445), .A2(KEYINPUT34), .ZN(n433) );
  INV_X1 U571 ( .A(n445), .ZN(n434) );
  INV_X1 U572 ( .A(n392), .ZN(n445) );
  NOR2_X1 U573 ( .A1(n475), .A2(n437), .ZN(n474) );
  NAND2_X1 U574 ( .A1(n786), .A2(n471), .ZN(n476) );
  XNOR2_X1 U575 ( .A(n438), .B(n743), .ZN(G51) );
  NAND2_X1 U576 ( .A1(n742), .A2(n759), .ZN(n438) );
  AND2_X2 U577 ( .A1(n650), .A2(n649), .ZN(n755) );
  XNOR2_X2 U578 ( .A(n440), .B(n628), .ZN(n439) );
  XNOR2_X1 U579 ( .A(n447), .B(n622), .ZN(n788) );
  XNOR2_X1 U580 ( .A(n508), .B(n443), .ZN(n744) );
  XNOR2_X1 U581 ( .A(n505), .B(n444), .ZN(n443) );
  NOR2_X1 U582 ( .A1(n744), .A2(G902), .ZN(n510) );
  XNOR2_X2 U583 ( .A(n459), .B(KEYINPUT32), .ZN(n791) );
  OR2_X1 U584 ( .A1(n562), .A2(n561), .ZN(n459) );
  NAND2_X1 U585 ( .A1(n674), .A2(n688), .ZN(n576) );
  XNOR2_X2 U586 ( .A(n462), .B(n461), .ZN(n674) );
  NAND2_X1 U587 ( .A1(n464), .A2(n463), .ZN(n462) );
  INV_X1 U588 ( .A(n708), .ZN(n463) );
  XNOR2_X1 U589 ( .A(n571), .B(n465), .ZN(n464) );
  INV_X1 U590 ( .A(KEYINPUT96), .ZN(n465) );
  NOR2_X1 U591 ( .A1(n598), .A2(n599), .ZN(n600) );
  NAND2_X1 U592 ( .A1(n564), .A2(n358), .ZN(n598) );
  XNOR2_X2 U593 ( .A(n774), .B(G146), .ZN(n470) );
  NAND2_X1 U594 ( .A1(n786), .A2(n791), .ZN(n478) );
  NAND2_X1 U595 ( .A1(n478), .A2(KEYINPUT44), .ZN(n473) );
  XNOR2_X1 U596 ( .A(n758), .B(n757), .ZN(n760) );
  NAND2_X1 U597 ( .A1(n658), .A2(n759), .ZN(n660) );
  XNOR2_X1 U598 ( .A(n654), .B(n653), .ZN(n658) );
  XNOR2_X2 U599 ( .A(n549), .B(n548), .ZN(n564) );
  NAND2_X1 U600 ( .A1(n393), .A2(G217), .ZN(n758) );
  NOR2_X2 U601 ( .A1(n562), .A2(n630), .ZN(n577) );
  XNOR2_X1 U602 ( .A(n538), .B(n507), .ZN(n508) );
  AND2_X1 U603 ( .A1(G217), .A2(n546), .ZN(n479) );
  XNOR2_X1 U604 ( .A(n694), .B(KEYINPUT77), .ZN(n595) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(n544) );
  INV_X1 U606 ( .A(KEYINPUT71), .ZN(n615) );
  XNOR2_X1 U607 ( .A(n747), .B(n746), .ZN(n748) );
  INV_X1 U608 ( .A(KEYINPUT118), .ZN(n659) );
  NAND2_X1 U609 ( .A1(n776), .A2(G224), .ZN(n481) );
  XNOR2_X1 U610 ( .A(n481), .B(KEYINPUT18), .ZN(n482) );
  XNOR2_X1 U611 ( .A(n483), .B(n482), .ZN(n486) );
  XNOR2_X2 U612 ( .A(G143), .B(KEYINPUT74), .ZN(n485) );
  INV_X1 U613 ( .A(G128), .ZN(n484) );
  XNOR2_X2 U614 ( .A(n485), .B(n484), .ZN(n515) );
  XNOR2_X2 U615 ( .A(n515), .B(KEYINPUT4), .ZN(n526) );
  XNOR2_X1 U616 ( .A(n488), .B(KEYINPUT15), .ZN(n581) );
  NAND2_X1 U617 ( .A1(n739), .A2(n581), .ZN(n490) );
  NAND2_X1 U618 ( .A1(n408), .A2(n489), .ZN(n491) );
  NAND2_X1 U619 ( .A1(n491), .A2(G214), .ZN(n632) );
  XOR2_X1 U620 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n494) );
  XNOR2_X1 U621 ( .A(n494), .B(n493), .ZN(n497) );
  NAND2_X1 U622 ( .A1(G952), .A2(n497), .ZN(n719) );
  NOR2_X1 U623 ( .A1(G953), .A2(n719), .ZN(n495) );
  XNOR2_X1 U624 ( .A(n495), .B(KEYINPUT89), .ZN(n587) );
  NOR2_X1 U625 ( .A1(G898), .A2(n776), .ZN(n496) );
  XOR2_X1 U626 ( .A(KEYINPUT90), .B(n496), .Z(n762) );
  INV_X1 U627 ( .A(n762), .ZN(n499) );
  NAND2_X1 U628 ( .A1(G902), .A2(n497), .ZN(n584) );
  INV_X1 U629 ( .A(n584), .ZN(n498) );
  NAND2_X1 U630 ( .A1(n499), .A2(n498), .ZN(n500) );
  NAND2_X1 U631 ( .A1(n587), .A2(n500), .ZN(n501) );
  XNOR2_X1 U632 ( .A(n503), .B(n504), .ZN(n505) );
  XNOR2_X1 U633 ( .A(n506), .B(KEYINPUT70), .ZN(n550) );
  NAND2_X1 U634 ( .A1(G214), .A2(n550), .ZN(n507) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n509) );
  NAND2_X1 U636 ( .A1(G217), .A2(n539), .ZN(n512) );
  XNOR2_X1 U637 ( .A(n356), .B(n513), .ZN(n514) );
  XNOR2_X1 U638 ( .A(n380), .B(n514), .ZN(n516) );
  XNOR2_X1 U639 ( .A(n518), .B(G478), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n581), .A2(G234), .ZN(n519) );
  XNOR2_X1 U641 ( .A(n519), .B(KEYINPUT20), .ZN(n520) );
  XNOR2_X1 U642 ( .A(KEYINPUT94), .B(n520), .ZN(n546) );
  AND2_X1 U643 ( .A1(n546), .A2(G221), .ZN(n522) );
  INV_X1 U644 ( .A(KEYINPUT21), .ZN(n521) );
  XNOR2_X1 U645 ( .A(n522), .B(n521), .ZN(n705) );
  AND2_X1 U646 ( .A1(n696), .A2(n466), .ZN(n523) );
  NAND2_X1 U647 ( .A1(n568), .A2(n523), .ZN(n524) );
  XNOR2_X1 U648 ( .A(n524), .B(KEYINPUT22), .ZN(n562) );
  XNOR2_X2 U649 ( .A(n526), .B(n525), .ZN(n774) );
  XNOR2_X1 U650 ( .A(n527), .B(n537), .ZN(n531) );
  NAND2_X1 U651 ( .A1(n776), .A2(G227), .ZN(n528) );
  XNOR2_X1 U652 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U653 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U654 ( .A(G469), .ZN(n533) );
  XNOR2_X1 U655 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U656 ( .A(n577), .B(KEYINPUT102), .ZN(n557) );
  XNOR2_X1 U657 ( .A(n536), .B(n535), .ZN(n545) );
  NAND2_X1 U658 ( .A1(G221), .A2(n539), .ZN(n543) );
  XNOR2_X1 U659 ( .A(n541), .B(n540), .ZN(n542) );
  NOR2_X1 U660 ( .A1(n756), .A2(G902), .ZN(n549) );
  XOR2_X1 U661 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n547) );
  XNOR2_X1 U662 ( .A(n547), .B(n479), .ZN(n548) );
  NAND2_X1 U663 ( .A1(G210), .A2(n550), .ZN(n552) );
  XNOR2_X1 U664 ( .A(G137), .B(KEYINPUT5), .ZN(n551) );
  XNOR2_X1 U665 ( .A(n552), .B(n551), .ZN(n554) );
  XNOR2_X1 U666 ( .A(n554), .B(n382), .ZN(n555) );
  NOR2_X1 U667 ( .A1(n612), .A2(n708), .ZN(n556) );
  NAND2_X1 U668 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U669 ( .A1(n563), .A2(n564), .ZN(n560) );
  NOR2_X1 U670 ( .A1(n564), .A2(n705), .ZN(n701) );
  NAND2_X1 U671 ( .A1(n672), .A2(n574), .ZN(n566) );
  XOR2_X1 U672 ( .A(n566), .B(KEYINPUT104), .Z(n620) );
  AND2_X1 U673 ( .A1(n392), .A2(n466), .ZN(n570) );
  NOR2_X1 U674 ( .A1(n564), .A2(n601), .ZN(n569) );
  NAND2_X1 U675 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U676 ( .A1(n701), .A2(n563), .ZN(n572) );
  OR2_X1 U677 ( .A1(n572), .A2(n463), .ZN(n711) );
  XNOR2_X1 U678 ( .A(n573), .B(KEYINPUT31), .ZN(n688) );
  INV_X1 U679 ( .A(n574), .ZN(n673) );
  NAND2_X1 U680 ( .A1(n576), .A2(n595), .ZN(n579) );
  NOR2_X1 U681 ( .A1(n394), .A2(n564), .ZN(n578) );
  NAND2_X1 U682 ( .A1(n379), .A2(n578), .ZN(n670) );
  AND2_X1 U683 ( .A1(n579), .A2(n670), .ZN(n580) );
  INV_X1 U684 ( .A(n581), .ZN(n642) );
  NAND2_X1 U685 ( .A1(n646), .A2(n642), .ZN(n582) );
  XNOR2_X1 U686 ( .A(n582), .B(KEYINPUT81), .ZN(n640) );
  NOR2_X1 U687 ( .A1(G900), .A2(n584), .ZN(n585) );
  NAND2_X1 U688 ( .A1(G953), .A2(n585), .ZN(n586) );
  XOR2_X1 U689 ( .A(n586), .B(KEYINPUT105), .Z(n588) );
  AND2_X1 U690 ( .A1(n588), .A2(n587), .ZN(n610) );
  INV_X1 U691 ( .A(n610), .ZN(n589) );
  NOR2_X1 U692 ( .A1(n590), .A2(n598), .ZN(n591) );
  NAND2_X1 U693 ( .A1(n591), .A2(n627), .ZN(n631) );
  XNOR2_X1 U694 ( .A(KEYINPUT108), .B(n631), .ZN(n593) );
  NOR2_X1 U695 ( .A1(n593), .A2(n592), .ZN(n594) );
  INV_X1 U696 ( .A(n630), .ZN(n703) );
  INV_X1 U697 ( .A(KEYINPUT47), .ZN(n596) );
  AND2_X1 U698 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U699 ( .A(KEYINPUT68), .B(n597), .ZN(n604) );
  XNOR2_X1 U700 ( .A(KEYINPUT28), .B(n600), .ZN(n602) );
  INV_X1 U701 ( .A(n601), .ZN(n613) );
  NAND2_X1 U702 ( .A1(n602), .A2(n613), .ZN(n621) );
  INV_X1 U703 ( .A(n621), .ZN(n603) );
  NAND2_X1 U704 ( .A1(n694), .A2(KEYINPUT76), .ZN(n605) );
  AND2_X1 U705 ( .A1(n605), .A2(n607), .ZN(n606) );
  NAND2_X1 U706 ( .A1(n683), .A2(n606), .ZN(n609) );
  NOR2_X1 U707 ( .A1(n705), .A2(n610), .ZN(n611) );
  AND2_X1 U708 ( .A1(n612), .A2(n611), .ZN(n614) );
  AND2_X1 U709 ( .A1(n614), .A2(n613), .ZN(n616) );
  XNOR2_X1 U710 ( .A(n616), .B(n615), .ZN(n626) );
  AND2_X1 U711 ( .A1(n623), .A2(n626), .ZN(n617) );
  INV_X1 U712 ( .A(n618), .ZN(n619) );
  XNOR2_X1 U713 ( .A(n618), .B(KEYINPUT38), .ZN(n624) );
  INV_X1 U714 ( .A(n624), .ZN(n693) );
  XNOR2_X1 U715 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n622) );
  INV_X1 U716 ( .A(n627), .ZN(n685) );
  NOR2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U719 ( .A(n634), .B(KEYINPUT43), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n635), .A2(n618), .ZN(n636) );
  XOR2_X1 U721 ( .A(KEYINPUT106), .B(n636), .Z(n785) );
  NAND2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U723 ( .A(KEYINPUT109), .B(n639), .Z(n790) );
  NAND2_X1 U724 ( .A1(n640), .A2(n725), .ZN(n641) );
  XNOR2_X1 U725 ( .A(n641), .B(KEYINPUT80), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n642), .A2(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n725), .A2(KEYINPUT2), .ZN(n648) );
  INV_X1 U729 ( .A(n764), .ZN(n647) );
  NOR2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n729) );
  NAND2_X1 U731 ( .A1(n755), .A2(G469), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n651), .B(KEYINPUT58), .ZN(n652) );
  INV_X1 U733 ( .A(G952), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n655), .A2(G953), .ZN(n657) );
  INV_X1 U735 ( .A(KEYINPUT87), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n660), .B(n659), .ZN(G54) );
  BUF_X1 U737 ( .A(n662), .Z(n663) );
  XNOR2_X1 U738 ( .A(n663), .B(G131), .ZN(G33) );
  NAND2_X1 U739 ( .A1(n393), .A2(G472), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n667), .A2(n759), .ZN(n669) );
  XOR2_X1 U742 ( .A(KEYINPUT85), .B(KEYINPUT63), .Z(n668) );
  XNOR2_X1 U743 ( .A(n669), .B(n668), .ZN(G57) );
  XNOR2_X1 U744 ( .A(G101), .B(n670), .ZN(G3) );
  NOR2_X1 U745 ( .A1(n685), .A2(n674), .ZN(n671) );
  XOR2_X1 U746 ( .A(G104), .B(n671), .Z(G6) );
  OR2_X1 U747 ( .A1(n673), .A2(n672), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n689), .A2(n674), .ZN(n679) );
  XOR2_X1 U749 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n676) );
  XNOR2_X1 U750 ( .A(G107), .B(KEYINPUT110), .ZN(n675) );
  XNOR2_X1 U751 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U752 ( .A(KEYINPUT26), .B(n677), .ZN(n678) );
  XNOR2_X1 U753 ( .A(n679), .B(n678), .ZN(G9) );
  XOR2_X1 U754 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n681) );
  NAND2_X1 U755 ( .A1(n683), .A2(n637), .ZN(n680) );
  XNOR2_X1 U756 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U757 ( .A(G128), .B(n682), .ZN(G30) );
  NAND2_X1 U758 ( .A1(n683), .A2(n627), .ZN(n684) );
  XNOR2_X1 U759 ( .A(n684), .B(G146), .ZN(G48) );
  NOR2_X1 U760 ( .A1(n685), .A2(n688), .ZN(n687) );
  XNOR2_X1 U761 ( .A(G113), .B(KEYINPUT113), .ZN(n686) );
  XNOR2_X1 U762 ( .A(n687), .B(n686), .ZN(G15) );
  NOR2_X1 U763 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U764 ( .A(G116), .B(n690), .Z(G18) );
  XNOR2_X1 U765 ( .A(G125), .B(n691), .ZN(n692) );
  XNOR2_X1 U766 ( .A(n692), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U767 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U768 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U769 ( .A1(n697), .A2(n457), .ZN(n698) );
  NOR2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U771 ( .A1(n381), .A2(n700), .ZN(n716) );
  INV_X1 U772 ( .A(n701), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U774 ( .A(n704), .B(KEYINPUT50), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n564), .A2(n705), .ZN(n706) );
  XNOR2_X1 U776 ( .A(KEYINPUT49), .B(n706), .ZN(n707) );
  NOR2_X1 U777 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U778 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U780 ( .A(KEYINPUT51), .B(n713), .ZN(n714) );
  NOR2_X1 U781 ( .A1(n721), .A2(n714), .ZN(n715) );
  NOR2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U783 ( .A(n717), .B(KEYINPUT52), .ZN(n718) );
  NOR2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U785 ( .A(n720), .B(KEYINPUT115), .ZN(n724) );
  OR2_X1 U786 ( .A1(n381), .A2(n721), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n734) );
  XOR2_X1 U788 ( .A(KEYINPUT2), .B(KEYINPUT75), .Z(n727) );
  NOR2_X1 U789 ( .A1(n775), .A2(n727), .ZN(n726) );
  XNOR2_X1 U790 ( .A(n726), .B(KEYINPUT79), .ZN(n731) );
  NOR2_X1 U791 ( .A1(n764), .A2(n727), .ZN(n728) );
  NOR2_X1 U792 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U793 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U794 ( .A1(n732), .A2(n776), .ZN(n733) );
  NOR2_X1 U795 ( .A1(n734), .A2(n733), .ZN(n736) );
  XNOR2_X1 U796 ( .A(KEYINPUT53), .B(KEYINPUT116), .ZN(n735) );
  XNOR2_X1 U797 ( .A(n736), .B(n735), .ZN(G75) );
  XNOR2_X1 U798 ( .A(KEYINPUT117), .B(KEYINPUT56), .ZN(n743) );
  NAND2_X1 U799 ( .A1(n755), .A2(G210), .ZN(n741) );
  XOR2_X1 U800 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n737) );
  XNOR2_X1 U801 ( .A(n737), .B(KEYINPUT86), .ZN(n738) );
  XNOR2_X1 U802 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U803 ( .A1(n755), .A2(G475), .ZN(n747) );
  XOR2_X1 U804 ( .A(KEYINPUT59), .B(KEYINPUT119), .Z(n745) );
  NAND2_X1 U805 ( .A1(n748), .A2(n759), .ZN(n750) );
  XOR2_X1 U806 ( .A(KEYINPUT60), .B(KEYINPUT120), .Z(n749) );
  XNOR2_X1 U807 ( .A(n750), .B(n749), .ZN(G60) );
  INV_X1 U808 ( .A(n759), .ZN(n754) );
  NAND2_X1 U809 ( .A1(n376), .A2(G478), .ZN(n752) );
  XNOR2_X1 U810 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U811 ( .A1(n754), .A2(n753), .ZN(G63) );
  INV_X1 U812 ( .A(n756), .ZN(n757) );
  NAND2_X1 U813 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U814 ( .A(n761), .B(KEYINPUT121), .ZN(G66) );
  NAND2_X1 U815 ( .A1(n763), .A2(n762), .ZN(n772) );
  NAND2_X1 U816 ( .A1(n764), .A2(n776), .ZN(n770) );
  NAND2_X1 U817 ( .A1(G224), .A2(G953), .ZN(n765) );
  XNOR2_X1 U818 ( .A(n765), .B(KEYINPUT122), .ZN(n766) );
  XNOR2_X1 U819 ( .A(KEYINPUT61), .B(n766), .ZN(n767) );
  NAND2_X1 U820 ( .A1(n767), .A2(G898), .ZN(n768) );
  XOR2_X1 U821 ( .A(KEYINPUT123), .B(n768), .Z(n769) );
  NAND2_X1 U822 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U823 ( .A(n772), .B(n771), .Z(G69) );
  XNOR2_X1 U824 ( .A(n774), .B(n773), .ZN(n778) );
  XNOR2_X1 U825 ( .A(n775), .B(n778), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n777), .A2(n776), .ZN(n783) );
  XOR2_X1 U827 ( .A(G227), .B(n778), .Z(n779) );
  NAND2_X1 U828 ( .A1(n779), .A2(G900), .ZN(n780) );
  XOR2_X1 U829 ( .A(KEYINPUT125), .B(n780), .Z(n781) );
  NAND2_X1 U830 ( .A1(G953), .A2(n781), .ZN(n782) );
  NAND2_X1 U831 ( .A1(n783), .A2(n782), .ZN(G72) );
  XOR2_X1 U832 ( .A(G140), .B(KEYINPUT114), .Z(n784) );
  XNOR2_X1 U833 ( .A(n785), .B(n784), .ZN(G42) );
  INV_X1 U834 ( .A(n383), .ZN(n787) );
  XOR2_X1 U835 ( .A(G122), .B(n787), .Z(G24) );
  XNOR2_X1 U836 ( .A(G137), .B(n788), .ZN(n789) );
  XNOR2_X1 U837 ( .A(n789), .B(KEYINPUT126), .ZN(G39) );
  XNOR2_X1 U838 ( .A(G134), .B(n790), .ZN(G36) );
  XNOR2_X1 U839 ( .A(n791), .B(G119), .ZN(G21) );
endmodule

