

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591;

  INV_X1 U321 ( .A(KEYINPUT27), .ZN(n420) );
  INV_X1 U322 ( .A(KEYINPUT10), .ZN(n439) );
  INV_X1 U323 ( .A(KEYINPUT95), .ZN(n425) );
  NOR2_X1 U324 ( .A1(n424), .A2(n423), .ZN(n426) );
  XNOR2_X1 U325 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U326 ( .A(n450), .B(n449), .ZN(n548) );
  XNOR2_X1 U327 ( .A(n448), .B(n447), .ZN(n449) );
  INV_X1 U328 ( .A(n434), .ZN(n414) );
  XNOR2_X1 U329 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U330 ( .A(n322), .B(n321), .Z(n289) );
  XOR2_X1 U331 ( .A(n400), .B(KEYINPUT21), .Z(n290) );
  AND2_X1 U332 ( .A1(n453), .A2(n452), .ZN(n291) );
  AND2_X1 U333 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n330), .B(n329), .ZN(n459) );
  INV_X1 U335 ( .A(KEYINPUT64), .ZN(n470) );
  XNOR2_X1 U336 ( .A(n443), .B(n292), .ZN(n389) );
  XNOR2_X1 U337 ( .A(n470), .B(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U338 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U339 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U340 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U341 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U342 ( .A(n398), .B(n397), .ZN(n402) );
  NOR2_X1 U343 ( .A1(n432), .A2(n431), .ZN(n486) );
  XNOR2_X1 U344 ( .A(KEYINPUT94), .B(n404), .ZN(n575) );
  XNOR2_X1 U345 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U346 ( .A(n479), .B(KEYINPUT121), .ZN(n562) );
  XNOR2_X1 U347 ( .A(n417), .B(n416), .ZN(n418) );
  BUF_X1 U348 ( .A(n562), .Z(n572) );
  NOR2_X1 U349 ( .A1(n520), .A2(n519), .ZN(n528) );
  XNOR2_X1 U350 ( .A(n480), .B(G176GAT), .ZN(n481) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n457) );
  XNOR2_X1 U352 ( .A(n482), .B(n481), .ZN(G1349GAT) );
  XNOR2_X1 U353 ( .A(n458), .B(n457), .ZN(G1330GAT) );
  XOR2_X1 U354 ( .A(KEYINPUT29), .B(G113GAT), .Z(n294) );
  XNOR2_X1 U355 ( .A(G141GAT), .B(G197GAT), .ZN(n293) );
  XNOR2_X1 U356 ( .A(n294), .B(n293), .ZN(n307) );
  XOR2_X1 U357 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n296) );
  NAND2_X1 U358 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U359 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U360 ( .A(n297), .B(KEYINPUT30), .Z(n302) );
  XOR2_X1 U361 ( .A(G29GAT), .B(G43GAT), .Z(n299) );
  XNOR2_X1 U362 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n438) );
  XNOR2_X1 U364 ( .A(G22GAT), .B(G15GAT), .ZN(n300) );
  XNOR2_X1 U365 ( .A(n300), .B(G1GAT), .ZN(n344) );
  XNOR2_X1 U366 ( .A(n438), .B(n344), .ZN(n301) );
  XNOR2_X1 U367 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U368 ( .A(G169GAT), .B(G8GAT), .Z(n413) );
  XOR2_X1 U369 ( .A(n303), .B(n413), .Z(n305) );
  XNOR2_X1 U370 ( .A(G36GAT), .B(G50GAT), .ZN(n304) );
  XNOR2_X1 U371 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U372 ( .A(n307), .B(n306), .Z(n578) );
  INV_X1 U373 ( .A(n578), .ZN(n563) );
  XNOR2_X1 U374 ( .A(G99GAT), .B(G85GAT), .ZN(n313) );
  INV_X1 U375 ( .A(KEYINPUT70), .ZN(n308) );
  NAND2_X1 U376 ( .A1(n308), .A2(G92GAT), .ZN(n311) );
  INV_X1 U377 ( .A(G92GAT), .ZN(n309) );
  NAND2_X1 U378 ( .A1(n309), .A2(KEYINPUT70), .ZN(n310) );
  NAND2_X1 U379 ( .A1(n311), .A2(n310), .ZN(n312) );
  XNOR2_X1 U380 ( .A(n313), .B(n312), .ZN(n435) );
  INV_X1 U381 ( .A(n435), .ZN(n314) );
  NAND2_X1 U382 ( .A1(n314), .A2(KEYINPUT33), .ZN(n317) );
  INV_X1 U383 ( .A(KEYINPUT33), .ZN(n315) );
  NAND2_X1 U384 ( .A1(n435), .A2(n315), .ZN(n316) );
  NAND2_X1 U385 ( .A1(n317), .A2(n316), .ZN(n319) );
  NAND2_X1 U386 ( .A1(G230GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U387 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U388 ( .A(n320), .B(KEYINPUT71), .Z(n322) );
  XOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT13), .Z(n340) );
  XNOR2_X1 U390 ( .A(G204GAT), .B(n340), .ZN(n321) );
  XOR2_X1 U391 ( .A(G176GAT), .B(G64GAT), .Z(n408) );
  XNOR2_X1 U392 ( .A(n289), .B(n408), .ZN(n330) );
  XOR2_X1 U393 ( .A(G120GAT), .B(G71GAT), .Z(n380) );
  XOR2_X1 U394 ( .A(G78GAT), .B(G148GAT), .Z(n324) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(KEYINPUT69), .ZN(n323) );
  XNOR2_X1 U396 ( .A(n324), .B(n323), .ZN(n390) );
  XNOR2_X1 U397 ( .A(n380), .B(n390), .ZN(n328) );
  XOR2_X1 U398 ( .A(KEYINPUT68), .B(KEYINPUT31), .Z(n326) );
  XNOR2_X1 U399 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n325) );
  XNOR2_X1 U400 ( .A(n326), .B(n325), .ZN(n327) );
  NAND2_X1 U401 ( .A1(n563), .A2(n459), .ZN(n488) );
  XOR2_X1 U402 ( .A(G64GAT), .B(G183GAT), .Z(n332) );
  XNOR2_X1 U403 ( .A(G8GAT), .B(G127GAT), .ZN(n331) );
  XNOR2_X1 U404 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U405 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n334) );
  XNOR2_X1 U406 ( .A(KEYINPUT74), .B(KEYINPUT12), .ZN(n333) );
  XNOR2_X1 U407 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U408 ( .A(n336), .B(n335), .ZN(n348) );
  XOR2_X1 U409 ( .A(G78GAT), .B(G155GAT), .Z(n338) );
  XNOR2_X1 U410 ( .A(G71GAT), .B(G211GAT), .ZN(n337) );
  XNOR2_X1 U411 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U412 ( .A(n340), .B(n339), .Z(n342) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U414 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U415 ( .A(n343), .B(KEYINPUT75), .Z(n346) );
  XNOR2_X1 U416 ( .A(n344), .B(KEYINPUT15), .ZN(n345) );
  XNOR2_X1 U417 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U418 ( .A(n348), .B(n347), .ZN(n566) );
  XOR2_X1 U419 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n350) );
  XNOR2_X1 U420 ( .A(KEYINPUT88), .B(KEYINPUT5), .ZN(n349) );
  XNOR2_X1 U421 ( .A(n350), .B(n349), .ZN(n369) );
  XOR2_X1 U422 ( .A(G85GAT), .B(G148GAT), .Z(n352) );
  XNOR2_X1 U423 ( .A(G29GAT), .B(G162GAT), .ZN(n351) );
  XNOR2_X1 U424 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U425 ( .A(KEYINPUT1), .B(G57GAT), .Z(n354) );
  XNOR2_X1 U426 ( .A(G1GAT), .B(G120GAT), .ZN(n353) );
  XNOR2_X1 U427 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U428 ( .A(n356), .B(n355), .Z(n367) );
  XNOR2_X1 U429 ( .A(G127GAT), .B(KEYINPUT79), .ZN(n357) );
  XNOR2_X1 U430 ( .A(n357), .B(KEYINPUT0), .ZN(n358) );
  XOR2_X1 U431 ( .A(n358), .B(KEYINPUT78), .Z(n360) );
  XNOR2_X1 U432 ( .A(G113GAT), .B(G134GAT), .ZN(n359) );
  XNOR2_X1 U433 ( .A(n360), .B(n359), .ZN(n388) );
  XOR2_X1 U434 ( .A(G155GAT), .B(KEYINPUT2), .Z(n362) );
  XNOR2_X1 U435 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n361) );
  XNOR2_X1 U436 ( .A(n362), .B(n361), .ZN(n392) );
  XOR2_X1 U437 ( .A(n392), .B(KEYINPUT4), .Z(n364) );
  NAND2_X1 U438 ( .A1(G225GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U439 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U440 ( .A(n388), .B(n365), .ZN(n366) );
  XNOR2_X1 U441 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U442 ( .A(n369), .B(n368), .Z(n521) );
  XOR2_X1 U443 ( .A(KEYINPUT82), .B(G190GAT), .Z(n371) );
  XNOR2_X1 U444 ( .A(G43GAT), .B(G99GAT), .ZN(n370) );
  XNOR2_X1 U445 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U446 ( .A(G176GAT), .B(KEYINPUT83), .Z(n373) );
  XNOR2_X1 U447 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n372) );
  XNOR2_X1 U448 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U449 ( .A(n375), .B(n374), .Z(n386) );
  XOR2_X1 U450 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n377) );
  XNOR2_X1 U451 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n376) );
  XNOR2_X1 U452 ( .A(n377), .B(n376), .ZN(n384) );
  XOR2_X1 U453 ( .A(G183GAT), .B(KEYINPUT17), .Z(n379) );
  XNOR2_X1 U454 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n378) );
  XNOR2_X1 U455 ( .A(n379), .B(n378), .ZN(n412) );
  XOR2_X1 U456 ( .A(n380), .B(n412), .Z(n382) );
  NAND2_X1 U457 ( .A1(G227GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U458 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U459 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U460 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U461 ( .A(n388), .B(n387), .ZN(n536) );
  XOR2_X1 U462 ( .A(G50GAT), .B(G162GAT), .Z(n443) );
  XOR2_X1 U463 ( .A(n391), .B(KEYINPUT86), .Z(n398) );
  XNOR2_X1 U464 ( .A(n392), .B(KEYINPUT23), .ZN(n396) );
  XOR2_X1 U465 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n394) );
  XNOR2_X1 U466 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U468 ( .A(G211GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n399), .B(KEYINPUT85), .ZN(n400) );
  XNOR2_X1 U470 ( .A(G197GAT), .B(G204GAT), .ZN(n401) );
  XOR2_X1 U471 ( .A(n290), .B(n401), .Z(n409) );
  XNOR2_X1 U472 ( .A(n402), .B(n409), .ZN(n476) );
  NOR2_X1 U473 ( .A1(n536), .A2(n476), .ZN(n403) );
  XOR2_X1 U474 ( .A(KEYINPUT26), .B(n403), .Z(n404) );
  XOR2_X1 U475 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n406) );
  NAND2_X1 U476 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U478 ( .A(KEYINPUT93), .B(n407), .Z(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT90), .B(n408), .Z(n411) );
  XOR2_X1 U480 ( .A(n409), .B(G92GAT), .Z(n410) );
  XNOR2_X1 U481 ( .A(n411), .B(n410), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U483 ( .A(G36GAT), .B(G190GAT), .Z(n434) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n525) );
  XNOR2_X1 U485 ( .A(n525), .B(n420), .ZN(n428) );
  NOR2_X1 U486 ( .A1(n575), .A2(n428), .ZN(n424) );
  NAND2_X1 U487 ( .A1(n536), .A2(n525), .ZN(n421) );
  NAND2_X1 U488 ( .A1(n476), .A2(n421), .ZN(n422) );
  XNOR2_X1 U489 ( .A(n422), .B(KEYINPUT25), .ZN(n423) );
  NOR2_X1 U490 ( .A1(n521), .A2(n427), .ZN(n432) );
  INV_X1 U491 ( .A(n521), .ZN(n429) );
  NOR2_X1 U492 ( .A1(n429), .A2(n428), .ZN(n533) );
  XNOR2_X1 U493 ( .A(KEYINPUT28), .B(n476), .ZN(n497) );
  NAND2_X1 U494 ( .A1(n533), .A2(n497), .ZN(n430) );
  NOR2_X1 U495 ( .A1(n430), .A2(n536), .ZN(n431) );
  NOR2_X1 U496 ( .A1(n566), .A2(n486), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n433), .B(KEYINPUT102), .ZN(n453) );
  XOR2_X1 U498 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U499 ( .A1(G232GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n438), .B(KEYINPUT11), .ZN(n440) );
  XOR2_X1 U502 ( .A(n444), .B(n443), .Z(n450) );
  XOR2_X1 U503 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n446) );
  XNOR2_X1 U504 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n445) );
  XOR2_X1 U505 ( .A(n446), .B(n445), .Z(n448) );
  XNOR2_X1 U506 ( .A(G134GAT), .B(G218GAT), .ZN(n447) );
  XOR2_X1 U507 ( .A(KEYINPUT36), .B(KEYINPUT101), .Z(n451) );
  XNOR2_X1 U508 ( .A(n548), .B(n451), .ZN(n589) );
  INV_X1 U509 ( .A(n589), .ZN(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n454) );
  XNOR2_X1 U511 ( .A(KEYINPUT37), .B(n454), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n291), .B(n455), .ZN(n520) );
  NOR2_X1 U513 ( .A1(n488), .A2(n520), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT38), .ZN(n505) );
  NAND2_X1 U515 ( .A1(n505), .A2(n536), .ZN(n458) );
  XOR2_X1 U516 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n464) );
  XNOR2_X1 U517 ( .A(n459), .B(KEYINPUT41), .ZN(n555) );
  AND2_X1 U518 ( .A1(n563), .A2(n555), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT46), .ZN(n461) );
  NOR2_X1 U520 ( .A1(n566), .A2(n461), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n462), .A2(n548), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(n469) );
  INV_X1 U523 ( .A(n566), .ZN(n586) );
  NOR2_X1 U524 ( .A1(n586), .A2(n589), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT45), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n466), .A2(n459), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n563), .A2(n467), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(n532) );
  AND2_X1 U530 ( .A1(n532), .A2(n525), .ZN(n474) );
  INV_X1 U531 ( .A(KEYINPUT54), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n475), .A2(n521), .ZN(n577) );
  NAND2_X1 U534 ( .A1(n577), .A2(n476), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(KEYINPUT55), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n478), .A2(n536), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n572), .A2(n555), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n484) );
  NAND2_X1 U540 ( .A1(n566), .A2(n548), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  NOR2_X1 U542 ( .A1(n486), .A2(n485), .ZN(n487) );
  XOR2_X1 U543 ( .A(KEYINPUT96), .B(n487), .Z(n510) );
  NOR2_X1 U544 ( .A1(n510), .A2(n488), .ZN(n498) );
  NAND2_X1 U545 ( .A1(n498), .A2(n521), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n489), .B(KEYINPUT97), .ZN(n490) );
  XOR2_X1 U547 ( .A(n490), .B(KEYINPUT98), .Z(n492) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n525), .A2(n498), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n495) );
  NAND2_X1 U553 ( .A1(n498), .A2(n536), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U555 ( .A(G15GAT), .B(n496), .Z(G1326GAT) );
  INV_X1 U556 ( .A(n497), .ZN(n535) );
  NAND2_X1 U557 ( .A1(n535), .A2(n498), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(KEYINPUT100), .ZN(n500) );
  XNOR2_X1 U559 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  NAND2_X1 U560 ( .A1(n505), .A2(n521), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n505), .A2(n525), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n535), .A2(n505), .ZN(n506) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(KEYINPUT108), .ZN(n508) );
  XOR2_X1 U570 ( .A(KEYINPUT107), .B(n508), .Z(n512) );
  NAND2_X1 U571 ( .A1(n555), .A2(n578), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(KEYINPUT106), .ZN(n519) );
  NOR2_X1 U573 ( .A1(n519), .A2(n510), .ZN(n515) );
  NAND2_X1 U574 ( .A1(n515), .A2(n521), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n525), .A2(n515), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n536), .A2(n515), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n535), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n518), .Z(G1335GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n523) );
  NAND2_X1 U585 ( .A1(n528), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n528), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n536), .A2(n528), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n530) );
  NAND2_X1 U593 ( .A1(n528), .A2(n535), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U595 ( .A(n531), .B(G106GAT), .Z(G1339GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n540) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(KEYINPUT114), .B(n534), .ZN(n552) );
  NOR2_X1 U599 ( .A1(n552), .A2(n535), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U601 ( .A(KEYINPUT115), .B(n538), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n549), .A2(n563), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U606 ( .A1(n549), .A2(n555), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n545) );
  NAND2_X1 U610 ( .A1(n549), .A2(n566), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  INV_X1 U614 ( .A(n548), .ZN(n571) );
  NAND2_X1 U615 ( .A1(n549), .A2(n571), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NOR2_X1 U617 ( .A1(n575), .A2(n552), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT120), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n563), .A2(n560), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n555), .A2(n560), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n566), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n571), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT122), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT123), .Z(n568) );
  NAND2_X1 U633 ( .A1(n572), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(KEYINPUT124), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(n570), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1351GAT) );
  INV_X1 U640 ( .A(n575), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n588) );
  NOR2_X1 U642 ( .A1(n578), .A2(n588), .ZN(n582) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT60), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT126), .B(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n459), .A2(n588), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n588), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

