//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G15gat), .B(G22gat), .Z(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G1gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n203), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n207), .B(new_n210), .Z(new_n211));
  XOR2_X1   g010(.A(G43gat), .B(G50gat), .Z(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NOR3_X1   g013(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT87), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT88), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n216), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n221), .A2(KEYINPUT88), .A3(new_n219), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G29gat), .A2(G36gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n214), .B1(new_n220), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n212), .A2(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(KEYINPUT89), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n234), .A3(new_n217), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n231), .B(new_n235), .C1(new_n213), .C2(new_n212), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n229), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n230), .B1(new_n229), .B2(new_n236), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n211), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n207), .B(new_n210), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n229), .A2(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n243), .B(KEYINPUT13), .Z(new_n247));
  INV_X1    g046(.A(new_n242), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n240), .A2(new_n241), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n239), .A2(KEYINPUT18), .A3(new_n242), .A4(new_n243), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT11), .B(G169gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G197gat), .ZN(new_n254));
  XOR2_X1   g053(.A(G113gat), .B(G141gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT12), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n246), .A2(new_n257), .A3(new_n250), .A4(new_n251), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G227gat), .ZN(new_n263));
  INV_X1    g062(.A(G233gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G169gat), .ZN(new_n266));
  INV_X1    g065(.A(G176gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT26), .ZN(new_n269));
  OR3_X1    g068(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n269), .B(new_n270), .C1(new_n266), .C2(new_n267), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT66), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT67), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT27), .B(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n278), .B(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n272), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n284), .A2(KEYINPUT24), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n286));
  NOR2_X1   g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n284), .B2(KEYINPUT24), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n266), .A2(new_n267), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(new_n268), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT65), .B(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT23), .A3(new_n266), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n290), .A2(new_n291), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n285), .A2(new_n288), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n298), .B(new_n294), .C1(new_n293), .C2(new_n268), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT25), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n283), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G113gat), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n303), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT69), .B1(new_n303), .B2(G120gat), .ZN(new_n305));
  INV_X1    g104(.A(G120gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n304), .B(new_n305), .C1(G113gat), .C2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G113gat), .B(G120gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT1), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n312), .A2(new_n309), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n302), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n283), .B2(new_n301), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n265), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT34), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI211_X1 g119(.A(KEYINPUT34), .B(new_n265), .C1(new_n316), .C2(new_n317), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n316), .A2(new_n265), .A3(new_n317), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT33), .ZN(new_n324));
  XNOR2_X1  g123(.A(G15gat), .B(G43gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(G71gat), .ZN(new_n326));
  INV_X1    g125(.A(G99gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n329), .B2(new_n328), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n323), .A2(KEYINPUT32), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n323), .B1(KEYINPUT32), .B2(new_n324), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n328), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n322), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n322), .B1(new_n332), .B2(new_n334), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT36), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340));
  XNOR2_X1  g139(.A(G141gat), .B(G148gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(G155gat), .B2(G162gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n340), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G155gat), .B(G162gat), .Z(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n314), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  AND2_X1   g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n344), .A2(new_n345), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n344), .A2(new_n345), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n353), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n346), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n315), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n346), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n356), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI221_X1 g161(.A(new_n350), .B1(new_n348), .B2(new_n347), .C1(new_n358), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n361), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n315), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n347), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n349), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n363), .A2(KEYINPUT5), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n347), .B(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT4), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n347), .B(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n348), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n358), .A2(new_n362), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n371), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT0), .B(G57gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT77), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n368), .A2(new_n376), .A3(new_n385), .A4(new_n381), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n377), .A2(new_n382), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(KEYINPUT78), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n377), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n383), .A2(new_n388), .A3(new_n384), .A4(new_n386), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT72), .Z(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n302), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT71), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n401));
  OR2_X1    g200(.A1(G197gat), .A2(G204gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n400), .B(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n283), .A2(new_n301), .B1(KEYINPUT29), .B2(new_n396), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n398), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n406), .B1(new_n398), .B2(new_n407), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(G8gat), .B(G36gat), .Z(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G64gat), .ZN(new_n413));
  INV_X1    g212(.A(G92gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n409), .B2(new_n410), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT30), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n411), .A2(new_n420), .A3(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n394), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n424), .B(G22gat), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n356), .B1(new_n405), .B2(KEYINPUT29), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n364), .ZN(new_n428));
  INV_X1    g227(.A(G228gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n264), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT75), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n346), .A2(new_n355), .A3(new_n356), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n428), .B(new_n430), .C1(new_n433), .C2(new_n406), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT79), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT31), .B(G50gat), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n433), .A2(new_n406), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n427), .A2(new_n353), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n430), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n436), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n434), .B(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n439), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n426), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n436), .B1(new_n435), .B2(new_n439), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n441), .A3(new_n444), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n425), .A3(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n446), .A2(KEYINPUT80), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT80), .B1(new_n446), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n339), .B1(new_n423), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(new_n449), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n422), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n349), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT39), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n366), .A2(new_n349), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n458), .B(new_n462), .C1(new_n461), .C2(new_n460), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT81), .B(KEYINPUT39), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n457), .A2(new_n349), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n465), .A3(new_n381), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n377), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n368), .A2(new_n376), .A3(KEYINPUT83), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n382), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT40), .A4(new_n381), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n456), .A2(new_n468), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n390), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n475), .A2(KEYINPUT85), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n472), .A2(new_n384), .A3(new_n383), .A4(new_n386), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(KEYINPUT85), .ZN(new_n478));
  OR3_X1    g277(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT37), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT37), .B1(new_n409), .B2(new_n410), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n479), .A2(new_n415), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n415), .A3(new_n482), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n417), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n455), .B(new_n474), .C1(new_n484), .C2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n387), .A2(new_n472), .B1(KEYINPUT85), .B2(new_n475), .ZN(new_n491));
  INV_X1    g290(.A(new_n487), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n476), .A4(new_n483), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(KEYINPUT86), .A3(new_n455), .A4(new_n474), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n453), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n423), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n335), .A2(new_n336), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(new_n454), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n422), .A3(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n496), .A2(new_n501), .B1(new_n503), .B2(new_n500), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n262), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n506));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G71gat), .B(G78gat), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n240), .B1(KEYINPUT21), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT92), .ZN(new_n513));
  XOR2_X1   g312(.A(G127gat), .B(G155gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(G183gat), .B(G211gat), .Z(new_n516));
  NAND2_X1  g315(.A1(G231gat), .A2(G233gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n515), .B(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n519), .B(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G99gat), .B(G106gat), .Z(new_n524));
  NAND2_X1  g323(.A1(G85gat), .A2(G92gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n414), .ZN(new_n529));
  NAND2_X1  g328(.A1(KEYINPUT93), .A2(G92gat), .ZN(new_n530));
  AOI21_X1  g329(.A(G85gat), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT8), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(G99gat), .B2(G106gat), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT94), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G85gat), .ZN(new_n535));
  AND2_X1   g334(.A1(KEYINPUT93), .A2(G92gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(KEYINPUT93), .A2(G92gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  INV_X1    g338(.A(G106gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT8), .B1(new_n327), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AOI211_X1 g341(.A(new_n524), .B(new_n527), .C1(new_n534), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n524), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n534), .A2(new_n542), .ZN(new_n545));
  INV_X1    g344(.A(new_n527), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n237), .A2(new_n238), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n547), .A2(new_n543), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n241), .ZN(new_n551));
  NAND3_X1  g350(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(KEYINPUT95), .A3(new_n552), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n549), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n556), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT95), .B1(new_n551), .B2(new_n552), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n548), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n558), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n561), .A2(new_n564), .B1(new_n569), .B2(new_n559), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(new_n559), .A3(KEYINPUT96), .A4(new_n564), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n523), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n509), .B(new_n510), .Z(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n547), .B2(new_n543), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n539), .B1(new_n538), .B2(new_n541), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n546), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n524), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n545), .A2(new_n544), .A3(new_n546), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n511), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n576), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n550), .A2(KEYINPUT10), .A3(new_n511), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n576), .A2(new_n582), .A3(KEYINPUT97), .A4(new_n583), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n576), .A2(new_n582), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT98), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(new_n306), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n574), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n505), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(new_n394), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n204), .ZN(G1324gat));
  NOR2_X1   g403(.A1(new_n602), .A2(new_n422), .ZN(new_n605));
  NAND2_X1  g404(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n208), .A2(new_n202), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT42), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n610), .B(new_n611), .C1(new_n202), .C2(new_n605), .ZN(G1325gat));
  INV_X1    g411(.A(G15gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n339), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n602), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n505), .A2(new_n337), .A3(new_n601), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n613), .B2(new_n616), .ZN(G1326gat));
  INV_X1    g416(.A(new_n452), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT43), .B(G22gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT99), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n619), .B(new_n621), .ZN(G1327gat));
  NAND2_X1  g421(.A1(new_n495), .A2(new_n504), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT44), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT96), .B1(new_n557), .B2(new_n558), .ZN(new_n626));
  INV_X1    g425(.A(new_n564), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n557), .A2(new_n558), .ZN(new_n628));
  AOI211_X1 g427(.A(new_n568), .B(new_n549), .C1(new_n555), .C2(new_n556), .ZN(new_n629));
  OAI22_X1  g428(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n625), .B1(new_n630), .B2(new_n571), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n625), .A3(new_n571), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n623), .A2(new_n624), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n573), .B1(new_n495), .B2(new_n504), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n635), .B1(new_n624), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n261), .A2(KEYINPUT100), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n259), .A2(new_n640), .A3(new_n260), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n523), .A2(new_n600), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G29gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n523), .A2(new_n600), .ZN(new_n646));
  INV_X1    g445(.A(new_n573), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n505), .A2(new_n223), .A3(new_n638), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT45), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(G1328gat));
  NAND2_X1  g455(.A1(new_n623), .A2(new_n261), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n648), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n422), .A2(G36gat), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT104), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n637), .A2(new_n456), .A3(new_n643), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G36gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n662), .A2(new_n664), .A3(new_n667), .ZN(G1329gat));
  AOI21_X1  g467(.A(new_n624), .B1(new_n623), .B2(new_n647), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n630), .A2(new_n625), .A3(new_n571), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n631), .ZN(new_n671));
  AOI211_X1 g470(.A(KEYINPUT44), .B(new_n671), .C1(new_n495), .C2(new_n504), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n339), .B(new_n643), .C1(new_n669), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(G43gat), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n657), .A2(G43gat), .A3(new_n497), .A4(new_n648), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT47), .B1(new_n677), .B2(KEYINPUT105), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n675), .B1(new_n673), .B2(G43gat), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n678), .A2(new_n682), .ZN(G1330gat));
  OAI211_X1 g482(.A(new_n454), .B(new_n643), .C1(new_n669), .C2(new_n672), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G50gat), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n618), .A2(G50gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n505), .A2(new_n649), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(KEYINPUT48), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n685), .A2(KEYINPUT107), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT107), .B1(new_n685), .B2(new_n688), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n687), .B(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n637), .A2(new_n452), .A3(new_n643), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(G50gat), .ZN(new_n694));
  OAI22_X1  g493(.A1(new_n689), .A2(new_n690), .B1(new_n694), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g494(.A(new_n574), .B1(new_n495), .B2(new_n504), .ZN(new_n696));
  INV_X1    g495(.A(new_n600), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n639), .A2(new_n641), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n638), .B(KEYINPUT108), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g504(.A(new_n422), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT109), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT110), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n701), .A2(new_n710), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1333gat));
  NAND3_X1  g513(.A1(new_n701), .A2(G71gat), .A3(new_n339), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n497), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(G71gat), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n452), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g519(.A1(new_n523), .A2(new_n698), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n636), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n724), .A2(new_n535), .A3(new_n638), .A4(new_n600), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n600), .B(new_n721), .C1(new_n669), .C2(new_n672), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(new_n394), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1336gat));
  NAND4_X1  g527(.A1(new_n637), .A2(new_n456), .A3(new_n600), .A4(new_n721), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n536), .A2(new_n537), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732));
  INV_X1    g531(.A(new_n724), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n456), .A2(new_n414), .A3(new_n600), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT111), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n722), .A2(KEYINPUT112), .A3(new_n723), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n723), .A2(KEYINPUT112), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n636), .A2(new_n721), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n729), .B2(new_n730), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n736), .B1(new_n732), .B2(new_n741), .ZN(G1337gat));
  NAND4_X1  g541(.A1(new_n724), .A2(new_n327), .A3(new_n337), .A4(new_n600), .ZN(new_n743));
  OAI21_X1  g542(.A(G99gat), .B1(new_n726), .B2(new_n614), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1338gat));
  OAI21_X1  g544(.A(G106gat), .B1(new_n726), .B2(new_n455), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n455), .A2(G106gat), .A3(new_n697), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n733), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n637), .A2(new_n452), .A3(new_n600), .A4(new_n721), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(G106gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n739), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n747), .B(KEYINPUT113), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n749), .A2(new_n750), .B1(new_n752), .B2(new_n755), .ZN(G1339gat));
  NOR3_X1   g555(.A1(new_n574), .A2(new_n600), .A3(new_n698), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758));
  INV_X1    g557(.A(new_n590), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n586), .A2(new_n759), .A3(new_n587), .A4(new_n588), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT54), .B1(new_n760), .B2(KEYINPUT114), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n591), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(new_n760), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n589), .A2(new_n765), .A3(new_n590), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n597), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n758), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n766), .A2(new_n597), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT114), .B1(new_n589), .B2(new_n590), .ZN(new_n770));
  INV_X1    g569(.A(new_n760), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n769), .B(KEYINPUT55), .C1(new_n772), .C2(new_n761), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n698), .A2(new_n598), .A3(new_n768), .A4(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n248), .A2(new_n249), .A3(new_n247), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n243), .B1(new_n239), .B2(new_n242), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n256), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n260), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n600), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT116), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n774), .A2(new_n782), .A3(new_n779), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n671), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n598), .A3(new_n778), .A4(new_n773), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n634), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT115), .B1(new_n671), .B2(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n523), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n757), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n497), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n638), .A2(new_n422), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(new_n618), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(G113gat), .B1(new_n797), .B2(new_n262), .ZN(new_n798));
  NOR4_X1   g597(.A1(new_n793), .A2(new_n499), .A3(new_n456), .A4(new_n702), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n303), .A3(new_n698), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1340gat));
  OAI21_X1  g600(.A(G120gat), .B1(new_n797), .B2(new_n697), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n306), .A3(new_n600), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1341gat));
  INV_X1    g603(.A(G127gat), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n797), .A2(new_n805), .A3(new_n792), .ZN(new_n806));
  AOI21_X1  g605(.A(G127gat), .B1(new_n799), .B2(new_n523), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(G1342gat));
  INV_X1    g607(.A(G134gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n799), .A2(new_n809), .A3(new_n647), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT56), .Z(new_n811));
  OAI21_X1  g610(.A(G134gat), .B1(new_n797), .B2(new_n573), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1343gat));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n614), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n774), .A2(new_n782), .A3(new_n779), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n782), .B1(new_n774), .B2(new_n779), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(new_n634), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n788), .A2(new_n789), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n792), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n757), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n455), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n814), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n779), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n769), .B(KEYINPUT117), .C1(new_n772), .C2(new_n761), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n758), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n771), .A2(new_n762), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(KEYINPUT54), .C1(new_n771), .C2(new_n770), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT117), .B1(new_n828), .B2(new_n769), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n598), .B(new_n773), .C1(new_n826), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n262), .B1(new_n830), .B2(KEYINPUT118), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n773), .A2(new_n598), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n832), .B(new_n833), .C1(new_n829), .C2(new_n826), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n824), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n790), .B1(new_n835), .B2(new_n647), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n757), .B1(new_n836), .B2(new_n792), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT57), .B1(new_n837), .B2(new_n618), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G141gat), .B1(new_n839), .B2(new_n262), .ZN(new_n840));
  XNOR2_X1  g639(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n702), .B1(new_n819), .B2(new_n820), .ZN(new_n842));
  INV_X1    g641(.A(G141gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n614), .A2(new_n454), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n842), .A2(new_n843), .A3(new_n422), .A4(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n840), .B(new_n841), .C1(new_n262), .C2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n823), .A2(new_n838), .A3(new_n698), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n848), .A2(KEYINPUT119), .A3(G141gat), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT119), .B1(new_n848), .B2(G141gat), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n846), .B2(new_n262), .ZN(new_n852));
  NOR4_X1   g651(.A1(new_n793), .A2(new_n456), .A3(new_n702), .A4(new_n844), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n853), .A2(KEYINPUT120), .A3(new_n843), .A4(new_n261), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n849), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n847), .B1(new_n856), .B2(new_n857), .ZN(G1344gat));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n859), .B(G148gat), .C1(new_n853), .C2(new_n600), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT57), .B1(new_n793), .B2(new_n455), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n785), .A2(new_n573), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n835), .B2(new_n647), .ZN(new_n864));
  AOI22_X1  g663(.A1(new_n864), .A2(new_n792), .B1(new_n262), .B2(new_n601), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n452), .A2(new_n822), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n859), .B(new_n697), .C1(new_n814), .C2(KEYINPUT122), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n868), .B(new_n869), .C1(KEYINPUT122), .C2(new_n814), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n859), .B1(new_n839), .B2(new_n697), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n860), .B1(new_n872), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g672(.A(G155gat), .B1(new_n853), .B2(new_n523), .ZN(new_n874));
  INV_X1    g673(.A(new_n839), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n523), .A2(G155gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(G1346gat));
  OAI21_X1  g676(.A(G162gat), .B1(new_n839), .B2(new_n671), .ZN(new_n878));
  INV_X1    g677(.A(G162gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n853), .A2(new_n879), .A3(new_n647), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n793), .A2(new_n638), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n499), .A2(new_n422), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n266), .A3(new_n698), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n702), .A2(new_n456), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n794), .A2(new_n618), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G169gat), .B1(new_n889), .B2(new_n262), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n886), .A2(new_n890), .ZN(G1348gat));
  AOI21_X1  g690(.A(G176gat), .B1(new_n885), .B2(new_n600), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n889), .A2(new_n295), .A3(new_n697), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(G1349gat));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  OAI21_X1  g694(.A(G183gat), .B1(new_n889), .B2(new_n792), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n882), .A2(new_n279), .A3(new_n523), .A4(new_n883), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AND4_X1   g698(.A1(new_n618), .A2(new_n794), .A3(new_n523), .A4(new_n888), .ZN(new_n900));
  INV_X1    g699(.A(G183gat), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n895), .B(new_n897), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(KEYINPUT60), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n904));
  INV_X1    g703(.A(new_n902), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n898), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n889), .B2(new_n573), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT61), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n885), .A2(new_n280), .A3(new_n634), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1351gat));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n867), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n861), .B(KEYINPUT125), .C1(new_n865), .C2(new_n866), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n887), .A2(new_n339), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n913), .A2(new_n914), .A3(new_n261), .A4(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n915), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n867), .B2(new_n912), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n920), .A2(KEYINPUT126), .A3(new_n261), .A4(new_n914), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n921), .A3(G197gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n844), .A2(new_n422), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT124), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT124), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n882), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n926), .A2(G197gat), .A3(new_n642), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n922), .A2(new_n927), .ZN(G1352gat));
  NOR3_X1   g727(.A1(new_n926), .A2(G204gat), .A3(new_n697), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n920), .A2(new_n600), .A3(new_n914), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G204gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1353gat));
  OR3_X1    g732(.A1(new_n926), .A2(G211gat), .A3(new_n792), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n868), .A2(new_n523), .A3(new_n915), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n647), .A3(new_n914), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G218gat), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n926), .A2(G218gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n671), .B2(new_n941), .ZN(G1355gat));
endmodule


