//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT77), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n193), .A3(KEYINPUT77), .A4(new_n194), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(G101), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n190), .A2(new_n193), .A3(new_n200), .A4(new_n194), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n201), .A2(KEYINPUT4), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT78), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n199), .A2(KEYINPUT4), .ZN(new_n205));
  INV_X1    g019(.A(G116), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G116), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT65), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(G116), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G119), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  AND3_X1   g029(.A1(KEYINPUT64), .A2(KEYINPUT2), .A3(G113), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n216), .A2(new_n217), .B1(KEYINPUT2), .B2(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(new_n212), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT78), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n199), .A2(new_n224), .A3(new_n202), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n204), .A2(new_n205), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n210), .A2(KEYINPUT5), .A3(new_n214), .ZN(new_n227));
  INV_X1    g041(.A(G113), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n207), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n192), .A2(KEYINPUT79), .A3(G104), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n192), .B2(G104), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n189), .A2(G107), .ZN(new_n235));
  OAI211_X1 g049(.A(G101), .B(new_n232), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n201), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n222), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n231), .A2(new_n238), .A3(KEYINPUT82), .A4(new_n222), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g057(.A(G110), .B(G122), .Z(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n226), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n231), .A2(new_n222), .A3(new_n237), .ZN(new_n247));
  XOR2_X1   g061(.A(new_n244), .B(KEYINPUT8), .Z(new_n248));
  NAND3_X1  g062(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT5), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n221), .B1(new_n230), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n247), .B(new_n248), .C1(new_n237), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G143), .B(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n257), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(G125), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G224), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n263), .A2(KEYINPUT85), .B1(KEYINPUT7), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT1), .B1(new_n254), .B2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n256), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n261), .A2(new_n270), .A3(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n263), .B1(new_n272), .B2(G125), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n266), .B(new_n273), .Z(new_n274));
  NAND3_X1  g088(.A1(new_n246), .A2(new_n251), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n226), .A2(new_n243), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n244), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT83), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n245), .B1(new_n226), .B2(new_n243), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT83), .A3(new_n280), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n280), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n283), .A2(new_n285), .B1(new_n286), .B2(new_n246), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n273), .B(new_n265), .Z(new_n288));
  AOI21_X1  g102(.A(KEYINPUT84), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n279), .A2(new_n244), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT6), .A3(new_n246), .ZN(new_n291));
  AND4_X1   g105(.A1(KEYINPUT83), .A2(new_n279), .A3(new_n280), .A4(new_n244), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT83), .B1(new_n284), .B2(new_n280), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n288), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n278), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT86), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n294), .A2(new_n295), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n283), .A2(new_n285), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n303), .A2(KEYINPUT84), .A3(new_n288), .A4(new_n291), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n277), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n298), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n188), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G217), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(G234), .B2(new_n276), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G128), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G119), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n208), .A2(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OR2_X1    g131(.A1(KEYINPUT24), .A2(G110), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT24), .A2(G110), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n315), .A2(new_n312), .ZN(new_n321));
  OAI22_X1  g135(.A1(new_n317), .A2(G110), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(G125), .A2(G140), .ZN(new_n326));
  NOR2_X1   g140(.A1(G125), .A2(G140), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT16), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n328), .A3(G146), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(G125), .A2(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n252), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n317), .A2(G110), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT16), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n331), .B2(new_n332), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n339), .A2(new_n252), .A3(new_n324), .ZN(new_n340));
  AOI21_X1  g154(.A(G146), .B1(new_n325), .B2(new_n328), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n318), .A2(new_n315), .A3(new_n312), .A4(new_n319), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT70), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n252), .B1(new_n339), .B2(new_n324), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n347), .A2(new_n329), .B1(G110), .B2(new_n317), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT70), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n343), .B(KEYINPUT69), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n336), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT22), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(G137), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT71), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n342), .A2(new_n345), .A3(KEYINPUT70), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n349), .B1(new_n348), .B2(new_n350), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n335), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT71), .ZN(new_n360));
  INV_X1    g174(.A(new_n355), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n335), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n352), .A2(KEYINPUT72), .A3(new_n355), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n363), .A2(new_n368), .A3(new_n276), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT73), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT25), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n363), .A2(new_n368), .A3(KEYINPUT25), .A4(new_n276), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT74), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n310), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT11), .ZN(new_n379));
  INV_X1    g193(.A(G134), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(G137), .ZN(new_n381));
  INV_X1    g195(.A(G137), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT11), .A3(G134), .ZN(new_n383));
  INV_X1    g197(.A(G131), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(G137), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n381), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n382), .A2(G134), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n380), .A2(G137), .ZN(new_n388));
  OAI21_X1  g202(.A(G131), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT66), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n272), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n381), .A2(new_n385), .A3(new_n383), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G131), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n386), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n260), .A2(new_n262), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n378), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n390), .B1(new_n269), .B2(new_n271), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n396), .A2(new_n386), .B1(new_n260), .B2(new_n262), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT30), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n223), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n221), .B1(new_n215), .B2(new_n218), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n394), .A2(new_n405), .A3(new_n399), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(G101), .ZN(new_n408));
  NOR2_X1   g222(.A1(G237), .A2(G953), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G210), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n408), .B(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT31), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT31), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n404), .A2(new_n414), .A3(new_n406), .A4(new_n411), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT67), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT28), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n406), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n223), .B1(new_n401), .B2(new_n402), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n406), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n416), .B1(new_n406), .B2(new_n417), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n413), .B(new_n415), .C1(new_n423), .C2(new_n411), .ZN(new_n424));
  NOR2_X1   g238(.A1(G472), .A2(G902), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT32), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT32), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n428), .A3(new_n425), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n394), .A2(new_n405), .A3(new_n399), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n405), .B1(new_n394), .B2(new_n399), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT28), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n430), .C2(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n421), .ZN(new_n437));
  INV_X1    g251(.A(new_n422), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT29), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .A4(new_n418), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n419), .A2(new_n422), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n436), .A2(new_n440), .A3(new_n411), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n411), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n404), .A2(new_n406), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n440), .B2(new_n411), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n442), .B(new_n276), .C1(new_n445), .C2(KEYINPUT29), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n427), .A2(new_n429), .B1(new_n446), .B2(G472), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n363), .A2(new_n368), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n449), .A2(G902), .A3(new_n309), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n377), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n409), .A2(G214), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n254), .A2(KEYINPUT87), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n384), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n452), .B1(KEYINPUT87), .B2(new_n254), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n453), .B1(G214), .B2(new_n409), .ZN(new_n458));
  OAI21_X1  g272(.A(G131), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n340), .A2(new_n341), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n460), .B(new_n461), .C1(new_n456), .C2(new_n459), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT18), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n454), .B1(new_n463), .B2(new_n384), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n333), .B(new_n252), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n464), .B(new_n465), .C1(new_n463), .C2(new_n459), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(G113), .B(G122), .Z(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT88), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n189), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n462), .A2(new_n470), .A3(new_n466), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n276), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n475), .A2(G475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n455), .A2(new_n459), .ZN(new_n477));
  XOR2_X1   g291(.A(new_n333), .B(KEYINPUT19), .Z(new_n478));
  OAI21_X1  g292(.A(new_n329), .B1(new_n478), .B2(G146), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n466), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n471), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n473), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n473), .A3(KEYINPUT89), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT20), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(KEYINPUT90), .B2(KEYINPUT20), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n482), .B(new_n489), .C1(KEYINPUT90), .C2(new_n485), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n476), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n264), .A2(G952), .ZN(new_n492));
  NAND2_X1  g306(.A1(G234), .A2(G237), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT21), .B(G898), .Z(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(G902), .A3(G953), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n311), .A2(G143), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n254), .A2(G128), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n380), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n498), .A2(KEYINPUT13), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT93), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n499), .B1(KEYINPUT13), .B2(new_n498), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT91), .B1(new_n206), .B2(G122), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n507));
  INV_X1    g321(.A(G122), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(G116), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n206), .A2(G122), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n510), .A2(KEYINPUT92), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT92), .B1(new_n510), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n192), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n512), .A2(new_n513), .A3(new_n192), .ZN(new_n516));
  OAI221_X1 g330(.A(new_n501), .B1(new_n505), .B2(new_n380), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n511), .B(KEYINPUT14), .ZN(new_n518));
  INV_X1    g332(.A(new_n510), .ZN(new_n519));
  OAI21_X1  g333(.A(G107), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n500), .B(new_n380), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT94), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n514), .A2(new_n524), .A3(new_n520), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT9), .B(G234), .Z(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n528), .A2(new_n308), .A3(G953), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n517), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n529), .B1(new_n517), .B2(new_n526), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n276), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G478), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n532), .A2(new_n534), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n491), .A2(new_n497), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G469), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n264), .A2(G227), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n330), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT75), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(G110), .Z(new_n543));
  NAND4_X1  g357(.A1(new_n204), .A2(new_n205), .A3(new_n398), .A4(new_n225), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT81), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT80), .B(KEYINPUT1), .C1(new_n254), .C2(G146), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G128), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT80), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n256), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n237), .B1(new_n271), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n545), .B1(new_n550), .B2(KEYINPUT10), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n256), .A2(KEYINPUT1), .A3(new_n311), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT80), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n267), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(G128), .A3(new_n546), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n553), .B1(new_n256), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT81), .B(new_n552), .C1(new_n557), .C2(new_n237), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n238), .A2(new_n272), .A3(KEYINPUT10), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n544), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n397), .ZN(new_n562));
  INV_X1    g376(.A(new_n397), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n544), .A2(new_n559), .A3(new_n563), .A4(new_n560), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n543), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n238), .A2(new_n272), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n397), .B1(new_n566), .B2(new_n550), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g383(.A(KEYINPUT12), .B(new_n397), .C1(new_n566), .C2(new_n550), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n564), .A2(new_n543), .A3(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n539), .B(new_n276), .C1(new_n565), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(G469), .A2(G902), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n564), .A2(new_n571), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n543), .A2(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n543), .A2(KEYINPUT76), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n562), .A2(new_n564), .A3(new_n543), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(G469), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G221), .B1(new_n528), .B2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n307), .A2(new_n451), .A3(new_n538), .A4(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  AOI21_X1  g400(.A(KEYINPUT95), .B1(new_n305), .B2(new_n298), .ZN(new_n587));
  INV_X1    g401(.A(new_n298), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n297), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n588), .B(new_n277), .C1(new_n302), .C2(new_n304), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n188), .B1(new_n591), .B2(KEYINPUT95), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n377), .A2(new_n450), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n424), .A2(new_n276), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n581), .A2(new_n597), .A3(new_n426), .A4(new_n582), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n593), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT97), .B1(new_n530), .B2(new_n531), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n531), .A2(KEYINPUT97), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT33), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n530), .B2(new_n531), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n602), .A2(G478), .A3(new_n276), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n532), .A2(new_n533), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n491), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n497), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n599), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  OR2_X1    g428(.A1(new_n487), .A2(KEYINPUT20), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n476), .B1(new_n615), .B2(new_n488), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n536), .A2(new_n535), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n610), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT98), .Z(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n599), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT99), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n621), .B(new_n623), .ZN(G9));
  NAND2_X1  g438(.A1(new_n597), .A2(new_n426), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n369), .A2(new_n371), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT73), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n448), .A2(KEYINPUT74), .A3(KEYINPUT25), .A4(new_n276), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT74), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n375), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n627), .A2(new_n628), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n309), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n361), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n359), .B(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n635), .A2(G902), .A3(new_n309), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n625), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n307), .A2(new_n538), .A3(new_n584), .A4(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT37), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G110), .ZN(G12));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  OR3_X1    g456(.A1(new_n496), .A2(new_n642), .A3(G900), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n642), .B1(new_n496), .B2(G900), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n494), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n618), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n590), .A2(new_n647), .A3(new_n592), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT101), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n590), .A2(new_n592), .A3(new_n650), .A4(new_n647), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n633), .A2(new_n637), .ZN(new_n652));
  INV_X1    g466(.A(new_n447), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n584), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n649), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  NAND2_X1  g471(.A1(new_n301), .A2(new_n306), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT102), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n305), .A2(new_n299), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n591), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n659), .A2(new_n663), .A3(KEYINPUT38), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT38), .B1(new_n659), .B2(new_n663), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n491), .B1(new_n535), .B2(new_n536), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n427), .A2(new_n429), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n443), .B1(new_n430), .B2(new_n431), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(KEYINPUT103), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n412), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(KEYINPUT103), .B2(new_n668), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n664), .A2(new_n665), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n652), .A2(new_n188), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n645), .B(KEYINPUT39), .Z(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n584), .A2(KEYINPUT104), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n583), .B2(new_n678), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n680), .A2(KEYINPUT40), .A3(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n659), .A2(new_n663), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT38), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n659), .A2(new_n663), .A3(KEYINPUT38), .ZN(new_n692));
  INV_X1    g506(.A(new_n674), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n687), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n677), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT105), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n254), .ZN(G45));
  NAND3_X1  g512(.A1(new_n607), .A2(new_n608), .A3(new_n645), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n593), .A2(new_n654), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT106), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n252), .ZN(G48));
  INV_X1    g516(.A(new_n451), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n276), .B1(new_n565), .B2(new_n572), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n582), .A3(new_n573), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n593), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n611), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n620), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  AOI21_X1  g529(.A(new_n636), .B1(new_n632), .B2(new_n309), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n716), .A2(new_n447), .A3(new_n537), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n592), .A3(new_n590), .A4(new_n708), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  AND4_X1   g533(.A1(new_n592), .A2(new_n708), .A3(new_n590), .A4(new_n666), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n377), .B2(new_n450), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n436), .A2(new_n441), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n443), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n413), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT108), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n724), .A2(new_n727), .A3(new_n413), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n415), .A3(new_n728), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n729), .A2(new_n425), .B1(G472), .B2(new_n596), .ZN(new_n730));
  INV_X1    g544(.A(new_n450), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n633), .A2(KEYINPUT109), .A3(new_n731), .ZN(new_n732));
  AND4_X1   g546(.A1(new_n497), .A2(new_n722), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n720), .A2(new_n733), .A3(KEYINPUT110), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n708), .A2(new_n590), .A3(new_n592), .A4(new_n666), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n722), .A2(new_n730), .A3(new_n732), .A4(new_n497), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT111), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n508), .ZN(G24));
  INV_X1    g555(.A(new_n593), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n730), .A2(new_n652), .ZN(new_n743));
  INV_X1    g557(.A(new_n699), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n708), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n661), .A3(new_n187), .A4(new_n584), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n722), .A2(new_n653), .A3(new_n732), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT42), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n301), .A2(new_n187), .A3(new_n306), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n699), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n451), .A4(new_n584), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n384), .ZN(G33));
  INV_X1    g569(.A(new_n750), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n451), .A3(new_n584), .A4(new_n647), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT112), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NAND2_X1  g573(.A1(new_n607), .A2(new_n491), .ZN(new_n760));
  NOR2_X1   g574(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n761), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n625), .B(new_n652), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n750), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n578), .A2(new_n579), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(G469), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n574), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(G469), .C1(new_n770), .C2(G902), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n573), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n582), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n678), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n768), .B(new_n777), .C1(new_n767), .C2(new_n766), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n582), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n594), .A2(new_n653), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n751), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  NOR2_X1   g600(.A1(G952), .A2(G953), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT119), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n705), .A2(new_n573), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n781), .B(new_n782), .C1(new_n582), .C2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n765), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n494), .B1(new_n791), .B2(new_n762), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n722), .A2(new_n732), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n792), .A2(new_n793), .A3(new_n730), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n790), .A2(new_n794), .A3(new_n756), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n188), .B1(new_n664), .B2(new_n665), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n792), .A2(new_n708), .A3(new_n793), .A4(new_n730), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT117), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT50), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT117), .B(new_n800), .C1(new_n796), .C2(new_n797), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n795), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n709), .A2(new_n750), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n792), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT118), .Z(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n743), .ZN(new_n806));
  INV_X1    g620(.A(new_n803), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n807), .A2(new_n595), .A3(new_n494), .A4(new_n673), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n491), .A3(new_n606), .A4(new_n605), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n802), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n802), .A2(KEYINPUT51), .A3(new_n806), .A4(new_n809), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n812), .A2(new_n492), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n794), .A2(new_n742), .A3(new_n708), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n808), .A2(new_n608), .A3(new_n607), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n590), .A2(new_n592), .A3(new_n666), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n645), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n377), .A2(new_n636), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n645), .A2(new_n819), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n822), .A3(new_n584), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n820), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n716), .A2(new_n584), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT116), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n818), .A2(new_n824), .A3(new_n673), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n742), .A2(new_n655), .A3(new_n744), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n656), .A2(new_n828), .A3(new_n745), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n654), .B1(new_n648), .B2(KEYINPUT101), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n700), .B1(new_n651), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n745), .A4(new_n828), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n710), .B1(new_n620), .B2(new_n611), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n377), .A2(new_n598), .A3(new_n450), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n617), .A2(new_n491), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n609), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n307), .A2(new_n838), .A3(new_n497), .A4(new_n840), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n585), .A2(new_n718), .A3(new_n841), .A4(new_n639), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n739), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n743), .A2(new_n751), .A3(new_n584), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n749), .A2(new_n753), .A3(new_n844), .A4(new_n757), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n617), .A2(new_n646), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n756), .A2(new_n616), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n756), .A2(KEYINPUT114), .A3(new_n616), .A4(new_n846), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n655), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n843), .A2(new_n845), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT53), .B1(new_n836), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n831), .A2(new_n835), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n718), .A2(new_n585), .A3(new_n841), .A4(new_n639), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n738), .B2(new_n734), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n749), .A2(new_n753), .A3(new_n844), .A4(new_n757), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n837), .A4(new_n851), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n855), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n817), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n836), .A2(new_n853), .A3(KEYINPUT53), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n860), .B1(new_n855), .B2(new_n859), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(KEYINPUT54), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n748), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n805), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT48), .Z(new_n870));
  OAI21_X1  g684(.A(new_n788), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n789), .B(KEYINPUT49), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n673), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n582), .B(new_n873), .C1(new_n664), .C2(new_n665), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n188), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n491), .A3(new_n607), .A4(new_n793), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(G75));
  NOR2_X1   g691(.A1(new_n264), .A2(G952), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n287), .B(new_n288), .Z(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT55), .Z(new_n880));
  AOI21_X1  g694(.A(new_n276), .B1(new_n863), .B2(new_n864), .ZN(new_n881));
  AOI211_X1 g695(.A(KEYINPUT56), .B(new_n880), .C1(new_n881), .C2(new_n300), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  INV_X1    g698(.A(new_n880), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n878), .B(new_n882), .C1(new_n886), .C2(new_n887), .ZN(G51));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n574), .B(KEYINPUT57), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n866), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n890), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n862), .A2(KEYINPUT121), .A3(new_n865), .A4(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n891), .B(new_n893), .C1(new_n565), .C2(new_n572), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n881), .A2(G469), .A3(new_n770), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n878), .B1(new_n894), .B2(new_n895), .ZN(G54));
  AND3_X1   g710(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n484), .A2(new_n486), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n878), .ZN(G60));
  INV_X1    g715(.A(new_n878), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n602), .A2(new_n604), .ZN(new_n903));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT59), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n862), .A2(new_n903), .A3(new_n865), .A4(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n906), .A2(KEYINPUT122), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(KEYINPUT122), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n902), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n862), .A2(new_n865), .A3(new_n905), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n911));
  INV_X1    g725(.A(new_n903), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n909), .A2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(new_n863), .A2(new_n864), .ZN(new_n917));
  INV_X1    g731(.A(new_n635), .ZN(new_n918));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT60), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n863), .B2(new_n864), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n922), .B(new_n902), .C1(new_n448), .C2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g739(.A(new_n264), .B1(new_n495), .B2(G224), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n843), .B2(new_n264), .ZN(new_n927));
  INV_X1    g741(.A(G898), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n287), .B1(new_n928), .B2(G953), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n927), .B(new_n929), .ZN(G69));
  NOR2_X1   g744(.A1(new_n400), .A2(new_n403), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n478), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n833), .A2(new_n745), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n688), .A2(new_n933), .A3(new_n696), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n688), .A2(new_n933), .A3(new_n696), .A4(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n683), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n756), .A3(new_n451), .A4(new_n840), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n778), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n778), .A2(KEYINPUT124), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n938), .A2(new_n785), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n932), .B1(new_n946), .B2(new_n264), .ZN(new_n947));
  INV_X1    g761(.A(new_n785), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n777), .A2(new_n818), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n868), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n933), .A2(new_n778), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n749), .A2(new_n753), .A3(new_n757), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT126), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n950), .A2(new_n951), .A3(new_n264), .A4(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(G900), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n954), .B(new_n932), .C1(new_n955), .C2(new_n264), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n947), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(G227), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n960), .B2(new_n955), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G72));
  INV_X1    g776(.A(new_n843), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n938), .A2(new_n785), .A3(new_n963), .A4(new_n945), .ZN(new_n964));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n443), .B1(new_n404), .B2(new_n406), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n963), .A2(new_n950), .A3(new_n951), .A4(new_n953), .ZN(new_n970));
  INV_X1    g784(.A(new_n966), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n444), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n444), .A2(new_n968), .A3(new_n971), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n917), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n969), .A2(new_n902), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT127), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n878), .B1(new_n967), .B2(new_n968), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n977), .A2(new_n978), .A3(new_n972), .A4(new_n974), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(G57));
endmodule


