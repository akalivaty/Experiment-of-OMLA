//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n205), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT66), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n205), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT64), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n214), .B(new_n224), .C1(KEYINPUT1), .C2(new_n212), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  INV_X1    g0036(.A(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(G50), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G222), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(G223), .A3(G1698), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n251), .B(new_n252), .C1(new_n202), .C2(new_n249), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  AOI21_X1  g0057(.A(G1), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n260), .A3(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G41), .A2(G45), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT69), .B1(new_n262), .B2(G1), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n264), .B(new_n265), .C1(G41), .C2(G45), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n263), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n261), .B1(new_n267), .B2(G226), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n255), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G169), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n272), .A2(new_n222), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT70), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(new_n205), .B2(new_n246), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT71), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(new_n221), .A3(new_n246), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n221), .A2(G33), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n283), .A2(new_n284), .B1(new_n221), .B2(new_n201), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n276), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n275), .A2(new_n222), .A3(new_n287), .A4(new_n272), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n265), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(KEYINPUT72), .A3(G50), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(KEYINPUT72), .B1(new_n289), .B2(G50), .ZN(new_n292));
  OR3_X1    g0092(.A1(new_n288), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n287), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n286), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n271), .B(new_n297), .C1(G179), .C2(new_n269), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n255), .A2(G190), .A3(new_n268), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n286), .A2(new_n293), .A3(KEYINPUT9), .A4(new_n296), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n269), .A2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n302), .A2(new_n308), .A3(new_n303), .A4(new_n305), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n299), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT74), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n249), .A2(G232), .A3(new_n250), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n249), .A2(G238), .A3(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(G107), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n249), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n254), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n261), .B1(new_n267), .B2(G244), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n270), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n280), .A2(new_n283), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT15), .B(G87), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n321), .A2(new_n284), .B1(new_n221), .B2(new_n202), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n276), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n288), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(G77), .A3(new_n289), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n323), .B(new_n325), .C1(G77), .C2(new_n287), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n316), .A2(new_n327), .A3(new_n317), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n319), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n318), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n316), .A2(KEYINPUT73), .A3(G190), .A4(new_n317), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n326), .B1(G200), .B2(new_n318), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n310), .A2(new_n311), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n311), .B1(new_n310), .B2(new_n336), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT75), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(KEYINPUT12), .ZN(new_n342));
  INV_X1    g0142(.A(G68), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n265), .A2(new_n343), .A3(G13), .A4(G20), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(KEYINPUT12), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT76), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n346), .B(KEYINPUT76), .C1(KEYINPUT12), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n289), .A2(G68), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n348), .C1(new_n288), .C2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n280), .A2(new_n295), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n284), .A2(new_n202), .B1(new_n221), .B2(G68), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n276), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT11), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(new_n276), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n350), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n258), .A2(new_n260), .A3(G274), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n263), .A2(G238), .A3(new_n260), .A4(new_n266), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G226), .A2(G1698), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n228), .B2(G1698), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n249), .B1(G33), .B2(G97), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n358), .B(new_n359), .C1(new_n362), .C2(new_n260), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G97), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n228), .A2(G1698), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G226), .B2(G1698), .ZN(new_n367));
  AND2_X1   g0167(.A1(KEYINPUT3), .A2(G33), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT3), .A2(G33), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n365), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n261), .B1(new_n371), .B2(new_n254), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT13), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n359), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n364), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n357), .B1(new_n331), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n364), .B2(new_n374), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n357), .ZN(new_n381));
  NAND2_X1  g0181(.A1(KEYINPUT77), .A2(KEYINPUT14), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n375), .A2(G169), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n364), .A2(new_n374), .A3(G179), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n382), .B1(new_n375), .B2(G169), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n247), .A2(new_n221), .A3(new_n248), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n248), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n343), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g0194(.A(G58), .B(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G20), .ZN(new_n396));
  INV_X1    g0196(.A(G159), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(new_n280), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n389), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n370), .B2(new_n221), .ZN(new_n400));
  INV_X1    g0200(.A(new_n393), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n278), .A2(new_n279), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n403), .A2(G159), .B1(new_n395), .B2(G20), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(new_n405), .A3(new_n276), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n283), .B1(new_n265), .B2(G20), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n324), .A2(new_n407), .B1(new_n294), .B2(new_n283), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n263), .A2(G232), .A3(new_n260), .A4(new_n266), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G223), .A2(G1698), .ZN(new_n411));
  INV_X1    g0211(.A(G226), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(G1698), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n249), .B1(G33), .B2(G87), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n358), .B(new_n410), .C1(new_n414), .C2(new_n260), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n327), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G223), .B2(G1698), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n419), .B2(new_n370), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n261), .B1(new_n420), .B2(new_n254), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n270), .B1(new_n421), .B2(new_n410), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT78), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n415), .A2(G169), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT78), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(new_n425), .C1(new_n327), .C2(new_n415), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n409), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n415), .A2(new_n377), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G190), .B2(new_n415), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n406), .A3(new_n408), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n430), .A2(new_n406), .A3(KEYINPUT17), .A4(new_n408), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n409), .A2(new_n423), .A3(new_n426), .A4(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n428), .A2(new_n433), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n388), .B1(KEYINPUT79), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n437), .A2(KEYINPUT79), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT80), .B1(new_n340), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n310), .A2(new_n336), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT74), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n337), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT80), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n439), .A4(new_n438), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT20), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n449), .A2(KEYINPUT84), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(KEYINPUT84), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  INV_X1    g0252(.A(G97), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n221), .C1(G33), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n275), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n272), .A2(new_n222), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n457), .A2(new_n458), .B1(new_n221), .B2(G116), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n450), .B(new_n451), .C1(new_n456), .C2(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n454), .B(KEYINPUT83), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n273), .A2(new_n275), .B1(G20), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n461), .A2(KEYINPUT84), .A3(new_n463), .A4(new_n449), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n287), .A2(G116), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n246), .A2(G1), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n288), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n467), .B2(G116), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n460), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n257), .A2(G1), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n254), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n260), .A2(G274), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n265), .A2(G45), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n471), .B2(new_n472), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n474), .A2(G270), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G264), .B(G1698), .C1(new_n368), .C2(new_n369), .ZN(new_n480));
  OAI211_X1 g0280(.A(G257), .B(new_n250), .C1(new_n368), .C2(new_n369), .ZN(new_n481));
  INV_X1    g0281(.A(G303), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(new_n481), .C1(new_n482), .C2(new_n249), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n254), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n270), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n469), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI211_X1 g0288(.A(new_n487), .B(new_n270), .C1(new_n479), .C2(new_n484), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n479), .A2(new_n484), .A3(G179), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n469), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n464), .A2(new_n468), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n479), .A2(new_n484), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G200), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n479), .A2(new_n484), .A3(G190), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n492), .A2(new_n494), .A3(new_n460), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n488), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(KEYINPUT85), .A2(G294), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT85), .A2(G294), .ZN(new_n499));
  OAI21_X1  g0299(.A(G33), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G257), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G1698), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G250), .B2(G1698), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n500), .B1(new_n503), .B2(new_n370), .ZN(new_n504));
  AOI22_X1  g0304(.A1(G264), .A2(new_n474), .B1(new_n504), .B2(new_n254), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT86), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n478), .A2(G274), .A3(new_n260), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n331), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n254), .ZN(new_n509));
  INV_X1    g0309(.A(new_n472), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n470), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(G264), .A3(new_n260), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n509), .A2(new_n331), .A3(new_n507), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT86), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n507), .A3(new_n513), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n377), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n508), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n221), .B(G87), .C1(new_n368), .C2(new_n369), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT22), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT22), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n249), .A2(new_n521), .A3(new_n221), .A4(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT24), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n246), .A2(new_n462), .A3(G20), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n221), .B2(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n314), .A2(KEYINPUT23), .A3(G20), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n524), .B1(new_n523), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n276), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n294), .A2(new_n314), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n533), .B(KEYINPUT25), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(G107), .B2(new_n467), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n518), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n505), .A2(new_n327), .A3(new_n507), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n516), .A2(new_n270), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n532), .B2(new_n535), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT87), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(new_n535), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n537), .A3(new_n538), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n518), .A2(new_n532), .A3(new_n535), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT87), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g0348(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n221), .B1(new_n549), .B2(new_n365), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  INV_X1    g0351(.A(G87), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n249), .A2(new_n221), .A3(G68), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n221), .A2(G33), .A3(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n276), .B1(new_n294), .B2(new_n321), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(G1698), .C1(new_n368), .C2(new_n369), .ZN(new_n560));
  OAI211_X1 g0360(.A(G238), .B(new_n250), .C1(new_n368), .C2(new_n369), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n246), .C2(new_n462), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n254), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n260), .A2(G250), .A3(new_n477), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n475), .B2(new_n477), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G200), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n467), .A2(G87), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n565), .B1(new_n562), .B2(new_n254), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G190), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n559), .A2(new_n568), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n276), .ZN(new_n573));
  OAI21_X1  g0373(.A(G107), .B1(new_n400), .B2(new_n401), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT6), .ZN(new_n575));
  AND2_X1   g0375(.A1(G97), .A2(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(new_n551), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n314), .A2(KEYINPUT6), .A3(G97), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(G20), .B1(G77), .B2(new_n403), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n573), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n467), .A2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n287), .A2(G97), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(new_n250), .C1(new_n368), .C2(new_n369), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n249), .A2(KEYINPUT4), .A3(G244), .A4(new_n250), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n249), .A2(G250), .A3(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n452), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n254), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n512), .A2(new_n260), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n507), .B1(new_n593), .B2(new_n501), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G200), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n254), .B2(new_n591), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G190), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n585), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n570), .A2(new_n327), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n321), .A2(new_n294), .ZN(new_n603));
  INV_X1    g0403(.A(new_n321), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n467), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n555), .A2(new_n557), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n550), .B2(new_n553), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n603), .B(new_n605), .C1(new_n607), .C2(new_n573), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT81), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n570), .A2(new_n609), .A3(new_n327), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n567), .A2(new_n270), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n602), .A2(new_n608), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n596), .A2(new_n270), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n598), .A2(new_n327), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n403), .A2(G77), .ZN(new_n615));
  INV_X1    g0415(.A(new_n578), .ZN(new_n616));
  XNOR2_X1  g0416(.A(G97), .B(G107), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n575), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n615), .B1(new_n618), .B2(new_n221), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n314), .B1(new_n392), .B2(new_n393), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n276), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n584), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n582), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n613), .A2(new_n614), .A3(new_n623), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n572), .A2(new_n600), .A3(new_n612), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n548), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n448), .A2(new_n497), .A3(new_n626), .ZN(G372));
  OAI21_X1  g0427(.A(new_n424), .B1(new_n327), .B2(new_n415), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n409), .A2(new_n435), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n435), .B1(new_n409), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n433), .A2(new_n434), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n380), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n375), .A2(G169), .ZN(new_n634));
  INV_X1    g0434(.A(new_n382), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n384), .A3(new_n383), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n329), .B1(new_n637), .B2(new_n381), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n631), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n307), .A2(new_n309), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n299), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n608), .A2(new_n601), .A3(new_n611), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n572), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n536), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n600), .A2(new_n624), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n543), .A2(new_n488), .A3(new_n491), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n612), .A2(new_n572), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n649), .B2(new_n624), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n643), .A2(new_n572), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n613), .A2(new_n614), .A3(new_n623), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n648), .A2(new_n643), .A3(new_n650), .A4(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n642), .B1(new_n448), .B2(new_n656), .ZN(G369));
  NAND3_X1  g0457(.A1(new_n265), .A2(new_n221), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n542), .A2(new_n663), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n548), .A2(new_n664), .B1(new_n540), .B2(new_n663), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n469), .A2(new_n663), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT88), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n488), .A2(new_n491), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n497), .B2(new_n667), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n663), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n547), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n540), .A2(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n215), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n553), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n220), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n655), .A2(new_n688), .A3(new_n674), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT26), .B1(new_n644), .B2(new_n624), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n653), .A2(new_n652), .A3(new_n572), .A4(new_n612), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n643), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT91), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT91), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n691), .A2(new_n692), .A3(new_n695), .A4(new_n643), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(new_n648), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n674), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n690), .B1(new_n698), .B2(KEYINPUT29), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n563), .A2(new_n509), .A3(new_n513), .A4(new_n566), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n490), .A3(KEYINPUT30), .A4(new_n598), .ZN(new_n702));
  AOI21_X1  g0502(.A(G179), .B1(new_n505), .B2(new_n507), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n596), .A3(new_n493), .A4(new_n567), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n479), .A2(new_n484), .A3(G179), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n596), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n702), .B(new_n704), .C1(new_n706), .C2(KEYINPUT30), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT31), .B1(new_n707), .B2(new_n663), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT90), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n708), .A2(KEYINPUT90), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n512), .A2(G270), .A3(new_n260), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n507), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n254), .B2(new_n483), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(G179), .A3(new_n505), .A4(new_n570), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n598), .A2(KEYINPUT30), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n493), .A2(new_n567), .A3(new_n327), .A4(new_n516), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(new_n598), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n700), .A2(new_n705), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT30), .B1(new_n719), .B2(new_n598), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT31), .B(new_n663), .C1(new_n718), .C2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n710), .A2(new_n711), .B1(KEYINPUT89), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n707), .A2(new_n663), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n722), .A2(KEYINPUT89), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(new_n709), .ZN(new_n730));
  AND4_X1   g0530(.A1(new_n488), .A2(new_n491), .A3(new_n496), .A4(new_n674), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n541), .A2(new_n625), .A3(new_n731), .A4(new_n546), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n723), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n699), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n687), .B1(new_n736), .B2(G1), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT92), .ZN(G364));
  INV_X1    g0538(.A(new_n671), .ZN(new_n739));
  INV_X1    g0539(.A(G13), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n265), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n682), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G330), .B2(new_n670), .ZN(new_n746));
  INV_X1    g0546(.A(new_n744), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n222), .B1(G20), .B2(new_n270), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n331), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n327), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT98), .Z(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(G20), .A2(G179), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(KEYINPUT95), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT95), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n755), .B2(new_n377), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n754), .A2(new_n453), .B1(new_n343), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n221), .A2(G179), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT97), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT97), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(KEYINPUT32), .A3(new_n397), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT96), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n760), .B2(new_n331), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n757), .A2(KEYINPUT96), .A3(G190), .A4(new_n759), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G50), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT32), .B1(new_n769), .B2(new_n397), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n764), .A2(new_n331), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n314), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n756), .A2(new_n765), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n750), .A2(new_n756), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n249), .B1(new_n780), .B2(new_n202), .C1(new_n237), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n779), .B(new_n782), .C1(G87), .C2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n771), .A2(new_n776), .A3(new_n777), .A4(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n781), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n249), .B1(new_n787), .B2(G322), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(new_n780), .ZN(new_n790));
  INV_X1    g0590(.A(new_n769), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(new_n791), .B2(G329), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n775), .A2(G326), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n498), .A2(new_n499), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n752), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n778), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G303), .B2(new_n784), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n761), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n792), .A2(new_n793), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n749), .B1(new_n786), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n748), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT93), .ZN(new_n807));
  OR2_X1    g0607(.A1(G355), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(G355), .A2(new_n807), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n808), .A2(new_n215), .A3(new_n249), .A4(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(G116), .B2(new_n215), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT94), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n240), .A2(G45), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n681), .A2(new_n249), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n220), .B2(G45), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n812), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n747), .B(new_n802), .C1(new_n806), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n805), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n670), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n746), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n329), .A2(new_n674), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n334), .A2(new_n335), .B1(new_n326), .B2(new_n663), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n329), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n656), .B2(new_n663), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n336), .A2(new_n674), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n648), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n650), .A2(new_n654), .A3(new_n643), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n744), .B1(new_n734), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n734), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n748), .A2(new_n803), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT99), .Z(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n747), .B1(new_n836), .B2(new_n202), .ZN(new_n837));
  INV_X1    g0637(.A(new_n824), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n370), .B1(new_n780), .B2(new_n462), .C1(new_n839), .C2(new_n781), .ZN(new_n840));
  INV_X1    g0640(.A(new_n778), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G87), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n314), .B2(new_n783), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n840), .B(new_n843), .C1(new_n791), .C2(G311), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n453), .B2(new_n754), .C1(new_n796), .C2(new_n762), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G303), .B2(new_n775), .ZN(new_n846));
  INV_X1    g0646(.A(new_n780), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G143), .A2(new_n787), .B1(new_n847), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(new_n775), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n848), .B1(new_n281), .B2(new_n762), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n769), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n370), .B1(new_n784), .B2(G50), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n841), .A2(G68), .ZN(new_n857));
  INV_X1    g0657(.A(new_n752), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n857), .C1(new_n237), .C2(new_n858), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n855), .B(new_n859), .C1(new_n851), .C2(new_n852), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n846), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n837), .B1(new_n804), .B2(new_n838), .C1(new_n861), .C2(new_n749), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n833), .A2(new_n862), .ZN(G384));
  NOR2_X1   g0663(.A1(new_n741), .A2(new_n265), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n697), .A2(new_n674), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n689), .B1(new_n865), .B2(new_n688), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n447), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n642), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT102), .Z(new_n869));
  NAND2_X1  g0669(.A1(new_n830), .A2(new_n822), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT101), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n830), .A2(new_n872), .A3(new_n822), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n661), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n409), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n437), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n427), .A2(new_n431), .A3(new_n876), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n431), .A2(KEYINPUT37), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n409), .B1(new_n628), .B2(new_n875), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n879), .A2(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n878), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n381), .A2(new_n663), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n380), .A2(new_n387), .A3(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n381), .B(new_n663), .C1(new_n637), .C2(new_n379), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n874), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n661), .B1(new_n629), .B2(new_n630), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n886), .A2(KEYINPUT39), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n637), .A2(new_n381), .A3(new_n674), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n876), .B1(new_n632), .B2(new_n631), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n879), .A2(new_n880), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n881), .A2(new_n882), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n897), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n894), .A2(new_n896), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n892), .A2(new_n893), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n869), .B(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n722), .A2(new_n708), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n732), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n824), .B1(new_n889), .B2(new_n890), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(new_n884), .C2(new_n885), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n904), .A2(KEYINPUT40), .A3(new_n912), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n912), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n448), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n447), .A2(new_n916), .A3(new_n912), .A4(new_n917), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(G330), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n864), .B1(new_n910), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n910), .B2(new_n922), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n222), .A2(new_n221), .A3(new_n462), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n579), .B2(KEYINPUT35), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT100), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n927), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT36), .Z(new_n931));
  OAI21_X1  g0731(.A(G77), .B1(new_n237), .B2(new_n343), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n220), .A2(new_n932), .B1(G50), .B2(new_n343), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(G1), .A3(new_n740), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n924), .A2(new_n931), .A3(new_n934), .ZN(G367));
  OAI21_X1  g0735(.A(new_n646), .B1(new_n585), .B2(new_n674), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n653), .A2(new_n663), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n676), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n936), .A2(new_n543), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n663), .B1(new_n942), .B2(new_n624), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n940), .B2(KEYINPUT42), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n559), .A2(new_n569), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n663), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n651), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n643), .B2(new_n946), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n941), .A2(new_n944), .B1(KEYINPUT43), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n949), .B(new_n950), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n672), .A2(new_n938), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n955));
  XNOR2_X1  g0755(.A(new_n682), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT44), .B1(new_n678), .B2(new_n939), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT104), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n678), .A2(KEYINPUT44), .A3(new_n939), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n938), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT45), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n678), .B2(new_n939), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n962), .A2(new_n964), .B1(new_n957), .B2(new_n958), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n672), .ZN(new_n967));
  INV_X1    g0767(.A(new_n664), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n675), .B1(new_n543), .B2(new_n674), .C1(new_n547), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n676), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n739), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n969), .A2(new_n671), .A3(new_n676), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n961), .A2(new_n965), .A3(new_n673), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n967), .A2(new_n736), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n956), .B1(new_n975), .B2(new_n736), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n953), .B(new_n954), .C1(new_n976), .C2(new_n743), .ZN(new_n977));
  INV_X1    g0777(.A(new_n806), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n681), .B2(new_n604), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n234), .A2(new_n814), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n747), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n784), .A2(G116), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT46), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n769), .A2(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n984), .B2(new_n983), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n370), .B1(new_n780), .B2(new_n796), .C1(new_n482), .C2(new_n781), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n858), .A2(new_n314), .B1(new_n778), .B2(new_n453), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n794), .C2(new_n761), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n986), .B(new_n989), .C1(new_n789), .C2(new_n849), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n249), .B1(new_n780), .B2(new_n295), .C1(new_n281), .C2(new_n781), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n237), .A2(new_n783), .B1(new_n778), .B2(new_n202), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n791), .C2(G137), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n753), .A2(G68), .B1(G159), .B2(new_n761), .ZN(new_n994));
  INV_X1    g0794(.A(G143), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n993), .B(new_n994), .C1(new_n995), .C2(new_n849), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n990), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  OAI221_X1 g0798(.A(new_n981), .B1(new_n818), .B2(new_n948), .C1(new_n998), .C2(new_n749), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n977), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT105), .ZN(G387));
  NAND3_X1  g0801(.A1(new_n973), .A2(new_n699), .A3(new_n734), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n682), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT113), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT113), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1005), .A3(new_n682), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n969), .A2(new_n671), .A3(new_n676), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n671), .B1(new_n969), .B2(new_n676), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n735), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT114), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n735), .A2(KEYINPUT114), .A3(new_n1009), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1004), .A2(new_n1006), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1009), .A2(new_n742), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT106), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(KEYINPUT106), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n781), .A2(new_n295), .B1(new_n780), .B2(new_n343), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n754), .A2(new_n321), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n283), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1018), .B(new_n1019), .C1(new_n1020), .C2(new_n761), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n370), .B1(new_n841), .B2(G97), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n202), .B2(new_n783), .C1(new_n769), .C2(new_n281), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT109), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(new_n397), .C2(new_n849), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n784), .A2(new_n794), .B1(new_n752), .B2(G283), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT110), .Z(new_n1027));
  AOI22_X1  g0827(.A1(G317), .A2(new_n787), .B1(new_n847), .B2(G303), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n762), .B2(new_n789), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G322), .B2(new_n775), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1027), .B1(new_n1030), .B2(KEYINPUT48), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT111), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1030), .A2(KEYINPUT48), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT112), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(KEYINPUT112), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n791), .A2(G326), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n249), .B1(new_n841), .B2(G116), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT49), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1025), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n748), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n249), .A2(new_n215), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1044), .A2(new_n684), .B1(G107), .B2(new_n215), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n681), .B(new_n249), .C1(new_n231), .C2(G45), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n684), .B(new_n257), .C1(new_n343), .C2(new_n202), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT107), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT50), .B1(new_n283), .B2(G50), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1045), .B1(new_n1046), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n744), .B1(new_n1054), .B2(new_n978), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT108), .Z(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n665), .B2(new_n805), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1016), .A2(new_n1017), .B1(new_n1043), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1014), .A2(new_n1058), .ZN(G393));
  INV_X1    g0859(.A(new_n974), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n673), .B1(new_n961), .B2(new_n965), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1002), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n975), .A3(new_n682), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n967), .A2(new_n743), .A3(new_n974), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n842), .B(new_n249), .C1(new_n283), .C2(new_n780), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n754), .A2(new_n202), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G50), .C2(new_n761), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n769), .A2(new_n995), .B1(new_n343), .B2(new_n783), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT115), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n775), .A2(G150), .B1(G159), .B2(new_n787), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT51), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1067), .B(new_n1069), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n775), .A2(G317), .B1(G311), .B2(new_n787), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n370), .B1(new_n780), .B2(new_n839), .C1(new_n778), .C2(new_n314), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n858), .A2(new_n462), .B1(new_n783), .B2(new_n796), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n791), .C2(G322), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n482), .B2(new_n762), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1076), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n748), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n978), .B1(G97), .B2(new_n681), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n243), .A2(new_n814), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n747), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1085), .B(new_n1088), .C1(new_n818), .C2(new_n938), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1064), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1063), .A2(new_n1090), .ZN(G390));
  NAND2_X1  g0891(.A1(new_n912), .A2(G330), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n891), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1092), .A2(new_n824), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n822), .ZN(new_n1095));
  AOI211_X1 g0895(.A(KEYINPUT101), .B(new_n1095), .C1(new_n655), .C2(new_n827), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n872), .B1(new_n830), .B2(new_n822), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n891), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1098), .A2(new_n895), .B1(new_n906), .B2(new_n894), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n895), .B(KEYINPUT117), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n904), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n823), .A2(new_n329), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n822), .B1(new_n698), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1101), .B1(new_n1103), .B2(new_n891), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1094), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1101), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1102), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1095), .B1(new_n865), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n1108), .B2(new_n1093), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n733), .A2(G330), .A3(new_n838), .A4(new_n891), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n896), .B1(new_n874), .B2(new_n891), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n894), .A2(new_n906), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1109), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1105), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1092), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n447), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n867), .A2(new_n1116), .A3(new_n642), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1093), .B1(new_n1092), .B2(new_n824), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1110), .A2(new_n1108), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n733), .A2(G330), .A3(new_n838), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1094), .B1(new_n1120), .B2(new_n1093), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n874), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1117), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1114), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1105), .A2(new_n1113), .A3(new_n1117), .A4(new_n1123), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n682), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1105), .A2(new_n1113), .A3(new_n743), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n747), .B1(new_n836), .B2(new_n283), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n775), .A2(G128), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n370), .B1(new_n847), .B2(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n295), .B2(new_n778), .C1(new_n854), .C2(new_n781), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G125), .B2(new_n791), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n783), .A2(new_n281), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n753), .A2(G159), .B1(G137), .B2(new_n761), .ZN(new_n1138));
  AND4_X1   g0938(.A1(new_n1130), .A2(new_n1135), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n249), .B1(new_n787), .B2(G116), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1140), .B(new_n857), .C1(new_n552), .C2(new_n783), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1141), .B(new_n1066), .C1(G294), .C2(new_n791), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n761), .A2(G107), .B1(G97), .B2(new_n847), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n849), .B2(new_n796), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT118), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1139), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1129), .B1(new_n749), .B2(new_n1146), .C1(new_n1112), .C2(new_n804), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1127), .A2(new_n1128), .A3(new_n1147), .ZN(G378));
  NAND2_X1  g0948(.A1(new_n297), .A2(new_n875), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n310), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n310), .A2(new_n1149), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n912), .A2(new_n913), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n885), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n903), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n917), .B(G330), .C1(new_n1159), .C2(KEYINPUT40), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT120), .ZN(new_n1161));
  INV_X1    g0961(.A(G330), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n914), .B2(new_n915), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT120), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n917), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1156), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n1163), .B2(new_n917), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1156), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n908), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  AND4_X1   g0970(.A1(new_n1164), .A2(new_n916), .A3(G330), .A4(new_n917), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1168), .B1(new_n1171), .B2(new_n1167), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n908), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1161), .A2(new_n1156), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1170), .A2(new_n1175), .A3(KEYINPUT121), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT121), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1172), .A2(new_n1173), .A3(new_n1177), .A4(new_n1174), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n743), .A3(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n744), .B1(new_n835), .B2(G50), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n370), .A2(new_n256), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n784), .B2(G77), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n237), .B2(new_n778), .C1(new_n769), .C2(new_n796), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT119), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G107), .A2(new_n787), .B1(new_n847), .B2(new_n604), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n754), .B2(new_n343), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G97), .B2(new_n761), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1184), .B(new_n1187), .C1(new_n462), .C2(new_n849), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G50), .B1(new_n246), .B2(new_n256), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1188), .A2(new_n1189), .B1(new_n1181), .B2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G128), .A2(new_n787), .B1(new_n847), .B2(G137), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n783), .B2(new_n1131), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n753), .B2(G150), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n775), .A2(G125), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n854), .C2(new_n762), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n791), .A2(G124), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n841), .C2(G159), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1191), .B1(new_n1189), .B2(new_n1188), .C1(new_n1197), .C2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1180), .B1(new_n1202), .B2(new_n748), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1156), .B2(new_n804), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1179), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1126), .A2(new_n1117), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1176), .A2(new_n1206), .A3(new_n1178), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT57), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1170), .A2(new_n1175), .A3(KEYINPUT122), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT122), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(new_n908), .C1(new_n1166), .C2(new_n1169), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n1206), .A3(KEYINPUT57), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n682), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1205), .B1(new_n1209), .B2(new_n1214), .ZN(G375));
  NAND2_X1  g1015(.A1(new_n775), .A2(G132), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT124), .Z(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n850), .B2(new_n781), .C1(new_n762), .C2(new_n1131), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT125), .Z(new_n1219));
  AOI21_X1  g1019(.A(new_n370), .B1(new_n847), .B2(G150), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n237), .B2(new_n778), .C1(new_n397), .C2(new_n783), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G128), .B2(new_n791), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1219), .B(new_n1222), .C1(new_n295), .C2(new_n754), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1019), .B1(G116), .B2(new_n761), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n370), .B1(new_n780), .B2(new_n314), .C1(new_n796), .C2(new_n781), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n202), .A2(new_n778), .B1(new_n783), .B2(new_n453), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n791), .C2(G303), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1224), .B(new_n1227), .C1(new_n839), .C2(new_n849), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n749), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n747), .B(new_n1229), .C1(new_n343), .C2(new_n836), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1093), .A2(new_n803), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1230), .A2(new_n1231), .B1(new_n1123), .B2(new_n743), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n956), .B(KEYINPUT123), .Z(new_n1233));
  NAND2_X1  g1033(.A1(new_n1124), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1117), .A2(new_n1123), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1232), .B1(new_n1234), .B2(new_n1235), .ZN(G381));
  NOR3_X1   g1036(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1237));
  INV_X1    g1037(.A(G378), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1014), .A2(new_n1058), .A3(new_n820), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  OR3_X1    g1041(.A1(G387), .A2(G375), .A3(new_n1241), .ZN(G407));
  NAND2_X1  g1042(.A1(new_n1238), .A2(new_n662), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(G375), .C2(new_n1243), .ZN(G409));
  AOI21_X1  g1044(.A(new_n820), .B1(new_n1014), .B2(new_n1058), .ZN(new_n1245));
  OAI21_X1  g1045(.A(G390), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT105), .B1(new_n1247), .B2(new_n1239), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1248), .B2(G390), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1000), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n977), .A2(new_n999), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n1246), .C1(G390), .C2(new_n1248), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G378), .B(new_n1205), .C1(new_n1209), .C2(new_n1214), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1210), .A2(new_n743), .A3(new_n1212), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1233), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1204), .B(new_n1255), .C1(new_n1207), .C2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1238), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1235), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n682), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1235), .B1(KEYINPUT60), .B2(new_n1124), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1232), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n833), .A3(new_n862), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G384), .B(new_n1232), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1254), .A2(KEYINPUT126), .A3(new_n1258), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n662), .A2(G213), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1261), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1259), .A2(new_n1271), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1268), .A2(new_n1273), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1272), .A2(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n662), .A2(G213), .A3(G2897), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1268), .B(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1253), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1272), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1261), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1279), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1268), .A2(new_n1282), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1259), .A2(new_n1271), .A3(new_n1287), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1250), .A2(new_n1252), .A3(new_n1277), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AND4_X1   g1091(.A1(KEYINPUT127), .A2(new_n1283), .A3(new_n1286), .A4(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1290), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT127), .B1(new_n1293), .B2(new_n1283), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1281), .B1(new_n1292), .B2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1238), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1254), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1297), .B(new_n1269), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(new_n1253), .ZN(G402));
endmodule


