//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(KEYINPUT10), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT78), .ZN(new_n188));
  XNOR2_X1  g002(.A(G104), .B(G107), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  OAI211_X1 g009(.A(KEYINPUT78), .B(G101), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n200), .A2(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n204), .B(new_n206), .C1(G128), .C2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n194), .A3(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n192), .A2(G107), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n190), .A4(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n197), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n209), .A2(new_n211), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n195), .A2(G101), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n191), .A2(new_n196), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT79), .B1(new_n219), .B2(new_n208), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n187), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n202), .A2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n225), .A2(new_n205), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n207), .A2(new_n226), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n190), .A2(KEYINPUT4), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n229), .A2(new_n230), .B1(new_n222), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT77), .B1(new_n224), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n224), .A2(KEYINPUT77), .A3(new_n232), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT65), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G134), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n241), .A3(G137), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n238), .A2(G137), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n237), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n241), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT11), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G131), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT65), .B(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n237), .B1(new_n251), .B2(G137), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n243), .B1(new_n251), .B2(G137), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n250), .B(new_n252), .C1(new_n253), .C2(new_n237), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n254), .A3(KEYINPUT66), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(G131), .C1(new_n245), .C2(new_n248), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n219), .A2(KEYINPUT10), .ZN(new_n259));
  AOI21_X1  g073(.A(G128), .B1(new_n201), .B2(new_n203), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n203), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT67), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n206), .B(new_n264), .C1(new_n207), .C2(G128), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n263), .A2(new_n265), .B1(new_n207), .B2(new_n199), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n221), .A2(new_n236), .A3(new_n258), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G227), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT76), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n219), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n266), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n216), .B2(new_n220), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n255), .A2(new_n257), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n276), .A2(KEYINPUT12), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT12), .B1(new_n276), .B2(new_n277), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n268), .B(new_n273), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n224), .A2(KEYINPUT77), .A3(new_n232), .ZN(new_n281));
  OAI22_X1  g095(.A1(new_n281), .A2(new_n233), .B1(new_n266), .B2(new_n259), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n214), .A2(new_n215), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n219), .A2(KEYINPUT79), .A3(new_n208), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT10), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n282), .A2(new_n285), .A3(new_n277), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n277), .B1(new_n282), .B2(new_n285), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT81), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT81), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n289), .B(new_n277), .C1(new_n282), .C2(new_n285), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n280), .B1(new_n291), .B2(new_n273), .ZN(new_n292));
  INV_X1    g106(.A(G469), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT72), .B(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n299));
  INV_X1    g113(.A(new_n273), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n268), .A2(new_n302), .A3(new_n273), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n221), .A2(new_n236), .A3(new_n267), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n289), .B1(new_n304), .B2(new_n277), .ZN(new_n305));
  INV_X1    g119(.A(new_n290), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n302), .B1(new_n268), .B2(new_n273), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n301), .B(G469), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n295), .A2(new_n298), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G210), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G110), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT8), .ZN(new_n317));
  INV_X1    g131(.A(G113), .ZN(new_n318));
  INV_X1    g132(.A(G116), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G119), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G116), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(G119), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT5), .ZN(new_n326));
  XNOR2_X1  g140(.A(G116), .B(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G113), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n322), .A2(new_n326), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n197), .A2(new_n332), .A3(new_n213), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n197), .B2(new_n213), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n317), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT85), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n229), .A2(new_n230), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G125), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n266), .B2(G125), .ZN(new_n340));
  INV_X1    g154(.A(G224), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(G953), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(KEYINPUT7), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n339), .B(new_n345), .C1(new_n266), .C2(G125), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(new_n317), .C1(new_n334), .C2(new_n335), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n337), .A2(new_n344), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n333), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT68), .B1(new_n331), .B2(new_n327), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n324), .A2(new_n325), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT2), .B(G113), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT68), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n222), .A2(new_n231), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n224), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n219), .A2(KEYINPUT83), .A3(new_n332), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n351), .A2(new_n359), .A3(new_n360), .A4(new_n316), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n296), .B1(new_n349), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n340), .B(new_n342), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(KEYINPUT6), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n351), .A2(new_n359), .A3(new_n360), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n316), .A2(KEYINPUT84), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(KEYINPUT6), .A3(new_n367), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n364), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n315), .B1(new_n363), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n340), .B(new_n343), .ZN(new_n373));
  AOI22_X1  g187(.A1(KEYINPUT6), .A2(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n374));
  INV_X1    g188(.A(new_n370), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n344), .A2(new_n346), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(new_n361), .A3(new_n337), .A4(new_n348), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n376), .A2(new_n378), .A3(new_n296), .A4(new_n314), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n372), .A2(KEYINPUT86), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n363), .A2(new_n371), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(new_n314), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G214), .B1(G237), .B2(G902), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n385), .B(KEYINPUT82), .Z(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n313), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n269), .A2(G952), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(G234), .B2(G237), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(KEYINPUT94), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI211_X1 g206(.A(new_n269), .B(new_n294), .C1(G234), .C2(G237), .ZN(new_n393));
  XOR2_X1   g207(.A(new_n393), .B(KEYINPUT95), .Z(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT21), .B(G898), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n319), .A2(KEYINPUT14), .A3(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(G116), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(G107), .B(new_n399), .C1(new_n401), .C2(KEYINPUT14), .ZN(new_n402));
  XNOR2_X1  g216(.A(G128), .B(G143), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n251), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n251), .A2(new_n403), .ZN(new_n405));
  OAI221_X1 g219(.A(new_n402), .B1(G107), .B2(new_n401), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n406), .A2(KEYINPUT93), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n400), .B(G107), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT92), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(KEYINPUT13), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n198), .A2(KEYINPUT13), .A3(G143), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n238), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n404), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n406), .A2(KEYINPUT93), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G217), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n311), .A2(new_n417), .A3(G953), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n418), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n407), .A2(new_n414), .A3(new_n415), .A4(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n294), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n424), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT87), .B(G143), .ZN(new_n430));
  INV_X1    g244(.A(G237), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n269), .A3(G214), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n434), .B2(new_n202), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(KEYINPUT18), .A2(G131), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n429), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT88), .B(new_n437), .C1(new_n433), .C2(new_n435), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n438), .ZN(new_n442));
  XNOR2_X1  g256(.A(G125), .B(G140), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n200), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(KEYINPUT73), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT73), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G125), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n449), .B2(new_n200), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n441), .A2(new_n442), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n436), .A2(new_n250), .ZN(new_n452));
  OAI21_X1  g266(.A(G131), .B1(new_n433), .B2(new_n435), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  MUX2_X1   g268(.A(new_n454), .B(new_n453), .S(KEYINPUT17), .Z(new_n455));
  AOI21_X1  g269(.A(KEYINPUT16), .B1(new_n447), .B2(G125), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT16), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n449), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G146), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n200), .B(new_n457), .C1(new_n449), .C2(new_n458), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(KEYINPUT74), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n463), .A3(G146), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n451), .B1(new_n455), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT89), .B(G104), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n467), .B(new_n468), .Z(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n441), .A2(new_n442), .A3(new_n450), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n443), .A2(KEYINPUT19), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n449), .B2(KEYINPUT19), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n454), .B(new_n460), .C1(G146), .C2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n469), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n475), .B1(new_n466), .B2(new_n469), .ZN(new_n481));
  INV_X1    g295(.A(new_n479), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT20), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n466), .A2(new_n469), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n466), .A2(new_n469), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n296), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT90), .B(G475), .Z(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n484), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n485), .B1(new_n484), .B2(new_n490), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n398), .B(new_n428), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n388), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n338), .A2(KEYINPUT64), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n338), .A2(KEYINPUT64), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n255), .A2(new_n257), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n251), .A2(G137), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n247), .A2(G134), .ZN(new_n499));
  OAI21_X1  g313(.A(G131), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n254), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n501), .A2(new_n266), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n255), .A2(new_n257), .A3(new_n338), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT30), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n505), .A2(new_n357), .A3(new_n356), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n356), .A2(new_n357), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT69), .Z(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n506), .A3(new_n502), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n513));
  NAND3_X1  g327(.A1(new_n431), .A2(new_n269), .A3(G210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT29), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n511), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n509), .B1(new_n497), .B2(new_n502), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT28), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n517), .B(KEYINPUT71), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n518), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n294), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n502), .A2(new_n506), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n509), .B(KEYINPUT69), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n511), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT28), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n523), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n517), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n536), .A2(KEYINPUT29), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n528), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G472), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n508), .A2(new_n511), .A3(new_n536), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n508), .A2(KEYINPUT31), .A3(new_n511), .A4(new_n536), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n524), .A2(new_n526), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n544), .A2(new_n545), .B1(new_n524), .B2(new_n526), .ZN(new_n551));
  INV_X1    g365(.A(new_n549), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n551), .A2(KEYINPUT32), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n540), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n323), .B2(G128), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n556), .B(new_n557), .C1(G119), .C2(new_n198), .ZN(new_n558));
  XNOR2_X1  g372(.A(G119), .B(G128), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  AOI22_X1  g374(.A1(new_n558), .A2(G110), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n462), .A2(new_n464), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n559), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n558), .A2(G110), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(KEYINPUT75), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(KEYINPUT75), .B2(new_n564), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n460), .A3(new_n444), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT22), .B(G137), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n569), .B(new_n570), .Z(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n562), .A2(new_n567), .A3(new_n571), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n294), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n417), .B1(new_n294), .B2(G234), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(G902), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n573), .A2(new_n574), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n577), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n554), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n494), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n190), .ZN(G3));
  NAND2_X1  g398(.A1(new_n548), .A2(new_n549), .ZN(new_n585));
  OAI21_X1  g399(.A(G472), .B1(new_n551), .B2(new_n528), .ZN(new_n586));
  AND4_X1   g400(.A1(new_n585), .A2(new_n313), .A3(new_n581), .A4(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT96), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n484), .A2(new_n490), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT91), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n484), .A2(new_n490), .A3(new_n485), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n419), .A2(new_n592), .A3(new_n421), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n407), .A2(new_n414), .A3(KEYINPUT98), .A4(new_n415), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n418), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT98), .B1(new_n420), .B2(KEYINPUT99), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n416), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT33), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n528), .A2(new_n423), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n595), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT100), .B(G478), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n422), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n590), .A2(new_n591), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n386), .B1(new_n372), .B2(new_n379), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n398), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n588), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND3_X1  g427(.A1(new_n484), .A2(new_n490), .A3(new_n427), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n609), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n588), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NAND2_X1  g432(.A1(new_n586), .A2(new_n585), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n388), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n577), .A2(new_n578), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n572), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n568), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n579), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n493), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT101), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n627), .B(new_n629), .ZN(G12));
  INV_X1    g444(.A(new_n608), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n554), .A2(new_n313), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n392), .B1(new_n395), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n614), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  NAND3_X1  g452(.A1(new_n590), .A2(new_n427), .A3(new_n591), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n621), .A2(new_n624), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n639), .A2(new_n386), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT102), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n384), .B(KEYINPUT38), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n635), .B(KEYINPUT39), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n313), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n645), .B2(KEYINPUT40), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(KEYINPUT40), .B2(new_n645), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n550), .A2(new_n553), .ZN(new_n648));
  INV_X1    g462(.A(new_n512), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n649), .A2(new_n536), .B1(new_n526), .B2(new_n532), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n650), .B2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n642), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n202), .ZN(G45));
  INV_X1    g469(.A(new_n635), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n590), .A2(new_n591), .A3(new_n606), .A4(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n633), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  INV_X1    g474(.A(new_n582), .ZN(new_n661));
  INV_X1    g475(.A(new_n292), .ZN(new_n662));
  OAI21_X1  g476(.A(G469), .B1(new_n662), .B2(new_n528), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n312), .A3(new_n295), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n661), .A2(new_n610), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NAND3_X1  g482(.A1(new_n661), .A2(new_n615), .A3(new_n665), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G116), .ZN(G18));
  NOR4_X1   g484(.A1(new_n493), .A2(new_n631), .A3(new_n625), .A4(new_n664), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n554), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G119), .ZN(G21));
  NOR3_X1   g487(.A1(new_n639), .A2(new_n609), .A3(new_n664), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n525), .B1(new_n534), .B2(KEYINPUT103), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(KEYINPUT103), .B2(new_n534), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n546), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n549), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n678), .A2(new_n581), .A3(new_n586), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G122), .ZN(G24));
  NAND3_X1  g495(.A1(new_n678), .A2(new_n586), .A3(new_n640), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n657), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n664), .A2(new_n631), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G125), .ZN(G27));
  INV_X1    g500(.A(new_n386), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n384), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT105), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n384), .A2(new_n690), .A3(new_n687), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n309), .A2(new_n298), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT104), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n295), .A2(new_n696), .A3(new_n298), .A4(new_n309), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n312), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT106), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n690), .B1(new_n384), .B2(new_n687), .ZN(new_n700));
  AOI211_X1 g514(.A(KEYINPUT105), .B(new_n386), .C1(new_n380), .C2(new_n383), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  INV_X1    g517(.A(new_n312), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n310), .B2(KEYINPUT104), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n702), .A2(new_n703), .A3(new_n697), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n661), .A3(new_n658), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n711), .A2(new_n707), .A3(new_n661), .A4(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n582), .B1(new_n699), .B2(new_n706), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n711), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n710), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  NAND3_X1  g531(.A1(new_n707), .A2(new_n661), .A3(new_n636), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G134), .ZN(G36));
  NOR2_X1   g533(.A1(new_n491), .A2(new_n492), .ZN(new_n720));
  INV_X1    g534(.A(new_n606), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n723), .A2(KEYINPUT109), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(KEYINPUT109), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n722), .B2(new_n725), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n619), .A3(new_n640), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT44), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n301), .B1(new_n307), .B2(new_n308), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n293), .B1(new_n730), .B2(new_n731), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n297), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n295), .B1(new_n734), .B2(KEYINPUT46), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n312), .B(new_n644), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n729), .A2(new_n702), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G137), .ZN(G39));
  NOR4_X1   g554(.A1(new_n554), .A2(new_n692), .A3(new_n657), .A4(new_n581), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n312), .B1(new_n735), .B2(new_n736), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n742), .A2(new_n744), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n741), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G140), .ZN(G42));
  AND4_X1   g563(.A1(new_n581), .A2(new_n722), .A3(new_n312), .A4(new_n687), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n663), .A2(new_n295), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT49), .Z(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(new_n643), .A3(new_n653), .A4(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n727), .A2(new_n392), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n679), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n643), .A2(new_n665), .A3(new_n386), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT116), .ZN(new_n760));
  NOR2_X1   g574(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n755), .A2(new_n758), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n764));
  OAI211_X1 g578(.A(KEYINPUT117), .B(KEYINPUT50), .C1(new_n755), .C2(new_n760), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n765), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT118), .B1(new_n767), .B2(new_n762), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n754), .A2(new_n679), .A3(new_n702), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT115), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n746), .A2(new_n747), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n312), .B2(new_n751), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n692), .A2(new_n664), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n754), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n682), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n581), .A2(new_n653), .A3(new_n392), .A4(new_n774), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n720), .A2(new_n606), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n766), .A2(new_n768), .A3(new_n773), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n773), .A2(new_n779), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n767), .A2(new_n762), .A3(new_n781), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n775), .A2(new_n582), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT48), .Z(new_n787));
  AND3_X1   g601(.A1(new_n777), .A2(new_n720), .A3(new_n606), .ZN(new_n788));
  INV_X1    g602(.A(new_n755), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n389), .B(new_n788), .C1(new_n789), .C2(new_n684), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n782), .A2(new_n785), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  INV_X1    g606(.A(new_n583), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n671), .A2(new_n554), .B1(new_n620), .B2(new_n626), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n491), .A2(new_n606), .A3(new_n492), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n427), .B1(new_n590), .B2(new_n591), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n387), .A2(new_n398), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n798), .A2(new_n587), .B1(new_n679), .B2(new_n674), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n661), .B(new_n665), .C1(new_n610), .C2(new_n615), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n793), .A2(new_n794), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n716), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n428), .A2(new_n484), .A3(new_n490), .A4(new_n656), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n625), .A2(new_n803), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n554), .A2(new_n313), .A3(new_n804), .A4(new_n702), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n707), .B2(new_n683), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n806), .A2(new_n807), .A3(new_n718), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n807), .B1(new_n806), .B2(new_n718), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n792), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n793), .A2(new_n794), .A3(new_n799), .A4(new_n800), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n707), .A2(new_n712), .A3(new_n661), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT108), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n714), .A2(new_n711), .A3(new_n712), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n812), .B1(new_n816), .B2(new_n710), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n806), .A2(new_n718), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT111), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n806), .A2(new_n807), .A3(new_n718), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n817), .A2(KEYINPUT112), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n633), .A2(new_n636), .B1(new_n683), .B2(new_n684), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n590), .A2(new_n427), .A3(new_n591), .A4(new_n608), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n698), .A2(new_n825), .A3(new_n640), .A4(new_n635), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n652), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n659), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n824), .A2(new_n827), .A3(new_n830), .A4(new_n659), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n823), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n637), .A2(new_n685), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n835), .B2(KEYINPUT52), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n832), .B(new_n836), .C1(new_n811), .C2(new_n822), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT54), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n716), .B(new_n801), .C1(new_n808), .C2(new_n809), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n835), .B2(KEYINPUT52), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n829), .A2(new_n831), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT113), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n829), .A2(new_n831), .A3(new_n841), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n817), .A3(new_n845), .A4(new_n821), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n832), .B1(new_n811), .B2(new_n822), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n838), .A2(KEYINPUT114), .A3(new_n850), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n850), .A2(KEYINPUT114), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n791), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(G952), .A2(G953), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT119), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n753), .B1(new_n853), .B2(new_n855), .ZN(G75));
  NOR2_X1   g670(.A1(new_n269), .A2(G952), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n843), .A2(new_n846), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n528), .B(new_n315), .C1(new_n834), .C2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n374), .A2(new_n375), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n364), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n376), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT55), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n858), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n866), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n862), .A2(KEYINPUT120), .A3(new_n866), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(G51));
  XNOR2_X1  g686(.A(new_n297), .B(KEYINPUT57), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n839), .A2(new_n792), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT112), .B1(new_n817), .B2(new_n821), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n833), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n840), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n848), .B1(new_n877), .B2(new_n847), .ZN(new_n878));
  INV_X1    g692(.A(new_n850), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n292), .B(KEYINPUT121), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n294), .B1(new_n877), .B2(new_n847), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n732), .A3(new_n733), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n857), .B1(new_n882), .B2(new_n884), .ZN(G54));
  AND2_X1   g699(.A1(KEYINPUT58), .A2(G475), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n857), .B1(new_n887), .B2(new_n481), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n883), .A2(KEYINPUT122), .A3(new_n477), .A4(new_n886), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n883), .A2(new_n477), .A3(new_n886), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(G60));
  AND2_X1   g707(.A1(new_n595), .A2(new_n601), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(G478), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT59), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n878), .B2(new_n879), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n858), .ZN(new_n900));
  INV_X1    g714(.A(new_n897), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n851), .A2(new_n852), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n895), .B2(new_n902), .ZN(G63));
  XNOR2_X1  g717(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n417), .A2(new_n296), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n623), .B(new_n906), .C1(new_n834), .C2(new_n859), .ZN(new_n907));
  INV_X1    g721(.A(new_n906), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n877), .B2(new_n847), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n858), .B(new_n907), .C1(new_n909), .C2(new_n580), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(G66));
  OAI21_X1  g726(.A(G953), .B1(new_n396), .B2(new_n341), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n801), .B2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n863), .B1(G898), .B2(new_n269), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G69));
  NAND2_X1  g730(.A1(new_n505), .A2(new_n507), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT124), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n473), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n824), .A2(new_n659), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT62), .B1(new_n654), .B2(new_n920), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n645), .A2(new_n795), .A3(new_n796), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n661), .A3(new_n702), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n739), .A2(new_n748), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n654), .A2(KEYINPUT62), .A3(new_n920), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n919), .B1(new_n926), .B2(G953), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT125), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n919), .C1(new_n926), .C2(G953), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n737), .A2(new_n582), .A3(new_n825), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n931), .B(new_n920), .C1(new_n636), .C2(new_n714), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n716), .A2(new_n739), .A3(new_n748), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n269), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n919), .B1(G900), .B2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n928), .A2(new_n930), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G72));
  NOR2_X1   g753(.A1(new_n649), .A2(new_n517), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n924), .A2(new_n925), .A3(new_n812), .ZN(new_n941));
  NAND2_X1  g755(.A1(G472), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT63), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n933), .B2(new_n801), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n512), .A2(new_n536), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT126), .Z(new_n947));
  OAI211_X1 g761(.A(new_n944), .B(new_n858), .C1(new_n945), .C2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n877), .B1(new_n876), .B2(new_n836), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n940), .A2(new_n946), .A3(new_n943), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(G57));
endmodule


