//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI211_X1 g034(.A(G137), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT70), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  NAND4_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G137), .A4(new_n457), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n457), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n461), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g052(.A(KEYINPUT69), .B(G2105), .C1(new_n470), .C2(new_n474), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n468), .B1(new_n477), .B2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n458), .A2(new_n459), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n457), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  MUX2_X1   g059(.A(G100), .B(G112), .S(G2105), .Z(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2104), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n457), .A2(G102), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2105), .ZN(new_n492));
  AOI211_X1 g067(.A(KEYINPUT71), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  INV_X1    g069(.A(G102), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n492), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n494), .B1(new_n496), .B2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n489), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .A4(new_n457), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT72), .Z(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n508), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n514), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n518), .A2(new_n519), .B1(new_n505), .B2(new_n506), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n516), .A2(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n511), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  OAI211_X1 g100(.A(G51), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(G89), .B1(new_n505), .B2(new_n506), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(new_n529), .B1(new_n513), .B2(new_n514), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G168));
  OR2_X1    g106(.A1(new_n505), .A2(new_n506), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n520), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n533), .A2(new_n540), .B1(new_n541), .B2(new_n520), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n517), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  INV_X1    g128(.A(G91), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n520), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n532), .A2(KEYINPUT75), .A3(G91), .A4(new_n515), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(KEYINPUT74), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n559), .B(G543), .C1(new_n506), .C2(new_n505), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n557), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n563), .B2(new_n517), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  OR2_X1    g143(.A1(new_n511), .A2(new_n522), .ZN(G303));
  INV_X1    g144(.A(new_n520), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n570), .A2(new_n571), .A3(G87), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n571), .B1(new_n570), .B2(G87), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n515), .A2(G74), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(new_n509), .B2(G49), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n570), .A2(G86), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n513), .B2(new_n514), .ZN(new_n580));
  AND2_X1   g155(.A1(G73), .A2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n509), .A2(G48), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(G305));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n533), .A2(new_n585), .B1(new_n586), .B2(new_n520), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n517), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT77), .B(G66), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n515), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g170(.A1(G79), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n515), .B2(new_n594), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n517), .B1(new_n598), .B2(KEYINPUT78), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n520), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n532), .A2(KEYINPUT10), .A3(G92), .A4(new_n515), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n603), .A2(new_n604), .B1(G54), .B2(new_n509), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT79), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n592), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n592), .B1(new_n607), .B2(G868), .ZN(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g185(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g186(.A(KEYINPUT80), .B(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(G860), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT81), .Z(G148));
  NAND2_X1  g189(.A1(new_n607), .A2(new_n612), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT82), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n481), .A2(G2104), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT13), .Z(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n481), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n483), .A2(G123), .ZN(new_n628));
  AND2_X1   g203(.A1(G111), .A2(G2105), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G99), .B2(new_n457), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n490), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(new_n626), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  INV_X1    g210(.A(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2427), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2427), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G2430), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n638), .A2(new_n639), .A3(G2430), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .A4(new_n649), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g232(.A1(new_n651), .A2(KEYINPUT84), .A3(new_n652), .A4(new_n654), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(G14), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n651), .A2(new_n652), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n661), .B2(new_n653), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n667), .B(KEYINPUT17), .Z(new_n670));
  INV_X1    g245(.A(new_n666), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n671), .A2(new_n665), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n669), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n666), .A2(new_n667), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n674), .A2(KEYINPUT85), .A3(new_n665), .ZN(new_n675));
  OAI21_X1  g250(.A(KEYINPUT85), .B1(new_n674), .B2(new_n665), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n671), .C2(new_n670), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n632), .A3(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n632), .B1(new_n673), .B2(new_n677), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n624), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n682), .A2(G2100), .A3(new_n678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT90), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT87), .Z(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n687), .B(KEYINPUT87), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT88), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT20), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n694), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n695), .A2(new_n696), .ZN(new_n704));
  AND4_X1   g279(.A1(new_n693), .A2(new_n691), .A3(new_n697), .A4(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n691), .B2(new_n693), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n708));
  AND3_X1   g283(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n703), .B2(new_n707), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n686), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n703), .A2(new_n707), .ZN(new_n712));
  INV_X1    g287(.A(new_n708), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n686), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1981), .B(G1986), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT89), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n711), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n711), .B2(new_n717), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(G229));
  NOR2_X1   g298(.A1(G16), .A2(G24), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n590), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1986), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G22), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT94), .Z(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G303), .B2(G16), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT95), .B(G1971), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G23), .ZN(new_n733));
  INV_X1    g308(.A(G288), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT33), .B(G1976), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT93), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n735), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G6), .A2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G305), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G16), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT32), .B(G1981), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n732), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n726), .B1(new_n744), .B2(KEYINPUT34), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G25), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n481), .A2(G131), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n483), .A2(G119), .ZN(new_n749));
  MUX2_X1   g324(.A(G95), .B(G107), .S(G2105), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2104), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT91), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT91), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n748), .A2(new_n749), .A3(new_n754), .A4(new_n751), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT92), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n747), .B1(new_n758), .B2(new_n746), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n745), .B(new_n761), .C1(KEYINPUT34), .C2(new_n744), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT36), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n727), .A2(G4), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n607), .B2(new_n727), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G35), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G162), .B2(G29), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT29), .Z(new_n770));
  INV_X1    g345(.A(G2090), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT102), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n727), .A2(G20), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT23), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n565), .B2(new_n727), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n773), .B2(KEYINPUT102), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n746), .A2(G33), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n481), .A2(G139), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT96), .B(KEYINPUT25), .ZN(new_n782));
  INV_X1    g357(.A(G103), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n782), .A2(new_n783), .A3(new_n465), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n782), .B1(new_n783), .B2(new_n465), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n462), .A2(G127), .ZN(new_n788));
  AND2_X1   g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n787), .B1(G2105), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n780), .B1(new_n791), .B2(new_n746), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G2072), .Z(new_n793));
  AND4_X1   g368(.A1(new_n767), .A2(new_n774), .A3(new_n779), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G27), .A2(G29), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G164), .B2(G29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2078), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n770), .A2(new_n771), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(new_n746), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G160), .B2(new_n746), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n797), .B(new_n798), .C1(G2084), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n631), .A2(new_n746), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT101), .Z(new_n805));
  INV_X1    g380(.A(G1961), .ZN(new_n806));
  NOR2_X1   g381(.A1(G171), .A2(new_n727), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G5), .B2(new_n727), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n727), .A2(G21), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G168), .B2(new_n727), .ZN(new_n811));
  INV_X1    g386(.A(G1966), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n809), .B(new_n813), .C1(G2084), .C2(new_n802), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n746), .A2(G26), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT28), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n481), .A2(G140), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n483), .A2(G128), .ZN(new_n818));
  MUX2_X1   g393(.A(G104), .B(G116), .S(G2105), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G2104), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n816), .B1(new_n822), .B2(new_n746), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2067), .ZN(new_n824));
  NOR2_X1   g399(.A1(G16), .A2(G19), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n545), .B2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1341), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT31), .B(G11), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT30), .B(G28), .Z(new_n829));
  OAI221_X1 g404(.A(new_n828), .B1(G29), .B2(new_n829), .C1(new_n808), .C2(new_n806), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n814), .A2(new_n824), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n746), .A2(G32), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n833));
  NAND3_X1  g408(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT99), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT26), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n483), .A2(G129), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n481), .A2(G141), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n466), .A2(G105), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n833), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n837), .A2(new_n841), .A3(new_n833), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n832), .B1(new_n845), .B2(new_n746), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT27), .B(G1996), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n794), .A2(new_n803), .A3(new_n831), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n763), .A2(new_n849), .ZN(G311));
  INV_X1    g425(.A(G311), .ZN(G150));
  AOI22_X1  g426(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n517), .ZN(new_n853));
  OAI211_X1 g428(.A(G55), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n520), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G860), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n545), .A2(new_n857), .ZN(new_n861));
  OAI22_X1  g436(.A1(new_n542), .A2(new_n544), .B1(new_n853), .B2(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n607), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n858), .B1(new_n867), .B2(KEYINPUT39), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n860), .B1(new_n868), .B2(new_n869), .ZN(G145));
  INV_X1    g445(.A(new_n844), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n822), .A3(new_n842), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n821), .B1(new_n843), .B2(new_n844), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n622), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n756), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n462), .A2(new_n457), .ZN(new_n877));
  INV_X1    g452(.A(G142), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  OAI22_X1  g455(.A1(new_n879), .A2(new_n880), .B1(G118), .B2(new_n457), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  OAI22_X1  g457(.A1(new_n877), .A2(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n483), .A2(G130), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n622), .A2(new_n753), .A3(new_n755), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n876), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n876), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n874), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n889), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n622), .B1(new_n753), .B2(new_n755), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n896), .A2(new_n890), .A3(new_n873), .A4(new_n872), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n791), .B(G164), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G160), .B(new_n487), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n631), .B(KEYINPUT103), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n791), .B(G164), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n897), .A3(new_n893), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n900), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n900), .B2(new_n905), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n906), .A2(new_n907), .A3(G37), .ZN(new_n908));
  XNOR2_X1  g483(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(G395));
  NOR3_X1   g485(.A1(new_n853), .A2(new_n856), .A3(G868), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(new_n740), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n734), .A2(new_n590), .ZN(new_n913));
  NAND2_X1  g488(.A1(G288), .A2(G290), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n912), .B(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n606), .A2(new_n565), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n600), .B(new_n605), .C1(new_n561), .C2(new_n564), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n606), .A2(new_n565), .A3(KEYINPUT107), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n921), .A2(new_n925), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n863), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n616), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n616), .A2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n616), .A2(new_n931), .ZN(new_n935));
  INV_X1    g510(.A(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n616), .A2(new_n931), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n920), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(new_n938), .A3(new_n920), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n940), .A2(KEYINPUT108), .A3(KEYINPUT42), .A4(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n943), .A2(new_n939), .B1(new_n917), .B2(new_n918), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n911), .B1(new_n945), .B2(G868), .ZN(G295));
  AOI21_X1  g521(.A(new_n911), .B1(new_n945), .B2(G868), .ZN(G331));
  INV_X1    g522(.A(new_n915), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(new_n912), .ZN(new_n949));
  OAI21_X1  g524(.A(G286), .B1(new_n538), .B2(new_n536), .ZN(new_n950));
  NAND2_X1  g525(.A1(G171), .A2(G168), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n863), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n950), .A2(new_n861), .A3(new_n951), .A4(new_n862), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n927), .A2(new_n955), .A3(new_n929), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n928), .A3(new_n954), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n949), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(G37), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n925), .A4(new_n926), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(KEYINPUT111), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(KEYINPUT111), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n964), .A2(new_n955), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n936), .B1(new_n955), .B2(KEYINPUT41), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n949), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT43), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n958), .A2(KEYINPUT109), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n956), .A2(new_n971), .A3(new_n957), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n916), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n969), .B1(new_n973), .B2(G37), .ZN(new_n974));
  INV_X1    g549(.A(new_n972), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n971), .B1(new_n956), .B2(new_n957), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n949), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G37), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(KEYINPUT110), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n959), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n968), .B1(new_n980), .B2(KEYINPUT43), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(KEYINPUT44), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n960), .ZN(new_n986));
  INV_X1    g561(.A(new_n967), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT43), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n983), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n982), .A2(new_n989), .ZN(G397));
  INV_X1    g565(.A(G2084), .ZN(new_n991));
  AND2_X1   g566(.A1(G160), .A2(G40), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n498), .B2(new_n503), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(KEYINPUT114), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(new_n993), .C1(new_n498), .C2(new_n503), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT50), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n991), .B(new_n992), .C1(new_n997), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n998), .B2(new_n1000), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  OAI211_X1 g579(.A(G160), .B(G40), .C1(new_n1004), .C2(new_n994), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n812), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT51), .B(G8), .C1(new_n1007), .C2(G286), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT124), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT124), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G168), .A2(new_n1011), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1010), .B(KEYINPUT51), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1012), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1013), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1009), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT123), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1015), .B2(G168), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1012), .A2(KEYINPUT123), .A3(G286), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n992), .B1(new_n997), .B2(new_n1001), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n994), .A2(new_n1004), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1005), .A2(new_n1028), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1026), .A2(G2090), .B1(G1971), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(G8), .B1(new_n511), .B2(new_n522), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n998), .A2(G40), .A3(G160), .A4(new_n1000), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n574), .A2(G1976), .A3(new_n576), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G305), .A2(G1981), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n578), .A2(new_n583), .A3(new_n1040), .A4(new_n582), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1039), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT49), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(G8), .A3(new_n1035), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT115), .B(G1976), .Z(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1047), .A2(G8), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1038), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1031), .B(KEYINPUT55), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n998), .B2(new_n1000), .ZN(new_n1053));
  OAI211_X1 g628(.A(G160), .B(G40), .C1(KEYINPUT50), .C2(new_n994), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n995), .A2(KEYINPUT45), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n992), .A2(new_n1056), .A3(new_n1027), .ZN(new_n1057));
  INV_X1    g632(.A(G1971), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1055), .A2(new_n771), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1051), .B1(new_n1059), .B2(new_n1011), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1034), .A2(new_n1050), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT125), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1034), .A2(new_n1050), .A3(new_n1060), .A4(KEYINPUT125), .ZN(new_n1064));
  INV_X1    g639(.A(G2078), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n1029), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1065), .A2(KEYINPUT53), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1026), .A2(new_n806), .ZN(new_n1070));
  AOI21_X1  g645(.A(G301), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1063), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1019), .A2(new_n1073), .A3(new_n1023), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1025), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n1076), .B(KEYINPUT116), .Z(new_n1077));
  AOI22_X1  g652(.A1(new_n1077), .A2(new_n1045), .B1(new_n1040), .B2(new_n740), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1035), .A2(G8), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1078), .A2(new_n1079), .B1(new_n1034), .B2(new_n1049), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1033), .B1(new_n1030), .B2(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1012), .A2(G168), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n1034), .A3(new_n1050), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1061), .B2(new_n1082), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1080), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1956), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1089));
  AND2_X1   g664(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1090));
  NOR2_X1   g665(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n565), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n565), .A2(new_n1091), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT56), .B(G2072), .Z(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n992), .A2(new_n1056), .A3(new_n1027), .A4(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1089), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1035), .A2(G2067), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1026), .B2(new_n766), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1100), .A2(new_n606), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1094), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1098), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT58), .B(G1341), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT118), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1035), .A2(KEYINPUT119), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1996), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n992), .A2(new_n1109), .A3(new_n1056), .A4(new_n1027), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT119), .B1(new_n1035), .B2(new_n1107), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT120), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1035), .A2(new_n1107), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1105), .B1(new_n1119), .B2(new_n545), .ZN(new_n1120));
  INV_X1    g695(.A(new_n545), .ZN(new_n1121));
  AOI211_X1 g696(.A(KEYINPUT59), .B(new_n1121), .C1(new_n1113), .C2(new_n1118), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT121), .B(new_n1124), .C1(new_n1098), .C2(new_n1102), .ZN(new_n1128));
  OR3_X1    g703(.A1(new_n1098), .A2(new_n1102), .A3(new_n1124), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1123), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1100), .A2(KEYINPUT60), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(new_n606), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1136), .A2(new_n1137), .B1(KEYINPUT60), .B2(new_n1100), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1104), .B1(new_n1131), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(G171), .B(KEYINPUT54), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1140), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1068), .A2(G40), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n475), .A2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n468), .B(new_n1144), .C1(new_n995), .C2(KEYINPUT45), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1142), .B(new_n1066), .C1(new_n1027), .C2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1070), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1024), .A2(new_n1063), .A3(new_n1064), .A4(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1075), .B(new_n1087), .C1(new_n1139), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n992), .A2(new_n1028), .ZN(new_n1150));
  OR3_X1    g725(.A1(new_n1150), .A2(KEYINPUT112), .A3(G1996), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT112), .B1(new_n1150), .B2(G1996), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n845), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1154), .A2(KEYINPUT113), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(KEYINPUT113), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1150), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n821), .A2(G2067), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n821), .A2(G2067), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n845), .B2(new_n1109), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1155), .A2(new_n1156), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n756), .B(new_n760), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1150), .B2(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(G290), .A2(G1986), .ZN(new_n1165));
  NAND2_X1  g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1150), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1149), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1150), .B1(new_n845), .B2(new_n1160), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1153), .B2(KEYINPUT46), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(KEYINPUT46), .B2(new_n1153), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT47), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1150), .A2(new_n1165), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT48), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1173), .B1(new_n1164), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1162), .A2(new_n758), .A3(new_n760), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1150), .B1(new_n1177), .B2(new_n1158), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1169), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1182));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n681), .A2(new_n683), .A3(G319), .ZN(new_n1184));
  INV_X1    g758(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n663), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g760(.A(KEYINPUT126), .B(new_n1184), .C1(new_n659), .C2(new_n662), .ZN(new_n1187));
  OAI21_X1  g761(.A(new_n722), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g762(.A1(new_n1188), .A2(new_n908), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1182), .B1(new_n981), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g764(.A(new_n968), .ZN(new_n1191));
  INV_X1    g765(.A(new_n959), .ZN(new_n1192));
  NOR3_X1   g766(.A1(new_n973), .A2(new_n969), .A3(G37), .ZN(new_n1193));
  AOI21_X1  g767(.A(KEYINPUT110), .B1(new_n977), .B2(new_n978), .ZN(new_n1194));
  OAI211_X1 g768(.A(KEYINPUT43), .B(new_n1192), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  AND4_X1   g769(.A1(new_n1182), .A2(new_n1189), .A3(new_n1191), .A4(new_n1195), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1190), .A2(new_n1196), .ZN(G308));
  NAND2_X1  g771(.A1(new_n981), .A2(new_n1189), .ZN(G225));
endmodule


