//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(KEYINPUT74), .A3(KEYINPUT2), .ZN(new_n206));
  AND2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n203), .A2(KEYINPUT75), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT75), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n202), .A2(new_n215), .A3(KEYINPUT2), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n214), .A2(new_n209), .A3(new_n211), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219));
  XOR2_X1   g018(.A(G211gat), .B(G218gat), .Z(new_n220));
  XOR2_X1   g019(.A(G197gat), .B(G204gat), .Z(new_n221));
  AOI21_X1  g020(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G211gat), .B(G218gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(G197gat), .B(G204gat), .ZN(new_n225));
  INV_X1    g024(.A(G211gat), .ZN(new_n226));
  INV_X1    g025(.A(G218gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n224), .B(new_n225), .C1(KEYINPUT22), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT29), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n219), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI211_X1 g031(.A(KEYINPUT79), .B(KEYINPUT29), .C1(new_n223), .C2(new_n229), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n218), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT80), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n218), .C1(new_n232), .C2(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n223), .A2(new_n229), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n213), .A2(new_n219), .A3(new_n217), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G228gat), .ZN(new_n244));
  INV_X1    g043(.A(G233gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G22gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n218), .B2(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n218), .A2(new_n230), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT81), .B1(new_n239), .B2(new_n240), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(new_n238), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT81), .A3(new_n240), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n249), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n241), .B1(new_n234), .B2(KEYINPUT80), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n246), .B1(new_n259), .B2(new_n237), .ZN(new_n260));
  OAI21_X1  g059(.A(G22gat), .B1(new_n260), .B2(new_n256), .ZN(new_n261));
  INV_X1    g060(.A(G78gat), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n258), .B2(new_n261), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT31), .B(G50gat), .ZN(new_n265));
  INV_X1    g064(.A(G106gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n263), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n249), .B1(new_n248), .B2(new_n257), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n260), .A2(G22gat), .A3(new_n256), .ZN(new_n271));
  OAI21_X1  g070(.A(G78gat), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n267), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G141gat), .B(G148gat), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT74), .B1(new_n202), .B2(KEYINPUT2), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n211), .B1(new_n278), .B2(new_n206), .ZN(new_n279));
  INV_X1    g078(.A(new_n217), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n282), .A2(KEYINPUT68), .B1(G127gat), .B2(G134gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(G127gat), .B2(G134gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(G113gat), .B2(G120gat), .ZN(new_n285));
  AND2_X1   g084(.A1(G113gat), .A2(G120gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OAI221_X1 g087(.A(new_n283), .B1(G127gat), .B2(G134gat), .C1(new_n285), .C2(new_n286), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n281), .A2(new_n290), .A3(new_n239), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n213), .A2(new_n217), .A3(new_n288), .A4(new_n289), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n290), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n295), .A2(KEYINPUT4), .A3(new_n213), .A4(new_n217), .ZN(new_n296));
  NAND2_X1  g095(.A1(G225gat), .A2(G233gat), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n291), .A2(new_n294), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT5), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n290), .B1(new_n279), .B2(new_n280), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n292), .ZN(new_n304));
  INV_X1    g103(.A(new_n297), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n218), .A2(KEYINPUT76), .A3(new_n290), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(KEYINPUT5), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(KEYINPUT5), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n298), .A3(new_n300), .ZN(new_n310));
  XNOR2_X1  g109(.A(G1gat), .B(G29gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT0), .ZN(new_n312));
  XNOR2_X1  g111(.A(G57gat), .B(G85gat), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n312), .B(new_n313), .Z(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n308), .A2(new_n310), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT85), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT85), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n308), .A2(new_n310), .A3(new_n318), .A4(new_n315), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G183gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT27), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G183gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT27), .B(G183gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT67), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(G190gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  INV_X1    g138(.A(G190gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n328), .A2(new_n330), .A3(new_n339), .A4(new_n340), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n336), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT26), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n345), .A2(KEYINPUT26), .ZN(new_n347));
  INV_X1    g146(.A(G169gat), .ZN(new_n348));
  INV_X1    g147(.A(G176gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI221_X1 g149(.A(new_n346), .B1(new_n327), .B2(new_n340), .C1(new_n347), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n345), .B2(KEYINPUT65), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n355), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n350), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n357), .A2(new_n362), .A3(KEYINPUT25), .A4(new_n363), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n344), .A2(new_n352), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G226gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(new_n245), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT70), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT70), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n366), .A2(new_n367), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT66), .B1(new_n331), .B2(G190gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n336), .A3(new_n342), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n351), .B1(new_n376), .B2(new_n338), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n373), .B(new_n370), .C1(new_n374), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n371), .B1(new_n368), .B2(KEYINPUT29), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n238), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n344), .A2(new_n352), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n370), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n385), .A3(new_n238), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT71), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT71), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n240), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n372), .A2(new_n378), .B1(new_n390), .B2(new_n371), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n389), .B(new_n386), .C1(new_n391), .C2(new_n238), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n326), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n379), .A2(new_n380), .ZN(new_n394));
  INV_X1    g193(.A(new_n238), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n326), .A3(new_n386), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT30), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n398), .A2(KEYINPUT30), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n320), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n291), .A2(new_n294), .A3(new_n296), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n305), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT82), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n405), .A3(new_n305), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT39), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT83), .B1(new_n407), .B2(new_n315), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n402), .A2(new_n405), .A3(new_n305), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n405), .B1(new_n402), .B2(new_n305), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n409), .B(new_n314), .C1(new_n412), .C2(KEYINPUT39), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n304), .A2(new_n306), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(KEYINPUT39), .C1(new_n305), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT84), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT40), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n417), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT40), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n308), .A2(new_n310), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT6), .B1(new_n424), .B2(new_n314), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n317), .A3(new_n319), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n316), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT37), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n396), .A2(new_n430), .A3(new_n386), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT38), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n325), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n238), .B1(new_n380), .B2(new_n385), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n379), .A2(new_n238), .A3(new_n380), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n391), .A2(KEYINPUT86), .A3(new_n238), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n430), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n397), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n423), .B1(new_n429), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(new_n438), .ZN(new_n444));
  INV_X1    g243(.A(new_n436), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT37), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n381), .A2(new_n387), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n433), .B1(new_n448), .B2(new_n430), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n398), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n450), .A2(KEYINPUT87), .A3(new_n428), .A4(new_n426), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n431), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n388), .A2(new_n392), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n326), .B1(new_n454), .B2(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n455), .B2(KEYINPUT88), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n430), .B1(new_n388), .B2(new_n392), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(new_n326), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n432), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n275), .B(new_n422), .C1(new_n452), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n424), .A2(new_n314), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n427), .A4(new_n316), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n428), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n425), .B2(new_n316), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n399), .B(new_n400), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n268), .B1(new_n263), .B2(new_n264), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n272), .A2(new_n273), .A3(new_n267), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n384), .A2(new_n290), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n368), .A2(new_n295), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G227gat), .A2(G233gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n475), .B(KEYINPUT64), .Z(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G43gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G71gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(G99gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n476), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n472), .A2(new_n486), .A3(new_n473), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT34), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n472), .A2(new_n489), .A3(new_n473), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT33), .B1(new_n474), .B2(new_n476), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n488), .B(new_n490), .C1(new_n493), .C2(new_n483), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n479), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n479), .A3(new_n494), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(KEYINPUT36), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n492), .A2(new_n479), .A3(new_n494), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(new_n495), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n471), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n461), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n500), .A2(new_n495), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n468), .A2(new_n505), .A3(new_n469), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n399), .A2(new_n400), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT35), .B1(new_n426), .B2(new_n428), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT35), .B1(new_n506), .B2(new_n467), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(KEYINPUT89), .A2(G43gat), .ZN(new_n514));
  INV_X1    g313(.A(G50gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(KEYINPUT89), .A2(G43gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT14), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n517), .A2(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527));
  OR2_X1    g326(.A1(G43gat), .A2(G50gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G43gat), .A2(G50gat), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n524), .A2(new_n525), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n530), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT17), .A4(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n534), .B1(new_n526), .B2(new_n530), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(KEYINPUT90), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT16), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(G1gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n540), .A2(G1gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(KEYINPUT91), .ZN(new_n544));
  INV_X1    g343(.A(G1gat), .ZN(new_n545));
  INV_X1    g344(.A(G15gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(G22gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n249), .A2(G15gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(G8gat), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT92), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n542), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G8gat), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n540), .B(KEYINPUT92), .C1(new_n541), .C2(G1gat), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n549), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n537), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n560), .A2(KEYINPUT18), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n558), .B(new_n561), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n563), .B(KEYINPUT13), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n560), .A2(new_n563), .A3(new_n562), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT93), .ZN(new_n572));
  XNOR2_X1  g371(.A(G113gat), .B(G141gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G197gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT11), .B(G169gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT12), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n568), .B(new_n571), .C1(new_n572), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n572), .A3(new_n567), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n569), .A2(new_n570), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n567), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n580), .B(new_n577), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  NAND2_X1  g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G64gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(G57gat), .ZN(new_n590));
  INV_X1    g389(.A(G57gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(G64gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n588), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n585), .B1(new_n593), .B2(KEYINPUT95), .ZN(new_n594));
  XNOR2_X1  g393(.A(G71gat), .B(G78gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(G64gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(G57gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n596), .A2(new_n597), .B1(new_n587), .B2(new_n586), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n598), .B2(KEYINPUT94), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n585), .B(new_n595), .C1(new_n593), .C2(KEYINPUT95), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n558), .B1(KEYINPUT21), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  XOR2_X1   g405(.A(G127gat), .B(G155gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT97), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT96), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n605), .A2(new_n606), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n605), .B2(new_n606), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n600), .A2(new_n601), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n621), .ZN(new_n624));
  OAI22_X1  g423(.A1(new_n614), .A2(new_n615), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n603), .B(new_n604), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n611), .ZN(new_n627));
  INV_X1    g426(.A(new_n624), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n627), .A2(new_n628), .A3(new_n622), .A4(new_n613), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634));
  XOR2_X1   g433(.A(G99gat), .B(G106gat), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(G85gat), .A2(G92gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT7), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT7), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n640), .A2(KEYINPUT99), .A3(G85gat), .A4(G92gat), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n637), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT8), .ZN(new_n643));
  NAND2_X1  g442(.A1(G99gat), .A2(G106gat), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n636), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n636), .B1(new_n642), .B2(new_n647), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n634), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n642), .A2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n635), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(KEYINPUT101), .A3(new_n648), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n633), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n602), .B1(new_n649), .B2(new_n650), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n600), .A2(new_n653), .A3(new_n601), .A4(new_n648), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT10), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n631), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n632), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n633), .A2(new_n655), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(KEYINPUT104), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n660), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n661), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n657), .A2(new_n667), .A3(new_n658), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  AND2_X1   g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n662), .A2(new_n632), .B1(new_n633), .B2(new_n655), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n668), .B1(new_n674), .B2(new_n667), .ZN(new_n675));
  INV_X1    g474(.A(new_n671), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G190gat), .B(G218gat), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n651), .A2(new_n654), .ZN(new_n681));
  AND2_X1   g480(.A1(G232gat), .A2(G233gat), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n539), .A2(new_n681), .B1(KEYINPUT41), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n655), .A2(new_n561), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n680), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n683), .A2(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT102), .ZN(new_n690));
  INV_X1    g489(.A(new_n680), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(G134gat), .B(G162gat), .Z(new_n694));
  AOI21_X1  g493(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(KEYINPUT103), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n688), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n696), .B(KEYINPUT103), .Z(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n688), .B2(new_n693), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n630), .B(new_n679), .C1(new_n699), .C2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n513), .A2(new_n584), .A3(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n465), .A2(new_n466), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(new_n545), .ZN(G1324gat));
  INV_X1    g507(.A(new_n507), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT105), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n705), .B2(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n555), .A2(KEYINPUT42), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT16), .B(G8gat), .Z(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n710), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n715), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1325gat));
  OAI21_X1  g523(.A(G15gat), .B1(new_n705), .B2(new_n502), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n505), .A2(new_n546), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n705), .B2(new_n726), .ZN(G1326gat));
  NOR2_X1   g526(.A1(new_n705), .A2(new_n275), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT43), .B(G22gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  NOR2_X1   g529(.A1(new_n699), .A2(new_n702), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n630), .A3(new_n678), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n513), .A2(new_n584), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n706), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n519), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT45), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n471), .A2(new_n502), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n454), .A2(KEYINPUT37), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(KEYINPUT88), .A3(new_n325), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n459), .A3(new_n431), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT38), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(new_n443), .A3(new_n451), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n418), .B1(new_n416), .B2(new_n417), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n470), .B1(new_n747), .B2(new_n401), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n739), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n275), .A2(new_n709), .A3(new_n706), .A4(new_n505), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n750), .A2(KEYINPUT35), .B1(new_n508), .B2(new_n509), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT108), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n504), .A2(new_n753), .A3(new_n512), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n749), .A2(new_n751), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n757), .B2(new_n732), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n678), .B(KEYINPUT107), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n584), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n761), .A2(new_n762), .A3(new_n630), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G29gat), .B1(new_n764), .B2(new_n706), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n738), .A2(new_n765), .ZN(G1328gat));
  OAI21_X1  g565(.A(G36gat), .B1(new_n764), .B2(new_n709), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n507), .A2(new_n523), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT46), .B1(new_n734), .B2(new_n768), .ZN(new_n769));
  OR3_X1    g568(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n768), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(G1329gat));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n514), .A2(new_n516), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n505), .A2(new_n773), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n734), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n734), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n764), .A2(new_n502), .ZN(new_n778));
  OAI211_X1 g577(.A(KEYINPUT47), .B(new_n777), .C1(new_n778), .C2(new_n773), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780));
  INV_X1    g579(.A(new_n777), .ZN(new_n781));
  INV_X1    g580(.A(new_n763), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n756), .B2(new_n758), .ZN(new_n783));
  INV_X1    g582(.A(new_n502), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n773), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n780), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n779), .A2(new_n786), .ZN(G1330gat));
  INV_X1    g586(.A(KEYINPUT48), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n759), .A2(new_n470), .A3(new_n763), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G50gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n470), .A2(new_n515), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n734), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n788), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AOI211_X1 g593(.A(KEYINPUT48), .B(new_n792), .C1(new_n789), .C2(G50gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(G1331gat));
  INV_X1    g595(.A(new_n630), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n760), .A2(new_n731), .A3(new_n797), .A4(new_n584), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n752), .A2(new_n754), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n752), .A2(new_n754), .A3(KEYINPUT110), .A4(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n736), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G57gat), .ZN(G1332gat));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n507), .A3(new_n802), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n806));
  XOR2_X1   g605(.A(KEYINPUT49), .B(G64gat), .Z(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n805), .B2(new_n807), .ZN(G1333gat));
  NAND3_X1  g607(.A1(new_n801), .A2(new_n784), .A3(new_n802), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G71gat), .ZN(new_n810));
  INV_X1    g609(.A(new_n505), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(G71gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n801), .A2(new_n802), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(KEYINPUT50), .A3(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1334gat));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n470), .A3(new_n802), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g619(.A1(new_n797), .A2(new_n762), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n679), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n759), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G85gat), .B1(new_n823), .B2(new_n706), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(KEYINPUT111), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n513), .A2(new_n731), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n825), .A2(KEYINPUT111), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n828), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n513), .A2(new_n731), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n706), .A2(G85gat), .A3(new_n679), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n824), .A2(new_n833), .ZN(G1336gat));
  INV_X1    g633(.A(G92gat), .ZN(new_n835));
  INV_X1    g634(.A(new_n822), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n756), .B2(new_n758), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(new_n507), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n709), .A2(G92gat), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n829), .A2(new_n761), .A3(new_n831), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n842), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT52), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1337gat));
  NOR3_X1   g645(.A1(new_n811), .A2(G99gat), .A3(new_n679), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n831), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT112), .B1(new_n823), .B2(new_n502), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G99gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n823), .A2(KEYINPUT112), .A3(new_n502), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(G1338gat));
  OAI21_X1  g651(.A(G106gat), .B1(new_n823), .B2(new_n275), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n275), .A2(G106gat), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n829), .A2(new_n761), .A3(new_n831), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n266), .B1(new_n837), .B2(new_n470), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n854), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT53), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n858), .A2(new_n861), .ZN(G1339gat));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n674), .B2(new_n667), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n666), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n674), .A2(new_n667), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n671), .B1(new_n866), .B2(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n865), .A2(KEYINPUT55), .A3(new_n867), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n673), .A3(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n571), .A2(new_n578), .A3(new_n567), .A4(new_n564), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n563), .B1(new_n560), .B2(new_n562), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n565), .A2(new_n566), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n576), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT114), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n731), .B1(new_n872), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n688), .A2(new_n693), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n700), .ZN(new_n884));
  INV_X1    g683(.A(new_n877), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n884), .A2(new_n698), .B1(new_n885), .B2(new_n678), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n584), .A3(new_n673), .A4(new_n871), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n888), .A3(new_n797), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n704), .A2(new_n762), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(new_n736), .A3(new_n508), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n584), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(G113gat), .ZN(G1340gat));
  AOI21_X1  g693(.A(G120gat), .B1(new_n892), .B2(new_n678), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n761), .A2(G120gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n892), .B2(new_n896), .ZN(G1341gat));
  NAND2_X1  g696(.A1(new_n892), .A2(new_n630), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g698(.A1(new_n892), .A2(new_n731), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n900), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(G134gat), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT56), .B1(new_n900), .B2(G134gat), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(KEYINPUT115), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(KEYINPUT115), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n901), .B(new_n902), .C1(new_n904), .C2(new_n905), .ZN(G1343gat));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n891), .B2(new_n470), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT57), .B(new_n275), .C1(new_n889), .C2(new_n890), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n784), .A2(new_n706), .A3(new_n507), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G141gat), .B1(new_n912), .B2(new_n762), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n703), .A2(new_n584), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n868), .A2(new_n869), .B1(new_n666), .B2(new_n672), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n915), .A2(new_n871), .A3(new_n878), .A4(new_n880), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n630), .B1(new_n916), .B2(new_n731), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n917), .B2(new_n888), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n275), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(new_n911), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n762), .A2(G141gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n913), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g723(.A(G148gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(new_n925), .A3(new_n678), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n470), .A2(KEYINPUT117), .A3(new_n907), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(new_n908), .B2(new_n909), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT57), .B1(new_n918), .B2(new_n275), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n891), .A2(new_n907), .A3(new_n470), .ZN(new_n931));
  INV_X1    g730(.A(new_n928), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n929), .A2(new_n678), .A3(new_n911), .A4(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n927), .B1(new_n934), .B2(G148gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n910), .A2(new_n678), .A3(new_n911), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n926), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT118), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n941), .B(new_n926), .C1(new_n935), .C2(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1345gat));
  OAI21_X1  g742(.A(G155gat), .B1(new_n912), .B2(new_n797), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n797), .A2(G155gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n921), .B2(new_n945), .ZN(G1346gat));
  INV_X1    g745(.A(G162gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n912), .A2(new_n947), .A3(new_n732), .ZN(new_n948));
  AOI21_X1  g747(.A(G162gat), .B1(new_n920), .B2(new_n731), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(G1347gat));
  NOR2_X1   g749(.A1(new_n918), .A2(new_n736), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT119), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n918), .B2(new_n736), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n506), .A2(new_n709), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT120), .A4(new_n955), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n958), .A2(new_n348), .A3(new_n584), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n951), .A2(new_n955), .ZN(new_n961));
  OAI21_X1  g760(.A(G169gat), .B1(new_n961), .B2(new_n762), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n963), .B(new_n964), .ZN(G1348gat));
  NAND4_X1  g764(.A1(new_n958), .A2(new_n349), .A3(new_n678), .A4(new_n959), .ZN(new_n966));
  OAI21_X1  g765(.A(G176gat), .B1(new_n961), .B2(new_n760), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1349gat));
  OAI21_X1  g767(.A(G183gat), .B1(new_n961), .B2(new_n797), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n630), .A2(new_n333), .A3(new_n335), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n956), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g770(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n972));
  XNOR2_X1  g771(.A(new_n971), .B(new_n972), .ZN(G1350gat));
  OAI21_X1  g772(.A(G190gat), .B1(new_n961), .B2(new_n732), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT123), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(KEYINPUT123), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(KEYINPUT61), .A3(new_n976), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n958), .A2(new_n340), .A3(new_n731), .A4(new_n959), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n974), .A2(KEYINPUT123), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(G1351gat));
  AOI21_X1  g780(.A(new_n932), .B1(new_n930), .B2(new_n931), .ZN(new_n982));
  AND4_X1   g781(.A1(KEYINPUT117), .A2(new_n918), .A3(new_n907), .A4(new_n470), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n502), .A2(new_n507), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(new_n706), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n984), .A2(new_n584), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g788(.A(KEYINPUT124), .B(G197gat), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n952), .A2(new_n954), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n985), .A2(new_n275), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n993), .A2(new_n584), .A3(new_n990), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT125), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n992), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n997), .A2(new_n999), .ZN(G1352gat));
  NOR2_X1   g799(.A1(new_n679), .A2(G204gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n993), .A2(new_n994), .A3(new_n1001), .ZN(new_n1002));
  XOR2_X1   g801(.A(new_n1002), .B(KEYINPUT62), .Z(new_n1003));
  NAND3_X1  g802(.A1(new_n984), .A2(new_n761), .A3(new_n988), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(G204gat), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n1005), .ZN(G1353gat));
  NAND4_X1  g805(.A1(new_n993), .A2(new_n226), .A3(new_n630), .A4(new_n994), .ZN(new_n1007));
  NOR4_X1   g806(.A1(new_n982), .A2(new_n983), .A3(new_n797), .A4(new_n987), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n226), .B1(new_n1008), .B2(KEYINPUT126), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n929), .A2(new_n630), .A3(new_n933), .A4(new_n988), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g811(.A(KEYINPUT63), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n984), .A2(KEYINPUT126), .A3(new_n630), .A4(new_n988), .ZN(new_n1014));
  AND4_X1   g813(.A1(KEYINPUT63), .A2(new_n1014), .A3(new_n1012), .A4(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1007), .B1(new_n1013), .B2(new_n1015), .ZN(G1354gat));
  NAND3_X1  g815(.A1(new_n993), .A2(new_n731), .A3(new_n994), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(new_n227), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1017), .A2(KEYINPUT127), .A3(new_n227), .ZN(new_n1021));
  NAND4_X1  g820(.A1(new_n984), .A2(G218gat), .A3(new_n731), .A4(new_n988), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(G1355gat));
endmodule


