

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590;

  XNOR2_X1 U322 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U323 ( .A(n445), .B(n322), .ZN(n324) );
  INV_X1 U324 ( .A(n361), .ZN(n328) );
  XNOR2_X1 U325 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U326 ( .A(n459), .B(KEYINPUT121), .ZN(n460) );
  XNOR2_X1 U327 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U328 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U329 ( .A(n466), .B(G190GAT), .ZN(n467) );
  XNOR2_X1 U330 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT0), .B(KEYINPUT81), .Z(n291) );
  XNOR2_X1 U332 ( .A(KEYINPUT80), .B(G127GAT), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U334 ( .A(G113GAT), .B(n292), .Z(n439) );
  XOR2_X1 U335 ( .A(G134GAT), .B(G190GAT), .Z(n294) );
  XNOR2_X1 U336 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n310) );
  XOR2_X1 U338 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n296) );
  XNOR2_X1 U339 ( .A(G120GAT), .B(KEYINPUT20), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U341 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n298) );
  XNOR2_X1 U342 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(KEYINPUT18), .B(n299), .Z(n416) );
  XOR2_X1 U345 ( .A(n300), .B(n416), .Z(n308) );
  XOR2_X1 U346 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n302) );
  XNOR2_X1 U347 ( .A(G15GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U349 ( .A(G176GAT), .B(G99GAT), .Z(n304) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G43GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U354 ( .A(n310), .B(n309), .Z(n312) );
  NAND2_X1 U355 ( .A1(G227GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U357 ( .A(n439), .B(n313), .ZN(n534) );
  XNOR2_X1 U358 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n355) );
  INV_X1 U359 ( .A(G148GAT), .ZN(n314) );
  NAND2_X1 U360 ( .A1(G78GAT), .A2(n314), .ZN(n317) );
  INV_X1 U361 ( .A(G78GAT), .ZN(n315) );
  NAND2_X1 U362 ( .A1(n315), .A2(G148GAT), .ZN(n316) );
  NAND2_X1 U363 ( .A1(n317), .A2(n316), .ZN(n319) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n445) );
  NAND2_X1 U366 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  INV_X1 U367 ( .A(KEYINPUT33), .ZN(n320) );
  INV_X1 U368 ( .A(KEYINPUT32), .ZN(n323) );
  NAND2_X1 U369 ( .A1(n324), .A2(n323), .ZN(n327) );
  INV_X1 U370 ( .A(n324), .ZN(n325) );
  NAND2_X1 U371 ( .A1(n325), .A2(KEYINPUT32), .ZN(n326) );
  NAND2_X1 U372 ( .A1(n327), .A2(n326), .ZN(n331) );
  XOR2_X1 U373 ( .A(G71GAT), .B(KEYINPUT13), .Z(n384) );
  XNOR2_X1 U374 ( .A(n384), .B(KEYINPUT31), .ZN(n329) );
  XOR2_X1 U375 ( .A(G99GAT), .B(G85GAT), .Z(n361) );
  XOR2_X1 U376 ( .A(G120GAT), .B(G57GAT), .Z(n431) );
  XOR2_X1 U377 ( .A(G64GAT), .B(G92GAT), .Z(n333) );
  XNOR2_X1 U378 ( .A(G176GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U379 ( .A(n333), .B(n332), .ZN(n407) );
  XNOR2_X1 U380 ( .A(n431), .B(n407), .ZN(n334) );
  XNOR2_X1 U381 ( .A(n335), .B(n334), .ZN(n579) );
  XNOR2_X1 U382 ( .A(KEYINPUT41), .B(n579), .ZN(n556) );
  XOR2_X1 U383 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n337) );
  XNOR2_X1 U384 ( .A(G197GAT), .B(G141GAT), .ZN(n336) );
  XNOR2_X1 U385 ( .A(n337), .B(n336), .ZN(n353) );
  XOR2_X1 U386 ( .A(G169GAT), .B(G8GAT), .Z(n404) );
  XOR2_X1 U387 ( .A(G113GAT), .B(G50GAT), .Z(n339) );
  XNOR2_X1 U388 ( .A(G36GAT), .B(G29GAT), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U390 ( .A(n404), .B(n340), .Z(n342) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U393 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n344) );
  XNOR2_X1 U394 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U396 ( .A(n346), .B(n345), .Z(n351) );
  XNOR2_X1 U397 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n347), .B(KEYINPUT8), .ZN(n363) );
  XOR2_X1 U399 ( .A(KEYINPUT69), .B(G1GAT), .Z(n349) );
  XNOR2_X1 U400 ( .A(G15GAT), .B(G22GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n388) );
  XNOR2_X1 U402 ( .A(n363), .B(n388), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U404 ( .A(n353), .B(n352), .Z(n551) );
  INV_X1 U405 ( .A(n551), .ZN(n575) );
  AND2_X1 U406 ( .A1(n556), .A2(n575), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n394) );
  XOR2_X1 U408 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n357) );
  XNOR2_X1 U409 ( .A(G92GAT), .B(KEYINPUT65), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(G50GAT), .B(G162GAT), .Z(n441) );
  XOR2_X1 U412 ( .A(n358), .B(n441), .Z(n360) );
  XNOR2_X1 U413 ( .A(G218GAT), .B(G106GAT), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n365) );
  XOR2_X1 U416 ( .A(G29GAT), .B(G134GAT), .Z(n435) );
  XOR2_X1 U417 ( .A(n363), .B(n435), .Z(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n374) );
  XOR2_X1 U419 ( .A(KEYINPUT74), .B(KEYINPUT64), .Z(n367) );
  XNOR2_X1 U420 ( .A(KEYINPUT73), .B(KEYINPUT9), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n372) );
  XNOR2_X1 U422 ( .A(G36GAT), .B(G190GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n368), .B(KEYINPUT76), .ZN(n412) );
  XOR2_X1 U424 ( .A(KEYINPUT10), .B(n412), .Z(n370) );
  NAND2_X1 U425 ( .A1(G232GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n563) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G57GAT), .Z(n376) );
  XNOR2_X1 U430 ( .A(G8GAT), .B(G155GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U432 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n378) );
  XNOR2_X1 U433 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n392) );
  XOR2_X1 U436 ( .A(G78GAT), .B(G211GAT), .Z(n382) );
  XNOR2_X1 U437 ( .A(G127GAT), .B(G183GAT), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U439 ( .A(n384), .B(n383), .Z(n386) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U442 ( .A(n387), .B(KEYINPUT79), .Z(n390) );
  XNOR2_X1 U443 ( .A(n388), .B(KEYINPUT15), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U445 ( .A(n392), .B(n391), .Z(n583) );
  INV_X1 U446 ( .A(n583), .ZN(n560) );
  NAND2_X1 U447 ( .A1(n563), .A2(n560), .ZN(n393) );
  OR2_X1 U448 ( .A1(n394), .A2(n393), .ZN(n395) );
  XNOR2_X1 U449 ( .A(KEYINPUT47), .B(n395), .ZN(n396) );
  XNOR2_X1 U450 ( .A(KEYINPUT113), .B(n396), .ZN(n402) );
  INV_X1 U451 ( .A(n563), .ZN(n544) );
  XOR2_X1 U452 ( .A(n544), .B(KEYINPUT36), .Z(n587) );
  NOR2_X1 U453 ( .A1(n560), .A2(n587), .ZN(n397) );
  XNOR2_X1 U454 ( .A(KEYINPUT45), .B(n397), .ZN(n398) );
  NAND2_X1 U455 ( .A1(n398), .A2(n579), .ZN(n399) );
  NOR2_X1 U456 ( .A1(n575), .A2(n399), .ZN(n400) );
  XOR2_X1 U457 ( .A(KEYINPUT114), .B(n400), .Z(n401) );
  AND2_X1 U458 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U459 ( .A(KEYINPUT48), .B(n403), .ZN(n549) );
  XOR2_X1 U460 ( .A(KEYINPUT99), .B(n404), .Z(n406) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U463 ( .A(n408), .B(n407), .Z(n414) );
  XOR2_X1 U464 ( .A(KEYINPUT91), .B(G218GAT), .Z(n410) );
  XNOR2_X1 U465 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U467 ( .A(G197GAT), .B(n411), .Z(n455) );
  XNOR2_X1 U468 ( .A(n455), .B(n412), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n523) );
  NOR2_X1 U471 ( .A1(n549), .A2(n523), .ZN(n419) );
  XOR2_X1 U472 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n417) );
  XNOR2_X1 U473 ( .A(KEYINPUT54), .B(n417), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n570) );
  XOR2_X1 U475 ( .A(KEYINPUT1), .B(G85GAT), .Z(n421) );
  XNOR2_X1 U476 ( .A(G148GAT), .B(G162GAT), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U478 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n423) );
  XNOR2_X1 U479 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U481 ( .A(n425), .B(n424), .Z(n430) );
  XOR2_X1 U482 ( .A(KEYINPUT97), .B(KEYINPUT6), .Z(n427) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(KEYINPUT4), .B(n428), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U487 ( .A(n432), .B(n431), .Z(n437) );
  XOR2_X1 U488 ( .A(G155GAT), .B(KEYINPUT2), .Z(n434) );
  XNOR2_X1 U489 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n440), .B(n435), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n475) );
  XOR2_X1 U494 ( .A(KEYINPUT98), .B(n475), .Z(n478) );
  XOR2_X1 U495 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U498 ( .A(n444), .B(KEYINPUT22), .Z(n447) );
  XNOR2_X1 U499 ( .A(n445), .B(KEYINPUT89), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U501 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n449) );
  XNOR2_X1 U502 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U504 ( .A(n451), .B(n450), .Z(n457) );
  XOR2_X1 U505 ( .A(KEYINPUT90), .B(G204GAT), .Z(n453) );
  XNOR2_X1 U506 ( .A(G22GAT), .B(KEYINPUT94), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(n479) );
  NOR2_X1 U510 ( .A1(n478), .A2(n479), .ZN(n458) );
  AND2_X1 U511 ( .A1(n570), .A2(n458), .ZN(n461) );
  INV_X1 U512 ( .A(KEYINPUT55), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n534), .A2(n462), .ZN(n567) );
  NAND2_X1 U514 ( .A1(n567), .A2(n556), .ZN(n465) );
  XOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(G176GAT), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  NAND2_X1 U518 ( .A1(n567), .A2(n544), .ZN(n468) );
  XOR2_X1 U519 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n466) );
  INV_X1 U520 ( .A(n478), .ZN(n571) );
  NOR2_X1 U521 ( .A1(n534), .A2(n523), .ZN(n469) );
  NOR2_X1 U522 ( .A1(n479), .A2(n469), .ZN(n470) );
  XNOR2_X1 U523 ( .A(n470), .B(KEYINPUT25), .ZN(n474) );
  NAND2_X1 U524 ( .A1(n534), .A2(n479), .ZN(n471) );
  XNOR2_X1 U525 ( .A(n471), .B(KEYINPUT26), .ZN(n472) );
  XOR2_X1 U526 ( .A(KEYINPUT100), .B(n472), .Z(n569) );
  XOR2_X1 U527 ( .A(KEYINPUT27), .B(n523), .Z(n477) );
  NAND2_X1 U528 ( .A1(n569), .A2(n477), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n476) );
  NAND2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n482) );
  NAND2_X1 U531 ( .A1(n478), .A2(n477), .ZN(n548) );
  XOR2_X1 U532 ( .A(n479), .B(KEYINPUT28), .Z(n530) );
  INV_X1 U533 ( .A(n530), .ZN(n480) );
  NOR2_X1 U534 ( .A1(n548), .A2(n480), .ZN(n536) );
  NAND2_X1 U535 ( .A1(n536), .A2(n534), .ZN(n481) );
  NAND2_X1 U536 ( .A1(n482), .A2(n481), .ZN(n496) );
  NAND2_X1 U537 ( .A1(n563), .A2(n583), .ZN(n483) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  AND2_X1 U539 ( .A1(n496), .A2(n484), .ZN(n510) );
  NAND2_X1 U540 ( .A1(n575), .A2(n579), .ZN(n485) );
  XOR2_X1 U541 ( .A(KEYINPUT72), .B(n485), .Z(n499) );
  NAND2_X1 U542 ( .A1(n510), .A2(n499), .ZN(n494) );
  NOR2_X1 U543 ( .A1(n571), .A2(n494), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NOR2_X1 U547 ( .A1(n523), .A2(n494), .ZN(n489) );
  XOR2_X1 U548 ( .A(G8GAT), .B(n489), .Z(G1325GAT) );
  NOR2_X1 U549 ( .A1(n494), .A2(n534), .ZN(n493) );
  XOR2_X1 U550 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n491) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  NOR2_X1 U554 ( .A1(n530), .A2(n494), .ZN(n495) );
  XOR2_X1 U555 ( .A(G22GAT), .B(n495), .Z(G1327GAT) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n502) );
  NOR2_X1 U557 ( .A1(n583), .A2(n587), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(KEYINPUT37), .B(n498), .ZN(n521) );
  NAND2_X1 U560 ( .A1(n521), .A2(n499), .ZN(n500) );
  XNOR2_X1 U561 ( .A(KEYINPUT38), .B(n500), .ZN(n506) );
  NOR2_X1 U562 ( .A1(n571), .A2(n506), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n506), .A2(n523), .ZN(n503) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  NOR2_X1 U566 ( .A1(n506), .A2(n534), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT40), .B(n504), .Z(n505) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  NOR2_X1 U569 ( .A1(n530), .A2(n506), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT104), .B(n507), .Z(n508) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  NAND2_X1 U572 ( .A1(n556), .A2(n551), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT105), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n520), .A2(n510), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n571), .A2(n517), .ZN(n511) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n523), .A2(n517), .ZN(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U582 ( .A1(n534), .A2(n517), .ZN(n516) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U584 ( .A1(n530), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n529) );
  NOR2_X1 U588 ( .A1(n571), .A2(n529), .ZN(n522) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n529), .ZN(n524) );
  XOR2_X1 U591 ( .A(KEYINPUT108), .B(n524), .Z(n525) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n525), .ZN(G1337GAT) );
  NOR2_X1 U593 ( .A1(n534), .A2(n529), .ZN(n527) );
  XNOR2_X1 U594 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(n528), .ZN(G1338GAT) );
  NOR2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U601 ( .A1(n534), .A2(n549), .ZN(n535) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT115), .B(n537), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n575), .A2(n545), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U607 ( .A1(n545), .A2(n556), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n542) );
  NAND2_X1 U610 ( .A1(n545), .A2(n583), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n569), .A2(n550), .ZN(n562) );
  NOR2_X1 U618 ( .A1(n551), .A2(n562), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n559) );
  INV_X1 U624 ( .A(n556), .ZN(n557) );
  NOR2_X1 U625 ( .A1(n557), .A2(n562), .ZN(n558) );
  XOR2_X1 U626 ( .A(n559), .B(n558), .Z(G1345GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n562), .ZN(n561) );
  XOR2_X1 U628 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  NAND2_X1 U631 ( .A1(n575), .A2(n567), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  NAND2_X1 U634 ( .A1(n583), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  INV_X1 U637 ( .A(n569), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(n574), .B(KEYINPUT124), .Z(n588) );
  INV_X1 U641 ( .A(n588), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n581) );
  OR2_X1 U646 ( .A1(n588), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(KEYINPUT126), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

