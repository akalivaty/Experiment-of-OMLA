//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919;
  AOI21_X1  g000(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT96), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204));
  INV_X1    g003(.A(G64gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT95), .B1(new_n205), .B2(G57gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT95), .ZN(new_n207));
  INV_X1    g006(.A(G57gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(G64gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n206), .B(new_n209), .C1(new_n208), .C2(G64gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n203), .A2(new_n204), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT97), .ZN(new_n212));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(new_n204), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT21), .ZN(new_n218));
  XOR2_X1   g017(.A(G15gat), .B(G22gat), .Z(new_n219));
  INV_X1    g018(.A(G1gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  INV_X1    g023(.A(G8gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n221), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT93), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n221), .A2(new_n224), .A3(KEYINPUT92), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n228), .B(G8gat), .C1(KEYINPUT92), .C2(new_n224), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n218), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G127gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n217), .A2(KEYINPUT21), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT98), .B(G211gat), .Z(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G231gat), .A2(G233gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n235), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G155gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n241), .B(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G50gat), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n245), .A2(G43gat), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT91), .B(G43gat), .Z(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n247), .B2(G50gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT15), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(G43gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n251), .A3(KEYINPUT15), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT89), .B(G29gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT90), .B(G36gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(G29gat), .A2(G36gat), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n254), .A2(new_n255), .B1(KEYINPUT14), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(KEYINPUT14), .B2(new_n256), .ZN(new_n258));
  MUX2_X1   g057(.A(new_n253), .B(new_n252), .S(new_n258), .Z(new_n259));
  INV_X1    g058(.A(G85gat), .ZN(new_n260));
  INV_X1    g059(.A(G92gat), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT99), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT99), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(G85gat), .A3(G92gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G99gat), .A2(G106gat), .ZN(new_n266));
  AOI22_X1  g065(.A1(KEYINPUT8), .A2(new_n266), .B1(new_n260), .B2(new_n261), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT7), .ZN(new_n268));
  OAI211_X1 g067(.A(KEYINPUT99), .B(new_n268), .C1(new_n260), .C2(new_n261), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G99gat), .B(G106gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT17), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n259), .B(new_n273), .Z(new_n274));
  NAND3_X1  g073(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G190gat), .B(G218gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT100), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G134gat), .B(G162gat), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n279), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n285), .A3(new_n283), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n244), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G78gat), .B(G106gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT31), .B(G50gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G22gat), .ZN(new_n292));
  INV_X1    g091(.A(G22gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT86), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT22), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G211gat), .B(G218gat), .Z(new_n303));
  OR2_X1    g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n303), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT3), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(new_n309), .B2(new_n308), .ZN(new_n311));
  INV_X1    g110(.A(G141gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G148gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT81), .B(G148gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(new_n312), .ZN(new_n315));
  OR2_X1    g114(.A1(KEYINPUT82), .A2(G162gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT82), .A2(G162gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(G155gat), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n319));
  OR2_X1    g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n315), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n321), .B(KEYINPUT80), .ZN(new_n324));
  XNOR2_X1  g123(.A(G141gat), .B(G148gat), .ZN(new_n325));
  AND2_X1   g124(.A1(KEYINPUT80), .A2(KEYINPUT2), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n324), .B(new_n320), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n306), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n307), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n311), .A2(new_n328), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G228gat), .ZN(new_n334));
  INV_X1    g133(.A(G233gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n306), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n332), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n328), .A2(KEYINPUT3), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n328), .A2(new_n306), .A3(new_n307), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n342), .A2(new_n336), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n296), .B1(new_n337), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n333), .A2(new_n336), .ZN(new_n346));
  INV_X1    g145(.A(new_n344), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n346), .A2(new_n347), .A3(new_n295), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT37), .ZN(new_n350));
  NOR2_X1   g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n363));
  AND2_X1   g162(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n364));
  AND2_X1   g163(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n363), .A2(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT66), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT65), .B(G190gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT27), .B(G183gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT66), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n373));
  AND3_X1   g172(.A1(new_n368), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT28), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT68), .B1(new_n367), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT68), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n369), .A2(new_n370), .A3(new_n377), .A4(KEYINPUT28), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n362), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n351), .A2(KEYINPUT23), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n358), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n232), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT24), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n360), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  OR3_X1    g191(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n393), .A2(new_n388), .A3(new_n389), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n392), .A2(KEYINPUT25), .B1(new_n397), .B2(new_n385), .ZN(new_n398));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n380), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n307), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n380), .B2(new_n398), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n400), .A2(new_n403), .A3(new_n329), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n306), .B(KEYINPUT77), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n376), .A2(new_n378), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n368), .A2(new_n372), .A3(new_n373), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n361), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n396), .A3(new_n395), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n384), .B1(new_n386), .B2(new_n390), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n396), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n401), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n380), .A2(new_n398), .A3(new_n399), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n405), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT78), .B1(new_n404), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n339), .B1(new_n400), .B2(new_n403), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n413), .A3(new_n306), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n350), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n350), .A3(new_n418), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT38), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n404), .A2(new_n414), .A3(new_n424), .ZN(new_n427));
  INV_X1    g226(.A(new_n425), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n306), .B1(new_n400), .B2(new_n403), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n339), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(KEYINPUT37), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT38), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G1gat), .B(G29gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(G85gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT0), .B(G57gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n440));
  INV_X1    g239(.A(G134gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(G127gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT1), .B1(new_n441), .B2(G127gat), .ZN(new_n444));
  INV_X1    g243(.A(G113gat), .ZN(new_n445));
  INV_X1    g244(.A(G120gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT70), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT70), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G120gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n446), .A2(G113gat), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n443), .B(new_n444), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n441), .A2(KEYINPUT69), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT69), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G134gat), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n234), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G113gat), .B(G120gat), .ZN(new_n457));
  OAI22_X1  g256(.A1(new_n456), .A2(new_n442), .B1(KEYINPUT1), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n328), .B(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT83), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n440), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n452), .A2(new_n458), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT4), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n323), .A4(new_n327), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT4), .B1(new_n328), .B2(new_n459), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n462), .B1(new_n328), .B2(new_n459), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n341), .A2(new_n459), .A3(new_n331), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n331), .A2(new_n459), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n341), .A2(new_n473), .B1(new_n466), .B2(new_n467), .ZN(new_n474));
  INV_X1    g273(.A(new_n462), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n440), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n439), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT84), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(KEYINPUT84), .A3(KEYINPUT6), .ZN(new_n480));
  INV_X1    g279(.A(new_n477), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n472), .A2(new_n476), .A3(new_n439), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n349), .B1(new_n435), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n424), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n418), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT79), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n417), .B1(new_n416), .B2(new_n418), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n424), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT30), .ZN(new_n494));
  INV_X1    g293(.A(new_n427), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT39), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n468), .A2(new_n470), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(new_n462), .ZN(new_n500));
  AOI211_X1 g299(.A(KEYINPUT87), .B(new_n475), .C1(new_n468), .C2(new_n470), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT87), .B1(new_n474), .B2(new_n475), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n498), .A3(new_n462), .ZN(new_n504));
  INV_X1    g303(.A(new_n460), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n497), .B1(new_n505), .B2(new_n475), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n439), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n502), .A2(new_n507), .A3(KEYINPUT40), .A4(new_n439), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n481), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT88), .B1(new_n486), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n345), .A2(new_n348), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n431), .A2(new_n432), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n495), .B1(new_n425), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT37), .B1(new_n491), .B2(new_n492), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n428), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n519), .B2(KEYINPUT38), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n483), .A2(new_n482), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n477), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n472), .A2(new_n476), .ZN(new_n523));
  INV_X1    g322(.A(new_n439), .ZN(new_n524));
  AND4_X1   g323(.A1(KEYINPUT84), .A2(new_n523), .A3(KEYINPUT6), .A4(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n522), .A2(new_n525), .A3(new_n478), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n515), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n488), .B(KEYINPUT79), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n415), .A2(new_n419), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n424), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n531), .B2(new_n427), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(new_n481), .A3(new_n511), .A4(new_n510), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n514), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n515), .B1(new_n526), .B2(new_n532), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n380), .A2(new_n398), .A3(new_n464), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n459), .B1(new_n408), .B2(new_n411), .ZN(new_n541));
  NAND2_X1  g340(.A1(G227gat), .A2(G233gat), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n380), .A2(new_n398), .A3(KEYINPUT71), .A4(new_n464), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT34), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT73), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n544), .B2(KEYINPUT73), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n551));
  INV_X1    g350(.A(new_n542), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT33), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT72), .B(G71gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G99gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(G15gat), .B(G43gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n553), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  AOI221_X4 g359(.A(new_n550), .B1(KEYINPUT33), .B2(new_n558), .C1(new_n551), .C2(new_n552), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n549), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT74), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n551), .A2(new_n552), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n559), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n553), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n561), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n544), .A2(KEYINPUT73), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT34), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n546), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n562), .A2(new_n563), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n549), .B(KEYINPUT74), .C1(new_n560), .C2(new_n561), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT36), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n578), .A3(new_n573), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n568), .A2(new_n569), .A3(new_n572), .A4(KEYINPUT76), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n536), .A2(new_n537), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n580), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n526), .A2(new_n532), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n349), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n515), .B1(new_n574), .B2(new_n575), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n589), .A2(new_n587), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n590), .B2(new_n586), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n288), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(new_n230), .B2(KEYINPUT94), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n259), .B2(KEYINPUT17), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n594), .A2(new_n259), .B1(new_n596), .B2(new_n230), .ZN(new_n597));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT18), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n230), .B(new_n259), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n598), .B(KEYINPUT13), .Z(new_n603));
  AND2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606));
  INV_X1    g405(.A(G197gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT11), .B(G169gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n217), .B(new_n272), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n217), .A2(KEYINPUT10), .A3(new_n272), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n620), .B2(KEYINPUT10), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n624), .A2(KEYINPUT101), .A3(new_n622), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT101), .B1(new_n624), .B2(new_n622), .ZN(new_n626));
  OAI221_X1 g425(.A(new_n619), .B1(new_n621), .B2(new_n622), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n624), .A2(new_n622), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n621), .A2(new_n622), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n618), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n592), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n526), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g434(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n223), .A2(new_n225), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n633), .A2(new_n532), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n225), .B1(new_n633), .B2(new_n532), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT102), .Z(G1325gat));
  AOI21_X1  g443(.A(G15gat), .B1(new_n633), .B2(new_n585), .ZN(new_n645));
  INV_X1    g444(.A(new_n583), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n633), .B2(new_n647), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n515), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT43), .B(G22gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  AOI21_X1  g450(.A(new_n287), .B1(new_n591), .B2(new_n584), .ZN(new_n652));
  INV_X1    g451(.A(new_n244), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n652), .A2(new_n632), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(new_n485), .A3(new_n254), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT45), .Z(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n658), .B(new_n287), .C1(new_n591), .C2(new_n584), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n584), .A2(KEYINPUT104), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n536), .A2(new_n661), .A3(new_n583), .A4(new_n537), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n591), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n287), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n659), .B1(new_n665), .B2(new_n658), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n244), .B(KEYINPUT103), .Z(new_n667));
  AND3_X1   g466(.A1(new_n666), .A2(new_n632), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n254), .B1(new_n669), .B2(new_n485), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n657), .A2(new_n670), .ZN(G1328gat));
  OAI21_X1  g470(.A(new_n255), .B1(new_n669), .B2(new_n496), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n655), .A2(new_n255), .A3(new_n496), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT46), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1329gat));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n247), .B1(new_n668), .B2(new_n646), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n654), .A2(new_n247), .A3(new_n585), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g479(.A(G50gat), .B1(new_n669), .B2(new_n349), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n654), .B(KEYINPUT106), .Z(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n245), .A3(new_n515), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT48), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1331gat));
  NOR2_X1   g485(.A1(new_n288), .A2(new_n614), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n663), .A2(new_n631), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n526), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g489(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n532), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT107), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1333gat));
  NAND3_X1  g494(.A1(new_n688), .A2(G71gat), .A3(new_n646), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n688), .A2(new_n585), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(G71gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g498(.A1(new_n688), .A2(new_n515), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT108), .B(G78gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1335gat));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n663), .B2(new_n664), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n653), .A2(new_n615), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(new_n659), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n631), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(new_n260), .A3(new_n485), .ZN(new_n707));
  INV_X1    g506(.A(new_n631), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n665), .A2(KEYINPUT109), .ZN(new_n709));
  INV_X1    g508(.A(new_n704), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n663), .A2(new_n711), .A3(new_n664), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n709), .A2(KEYINPUT51), .A3(new_n710), .A4(new_n712), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n708), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n526), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n707), .B1(new_n718), .B2(new_n260), .ZN(G1336gat));
  NOR2_X1   g518(.A1(new_n496), .A2(G92gat), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n663), .A2(new_n711), .A3(new_n664), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n711), .B1(new_n663), .B2(new_n664), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT51), .B1(new_n723), .B2(new_n710), .ZN(new_n724));
  INV_X1    g523(.A(new_n716), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n631), .B(new_n720), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n666), .A2(new_n631), .A3(new_n532), .A4(new_n710), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(G92gat), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT52), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT52), .B1(new_n717), .B2(new_n720), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n705), .A2(KEYINPUT110), .A3(new_n631), .A4(new_n532), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(G92gat), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n731), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738));
  AND4_X1   g537(.A1(new_n731), .A2(new_n726), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n730), .B1(new_n737), .B2(new_n739), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n706), .B2(new_n583), .ZN(new_n741));
  INV_X1    g540(.A(new_n717), .ZN(new_n742));
  INV_X1    g541(.A(new_n585), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(G99gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n742), .B2(new_n744), .ZN(G1338gat));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n666), .A2(new_n631), .A3(new_n515), .A4(new_n710), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G106gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n724), .A2(new_n725), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n708), .A2(G106gat), .A3(new_n349), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n746), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(KEYINPUT112), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n748), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT113), .B1(new_n754), .B2(KEYINPUT53), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n715), .B2(new_n716), .ZN(new_n756));
  INV_X1    g555(.A(new_n748), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT113), .B(KEYINPUT53), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n751), .B1(new_n755), .B2(new_n759), .ZN(G1339gat));
  NOR2_X1   g559(.A1(new_n532), .A2(new_n485), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n624), .A2(new_n622), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT54), .B(new_n763), .C1(new_n625), .C2(new_n626), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n628), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n618), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n764), .A2(KEYINPUT55), .A3(new_n618), .A4(new_n766), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n627), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT115), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n769), .A2(new_n773), .A3(new_n627), .A4(new_n770), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n614), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n597), .A2(new_n599), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n603), .B2(new_n602), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n605), .A2(new_n611), .B1(new_n610), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n631), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n664), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n778), .A2(new_n284), .A3(new_n286), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n772), .A2(new_n781), .A3(new_n774), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n667), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n288), .A2(new_n631), .A3(new_n614), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n762), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n589), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n445), .A3(new_n614), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n743), .A2(new_n515), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n787), .A2(KEYINPUT116), .A3(new_n790), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n614), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n795), .A2(KEYINPUT117), .A3(G113gat), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT117), .B1(new_n795), .B2(G113gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n789), .B1(new_n796), .B2(new_n797), .ZN(G1340gat));
  NAND2_X1  g597(.A1(new_n447), .A2(new_n449), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n788), .A2(new_n799), .A3(new_n631), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n793), .A2(new_n794), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n631), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n802), .B2(new_n446), .ZN(G1341gat));
  AOI21_X1  g602(.A(G127gat), .B1(new_n788), .B2(new_n244), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n667), .A2(new_n234), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n801), .B2(new_n805), .ZN(G1342gat));
  NAND2_X1  g605(.A1(new_n453), .A2(new_n455), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n807), .A3(new_n664), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT56), .Z(new_n809));
  NAND2_X1  g608(.A1(new_n801), .A2(new_n664), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G134gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1343gat));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n349), .B1(new_n784), .B2(new_n786), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n646), .A2(new_n762), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n779), .B1(new_n615), .B2(new_n771), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n287), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n244), .B1(new_n820), .B2(new_n782), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n515), .B1(new_n821), .B2(new_n785), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n818), .B1(new_n822), .B2(KEYINPUT57), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n816), .A2(new_n823), .A3(new_n614), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n784), .A2(new_n786), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n515), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(G141gat), .A3(new_n818), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n824), .A2(G141gat), .B1(new_n827), .B2(new_n614), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n813), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n824), .A2(G141gat), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n312), .A3(new_n614), .A4(new_n817), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(KEYINPUT118), .A3(KEYINPUT58), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT58), .B1(new_n832), .B2(KEYINPUT119), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n831), .B(new_n835), .C1(KEYINPUT119), .C2(new_n832), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n830), .A2(new_n834), .A3(new_n836), .ZN(G1344gat));
  NAND3_X1  g636(.A1(new_n816), .A2(new_n823), .A3(new_n631), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n839), .A3(new_n314), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n781), .A2(new_n627), .A3(new_n769), .A4(new_n770), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n244), .B1(new_n820), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n815), .B(new_n515), .C1(new_n844), .C2(new_n785), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n631), .B(new_n845), .C1(new_n814), .C2(new_n815), .ZN(new_n846));
  OAI21_X1  g645(.A(G148gat), .B1(new_n846), .B2(new_n818), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT59), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n838), .A2(KEYINPUT121), .A3(new_n839), .A4(new_n314), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n842), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR4_X1   g649(.A1(new_n826), .A2(new_n314), .A3(new_n708), .A4(new_n818), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT120), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1345gat));
  AND2_X1   g652(.A1(new_n816), .A2(new_n823), .ZN(new_n854));
  INV_X1    g653(.A(G155gat), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n667), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n814), .A2(new_n244), .A3(new_n817), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n814), .A2(KEYINPUT122), .A3(new_n244), .A4(new_n817), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n855), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT123), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n857), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1346gat));
  NAND2_X1  g666(.A1(new_n316), .A2(new_n317), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n287), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n814), .A2(new_n664), .A3(new_n817), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n854), .A2(new_n869), .B1(new_n868), .B2(new_n870), .ZN(G1347gat));
  AOI21_X1  g670(.A(new_n526), .B1(new_n784), .B2(new_n786), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n532), .A3(new_n790), .ZN(new_n873));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873), .B2(new_n615), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n872), .A2(new_n589), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n532), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n614), .A2(new_n355), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(G1348gat));
  NOR3_X1   g677(.A1(new_n873), .A2(new_n356), .A3(new_n708), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n875), .A2(new_n631), .A3(new_n532), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n356), .ZN(G1349gat));
  OAI21_X1  g680(.A(G183gat), .B1(new_n873), .B2(new_n667), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n875), .A2(new_n370), .A3(new_n532), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n653), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g684(.A(G190gat), .B1(new_n873), .B2(new_n287), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n876), .A2(new_n287), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT124), .B1(new_n890), .B2(new_n369), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892));
  INV_X1    g691(.A(new_n369), .ZN(new_n893));
  NOR4_X1   g692(.A1(new_n876), .A2(new_n892), .A3(new_n893), .A4(new_n287), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n888), .B(new_n889), .C1(new_n891), .C2(new_n894), .ZN(G1351gat));
  NAND3_X1  g694(.A1(new_n583), .A2(new_n485), .A3(new_n532), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n897), .B(new_n845), .C1(new_n814), .C2(new_n815), .ZN(new_n898));
  OAI21_X1  g697(.A(G197gat), .B1(new_n898), .B2(new_n615), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n826), .A2(new_n896), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n607), .A3(new_n614), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1352gat));
  NOR4_X1   g701(.A1(new_n826), .A2(G204gat), .A3(new_n708), .A4(new_n896), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT62), .ZN(new_n904));
  OAI21_X1  g703(.A(G204gat), .B1(new_n846), .B2(new_n896), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1353gat));
  OAI21_X1  g705(.A(G211gat), .B1(new_n898), .B2(new_n653), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT63), .B(G211gat), .C1(new_n898), .C2(new_n653), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(KEYINPUT125), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n900), .A2(new_n299), .A3(new_n244), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n907), .A2(new_n913), .A3(new_n908), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(G1354gat));
  NOR3_X1   g714(.A1(new_n826), .A2(new_n287), .A3(new_n896), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n287), .A2(new_n300), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT126), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n916), .A2(G218gat), .B1(new_n898), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT127), .Z(G1355gat));
endmodule


