

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(n727), .ZN(n523) );
  OR2_X1 U556 ( .A1(n965), .A2(n700), .ZN(n701) );
  NAND2_X1 U557 ( .A1(n767), .A2(n766), .ZN(n806) );
  AND2_X1 U558 ( .A1(n765), .A2(n528), .ZN(n766) );
  NOR2_X1 U559 ( .A1(G651), .A2(n654), .ZN(n656) );
  AND2_X1 U560 ( .A1(n525), .A2(n805), .ZN(n524) );
  XOR2_X1 U561 ( .A(KEYINPUT98), .B(n803), .Z(n525) );
  AND2_X1 U562 ( .A1(n551), .A2(n550), .ZN(n526) );
  XOR2_X1 U563 ( .A(KEYINPUT14), .B(n559), .Z(n527) );
  OR2_X1 U564 ( .A1(n764), .A2(n763), .ZN(n528) );
  AND2_X1 U565 ( .A1(n711), .A2(n710), .ZN(n712) );
  INV_X1 U566 ( .A(KEYINPUT103), .ZN(n741) );
  NAND2_X1 U567 ( .A1(n769), .A2(n690), .ZN(n727) );
  AND2_X1 U568 ( .A1(n531), .A2(G2104), .ZN(n873) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n558), .Z(n660) );
  AND2_X1 U570 ( .A1(n872), .A2(G138), .ZN(n554) );
  NAND2_X1 U571 ( .A1(n568), .A2(n567), .ZN(n980) );
  NOR2_X1 U572 ( .A1(n539), .A2(n538), .ZN(G160) );
  INV_X1 U573 ( .A(KEYINPUT23), .ZN(n530) );
  INV_X1 U574 ( .A(G2105), .ZN(n531) );
  NAND2_X1 U575 ( .A1(n873), .A2(G101), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n530), .B(n529), .ZN(n533) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n531), .ZN(n876) );
  NAND2_X1 U578 ( .A1(n876), .A2(G125), .ZN(n532) );
  NAND2_X1 U579 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U580 ( .A(KEYINPUT64), .B(n534), .ZN(n539) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n535) );
  XOR2_X2 U582 ( .A(KEYINPUT17), .B(n535), .Z(n872) );
  NAND2_X1 U583 ( .A1(G137), .A2(n872), .ZN(n537) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n877) );
  NAND2_X1 U585 ( .A1(G113), .A2(n877), .ZN(n536) );
  NAND2_X1 U586 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U587 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U588 ( .A1(G135), .A2(n872), .ZN(n540) );
  XNOR2_X1 U589 ( .A(n540), .B(KEYINPUT76), .ZN(n548) );
  NAND2_X1 U590 ( .A1(n876), .A2(G123), .ZN(n541) );
  XNOR2_X1 U591 ( .A(n541), .B(KEYINPUT18), .ZN(n543) );
  NAND2_X1 U592 ( .A1(G111), .A2(n877), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U594 ( .A1(G99), .A2(n873), .ZN(n544) );
  XNOR2_X1 U595 ( .A(KEYINPUT77), .B(n544), .ZN(n545) );
  NOR2_X1 U596 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n548), .A2(n547), .ZN(n999) );
  XNOR2_X1 U598 ( .A(G2096), .B(n999), .ZN(n549) );
  OR2_X1 U599 ( .A1(G2100), .A2(n549), .ZN(G156) );
  INV_X1 U600 ( .A(G57), .ZN(G237) );
  NAND2_X1 U601 ( .A1(G114), .A2(n877), .ZN(n551) );
  NAND2_X1 U602 ( .A1(G102), .A2(n873), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G126), .A2(n876), .ZN(n552) );
  NAND2_X1 U604 ( .A1(n526), .A2(n552), .ZN(n553) );
  NOR2_X1 U605 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U606 ( .A(KEYINPUT89), .B(n555), .Z(G164) );
  NAND2_X1 U607 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U608 ( .A(n556), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U609 ( .A(G223), .ZN(n823) );
  NAND2_X1 U610 ( .A1(n823), .A2(G567), .ZN(n557) );
  XOR2_X1 U611 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  INV_X1 U612 ( .A(G651), .ZN(n561) );
  NOR2_X1 U613 ( .A1(G543), .A2(n561), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n660), .A2(G56), .ZN(n559) );
  NOR2_X1 U615 ( .A1(G543), .A2(G651), .ZN(n644) );
  NAND2_X1 U616 ( .A1(n644), .A2(G81), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n560), .B(KEYINPUT12), .ZN(n563) );
  XOR2_X1 U618 ( .A(G543), .B(KEYINPUT0), .Z(n654) );
  NOR2_X1 U619 ( .A1(n654), .A2(n561), .ZN(n645) );
  NAND2_X1 U620 ( .A1(G68), .A2(n645), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT13), .B(n564), .Z(n565) );
  NOR2_X1 U623 ( .A1(n527), .A2(n565), .ZN(n566) );
  XNOR2_X1 U624 ( .A(n566), .B(KEYINPUT70), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G43), .A2(n656), .ZN(n567) );
  INV_X1 U626 ( .A(G860), .ZN(n610) );
  OR2_X1 U627 ( .A1(n980), .A2(n610), .ZN(G153) );
  NAND2_X1 U628 ( .A1(G52), .A2(n656), .ZN(n570) );
  NAND2_X1 U629 ( .A1(G64), .A2(n660), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U631 ( .A(KEYINPUT67), .B(n571), .Z(n576) );
  NAND2_X1 U632 ( .A1(G90), .A2(n644), .ZN(n573) );
  NAND2_X1 U633 ( .A1(G77), .A2(n645), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT9), .B(n574), .Z(n575) );
  NOR2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U637 ( .A(KEYINPUT68), .B(n577), .ZN(G171) );
  XNOR2_X1 U638 ( .A(KEYINPUT71), .B(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n578) );
  XNOR2_X1 U640 ( .A(n578), .B(KEYINPUT72), .ZN(n589) );
  INV_X1 U641 ( .A(G868), .ZN(n672) );
  NAND2_X1 U642 ( .A1(n644), .A2(G92), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT73), .B(n579), .Z(n581) );
  NAND2_X1 U644 ( .A1(n660), .A2(G66), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT74), .B(n582), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G54), .A2(n656), .ZN(n584) );
  NAND2_X1 U648 ( .A1(G79), .A2(n645), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT15), .B(n587), .Z(n965) );
  INV_X1 U652 ( .A(n965), .ZN(n832) );
  NAND2_X1 U653 ( .A1(n672), .A2(n832), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G91), .A2(n644), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G78), .A2(n645), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G65), .A2(n660), .ZN(n592) );
  XNOR2_X1 U659 ( .A(KEYINPUT69), .B(n592), .ZN(n593) );
  NOR2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U661 ( .A1(n656), .A2(G53), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(G299) );
  NAND2_X1 U663 ( .A1(n644), .A2(G89), .ZN(n597) );
  XNOR2_X1 U664 ( .A(n597), .B(KEYINPUT4), .ZN(n599) );
  NAND2_X1 U665 ( .A1(G76), .A2(n645), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U667 ( .A(KEYINPUT5), .B(n600), .ZN(n606) );
  NAND2_X1 U668 ( .A1(n660), .A2(G63), .ZN(n601) );
  XOR2_X1 U669 ( .A(KEYINPUT75), .B(n601), .Z(n603) );
  NAND2_X1 U670 ( .A1(n656), .A2(G51), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U672 ( .A(KEYINPUT6), .B(n604), .Z(n605) );
  NAND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U674 ( .A(KEYINPUT7), .B(n607), .ZN(G168) );
  XOR2_X1 U675 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U677 ( .A1(G286), .A2(n672), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n611), .A2(n965), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n980), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G868), .A2(n965), .ZN(n613) );
  NOR2_X1 U684 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U686 ( .A1(n660), .A2(G67), .ZN(n616) );
  XOR2_X1 U687 ( .A(KEYINPUT79), .B(n616), .Z(n618) );
  NAND2_X1 U688 ( .A1(n656), .A2(G55), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U690 ( .A(KEYINPUT80), .B(n619), .ZN(n624) );
  NAND2_X1 U691 ( .A1(n644), .A2(G93), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n620), .B(KEYINPUT78), .ZN(n622) );
  NAND2_X1 U693 ( .A1(G80), .A2(n645), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  OR2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n671) );
  NAND2_X1 U696 ( .A1(n965), .A2(G559), .ZN(n669) );
  XNOR2_X1 U697 ( .A(n980), .B(n669), .ZN(n625) );
  NOR2_X1 U698 ( .A1(G860), .A2(n625), .ZN(n626) );
  XOR2_X1 U699 ( .A(KEYINPUT81), .B(n626), .Z(n627) );
  XOR2_X1 U700 ( .A(n671), .B(n627), .Z(G145) );
  NAND2_X1 U701 ( .A1(G86), .A2(n644), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G61), .A2(n660), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n645), .A2(G73), .ZN(n630) );
  XOR2_X1 U705 ( .A(KEYINPUT2), .B(n630), .Z(n631) );
  NOR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U707 ( .A(KEYINPUT83), .B(n633), .Z(n635) );
  NAND2_X1 U708 ( .A1(n656), .A2(G48), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G50), .A2(n656), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT84), .ZN(n643) );
  NAND2_X1 U712 ( .A1(G88), .A2(n644), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G62), .A2(n660), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G75), .A2(n645), .ZN(n639) );
  XNOR2_X1 U716 ( .A(KEYINPUT85), .B(n639), .ZN(n640) );
  NOR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(G303) );
  INV_X1 U719 ( .A(G303), .ZN(G166) );
  NAND2_X1 U720 ( .A1(n660), .A2(G60), .ZN(n652) );
  NAND2_X1 U721 ( .A1(G85), .A2(n644), .ZN(n647) );
  NAND2_X1 U722 ( .A1(G72), .A2(n645), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G47), .A2(n656), .ZN(n648) );
  XNOR2_X1 U725 ( .A(KEYINPUT65), .B(n648), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT66), .ZN(G290) );
  NAND2_X1 U729 ( .A1(G87), .A2(n654), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n655), .B(KEYINPUT82), .ZN(n662) );
  NAND2_X1 U731 ( .A1(G49), .A2(n656), .ZN(n658) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n662), .A2(n661), .ZN(G288) );
  XOR2_X1 U736 ( .A(G305), .B(n671), .Z(n664) );
  INV_X1 U737 ( .A(G299), .ZN(n968) );
  XNOR2_X1 U738 ( .A(G166), .B(n968), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(n980), .ZN(n668) );
  XNOR2_X1 U741 ( .A(G290), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n666), .B(G288), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n668), .B(n667), .ZN(n831) );
  XNOR2_X1 U744 ( .A(n669), .B(n831), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U747 ( .A1(n674), .A2(n673), .ZN(G295) );
  XOR2_X1 U748 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n676) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XNOR2_X1 U750 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U753 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n681) );
  NAND2_X1 U756 ( .A1(G132), .A2(G82), .ZN(n680) );
  XNOR2_X1 U757 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U758 ( .A(n682), .B(KEYINPUT87), .ZN(n683) );
  NOR2_X1 U759 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U760 ( .A1(G96), .A2(n684), .ZN(n829) );
  NAND2_X1 U761 ( .A1(n829), .A2(G2106), .ZN(n688) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U763 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U764 ( .A1(G108), .A2(n686), .ZN(n830) );
  NAND2_X1 U765 ( .A1(n830), .A2(G567), .ZN(n687) );
  NAND2_X1 U766 ( .A1(n688), .A2(n687), .ZN(n914) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U768 ( .A1(n914), .A2(n689), .ZN(n828) );
  NAND2_X1 U769 ( .A1(n828), .A2(G36), .ZN(G176) );
  XOR2_X1 U770 ( .A(KEYINPUT32), .B(KEYINPUT104), .Z(n735) );
  XNOR2_X1 U771 ( .A(G1996), .B(KEYINPUT100), .ZN(n941) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n768) );
  INV_X1 U774 ( .A(n768), .ZN(n690) );
  NAND2_X1 U775 ( .A1(n941), .A2(n523), .ZN(n691) );
  XNOR2_X1 U776 ( .A(n691), .B(KEYINPUT26), .ZN(n694) );
  AND2_X1 U777 ( .A1(n727), .A2(G1341), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n692), .A2(n980), .ZN(n693) );
  AND2_X1 U779 ( .A1(n694), .A2(n693), .ZN(n700) );
  NAND2_X1 U780 ( .A1(n700), .A2(n965), .ZN(n699) );
  INV_X1 U781 ( .A(G2067), .ZN(n945) );
  NOR2_X1 U782 ( .A1(n727), .A2(n945), .ZN(n695) );
  XNOR2_X1 U783 ( .A(n695), .B(KEYINPUT101), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n727), .A2(G1348), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U787 ( .A1(n702), .A2(n701), .ZN(n707) );
  NAND2_X1 U788 ( .A1(n523), .A2(G2072), .ZN(n703) );
  XNOR2_X1 U789 ( .A(n703), .B(KEYINPUT27), .ZN(n705) );
  INV_X1 U790 ( .A(G1956), .ZN(n920) );
  NOR2_X1 U791 ( .A1(n920), .A2(n523), .ZN(n704) );
  NOR2_X1 U792 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U793 ( .A1(n968), .A2(n708), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U795 ( .A1(n708), .A2(n968), .ZN(n709) );
  XOR2_X1 U796 ( .A(n709), .B(KEYINPUT28), .Z(n710) );
  XNOR2_X1 U797 ( .A(n712), .B(KEYINPUT29), .ZN(n716) );
  INV_X1 U798 ( .A(G1961), .ZN(n931) );
  NAND2_X1 U799 ( .A1(n727), .A2(n931), .ZN(n714) );
  XNOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .ZN(n948) );
  NAND2_X1 U801 ( .A1(n523), .A2(n948), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n718) );
  NAND2_X1 U803 ( .A1(G171), .A2(n718), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U805 ( .A(n717), .B(KEYINPUT102), .ZN(n726) );
  NOR2_X1 U806 ( .A1(G171), .A2(n718), .ZN(n723) );
  NAND2_X1 U807 ( .A1(G8), .A2(n727), .ZN(n763) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n763), .ZN(n740) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n727), .ZN(n736) );
  NOR2_X1 U810 ( .A1(n740), .A2(n736), .ZN(n719) );
  NAND2_X1 U811 ( .A1(G8), .A2(n719), .ZN(n720) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n720), .ZN(n721) );
  NOR2_X1 U813 ( .A1(G168), .A2(n721), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U815 ( .A(KEYINPUT31), .B(n724), .Z(n725) );
  NAND2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n738) );
  NAND2_X1 U817 ( .A1(G286), .A2(n738), .ZN(n732) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n763), .ZN(n729) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n730), .A2(G303), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U823 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U824 ( .A(n735), .B(n734), .ZN(n744) );
  NAND2_X1 U825 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U827 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U828 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U829 ( .A1(n744), .A2(n743), .ZN(n758) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NOR2_X1 U831 ( .A1(n758), .A2(n971), .ZN(n747) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n745) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT105), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n750) );
  INV_X1 U835 ( .A(n763), .ZN(n748) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n972) );
  AND2_X1 U837 ( .A1(n748), .A2(n972), .ZN(n749) );
  AND2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U839 ( .A1(KEYINPUT33), .A2(n751), .ZN(n754) );
  NAND2_X1 U840 ( .A1(n971), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n752), .A2(n763), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U843 ( .A(G1981), .B(G305), .Z(n983) );
  NAND2_X1 U844 ( .A1(n755), .A2(n983), .ZN(n767) );
  NAND2_X1 U845 ( .A1(G166), .A2(G8), .ZN(n756) );
  NOR2_X1 U846 ( .A1(G2090), .A2(n756), .ZN(n757) );
  NOR2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U848 ( .A(KEYINPUT106), .B(n759), .Z(n760) );
  NAND2_X1 U849 ( .A1(n760), .A2(n763), .ZN(n765) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XNOR2_X1 U851 ( .A(n761), .B(KEYINPUT99), .ZN(n762) );
  XNOR2_X1 U852 ( .A(n762), .B(KEYINPUT24), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U854 ( .A(KEYINPUT91), .B(n770), .ZN(n801) );
  INV_X1 U855 ( .A(n801), .ZN(n818) );
  XOR2_X1 U856 ( .A(KEYINPUT37), .B(G2067), .Z(n815) );
  NAND2_X1 U857 ( .A1(G128), .A2(n876), .ZN(n772) );
  NAND2_X1 U858 ( .A1(G116), .A2(n877), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U860 ( .A(KEYINPUT35), .B(n773), .ZN(n779) );
  NAND2_X1 U861 ( .A1(G140), .A2(n872), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G104), .A2(n873), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n777) );
  XOR2_X1 U864 ( .A(KEYINPUT34), .B(KEYINPUT92), .Z(n776) );
  XNOR2_X1 U865 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n780), .ZN(n861) );
  NAND2_X1 U868 ( .A1(n815), .A2(n861), .ZN(n781) );
  XNOR2_X1 U869 ( .A(n781), .B(KEYINPUT93), .ZN(n1009) );
  NAND2_X1 U870 ( .A1(n818), .A2(n1009), .ZN(n813) );
  NAND2_X1 U871 ( .A1(G119), .A2(n876), .ZN(n783) );
  NAND2_X1 U872 ( .A1(G107), .A2(n877), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT94), .B(n784), .Z(n788) );
  NAND2_X1 U875 ( .A1(G131), .A2(n872), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G95), .A2(n873), .ZN(n785) );
  AND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n860) );
  AND2_X1 U879 ( .A1(n860), .A2(G1991), .ZN(n800) );
  NAND2_X1 U880 ( .A1(G141), .A2(n872), .ZN(n789) );
  XNOR2_X1 U881 ( .A(n789), .B(KEYINPUT96), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G105), .A2(n873), .ZN(n790) );
  XNOR2_X1 U883 ( .A(n790), .B(KEYINPUT38), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n876), .A2(G129), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G117), .A2(n877), .ZN(n793) );
  XNOR2_X1 U887 ( .A(KEYINPUT95), .B(n793), .ZN(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U890 ( .A(KEYINPUT97), .B(n798), .ZN(n856) );
  INV_X1 U891 ( .A(G1996), .ZN(n807) );
  NOR2_X1 U892 ( .A1(n856), .A2(n807), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n1007) );
  NOR2_X1 U894 ( .A1(n1007), .A2(n801), .ZN(n810) );
  INV_X1 U895 ( .A(n810), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n813), .A2(n802), .ZN(n803) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n804) );
  XNOR2_X1 U898 ( .A(n804), .B(KEYINPUT90), .ZN(n967) );
  NAND2_X1 U899 ( .A1(n967), .A2(n818), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n524), .ZN(n821) );
  AND2_X1 U901 ( .A1(n807), .A2(n856), .ZN(n1002) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n860), .ZN(n998) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n998), .A2(n808), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n1002), .A2(n811), .ZN(n812) );
  XNOR2_X1 U907 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n817) );
  NOR2_X1 U909 ( .A1(n815), .A2(n861), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n816), .B(KEYINPUT107), .ZN(n1011) );
  NAND2_X1 U911 ( .A1(n817), .A2(n1011), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U914 ( .A(KEYINPUT40), .B(n822), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n823), .ZN(G217) );
  NAND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n825) );
  INV_X1 U917 ( .A(G661), .ZN(n824) );
  NOR2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(KEYINPUT111), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(G188) );
  XOR2_X1 U922 ( .A(G96), .B(KEYINPUT112), .Z(G221) );
  INV_X1 U924 ( .A(G132), .ZN(G219) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G82), .ZN(G220) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U930 ( .A(n831), .B(G171), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n834), .B(G286), .ZN(n835) );
  NOR2_X1 U933 ( .A1(G37), .A2(n835), .ZN(G397) );
  XNOR2_X1 U934 ( .A(KEYINPUT109), .B(G2427), .ZN(n845) );
  XOR2_X1 U935 ( .A(G2443), .B(G2438), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2430), .B(G2454), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(KEYINPUT108), .B(G2435), .Z(n839) );
  XNOR2_X1 U939 ( .A(G1341), .B(G1348), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U942 ( .A(G2446), .B(G2451), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  NAND2_X1 U945 ( .A1(n846), .A2(G14), .ZN(n847) );
  XOR2_X1 U946 ( .A(KEYINPUT110), .B(n847), .Z(G401) );
  NAND2_X1 U947 ( .A1(G100), .A2(n873), .ZN(n854) );
  NAND2_X1 U948 ( .A1(G136), .A2(n872), .ZN(n849) );
  NAND2_X1 U949 ( .A1(G112), .A2(n877), .ZN(n848) );
  NAND2_X1 U950 ( .A1(n849), .A2(n848), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n876), .A2(G124), .ZN(n850) );
  XOR2_X1 U952 ( .A(KEYINPUT44), .B(n850), .Z(n851) );
  NOR2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n853) );
  NAND2_X1 U954 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n855), .B(KEYINPUT115), .ZN(G162) );
  XOR2_X1 U956 ( .A(G162), .B(n856), .Z(n858) );
  XNOR2_X1 U957 ( .A(G164), .B(G160), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n999), .B(n859), .ZN(n863) );
  XOR2_X1 U960 ( .A(n861), .B(n860), .Z(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n887) );
  NAND2_X1 U962 ( .A1(G130), .A2(n876), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G118), .A2(n877), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U965 ( .A1(G142), .A2(n872), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G106), .A2(n873), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(KEYINPUT45), .B(n868), .Z(n869) );
  NOR2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U970 ( .A(n871), .B(KEYINPUT46), .Z(n885) );
  NAND2_X1 U971 ( .A1(G139), .A2(n872), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G103), .A2(n873), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n883) );
  NAND2_X1 U974 ( .A1(G127), .A2(n876), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G115), .A2(n877), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  XNOR2_X1 U978 ( .A(KEYINPUT116), .B(n881), .ZN(n882) );
  NOR2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n992) );
  XNOR2_X1 U980 ( .A(n992), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U981 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U983 ( .A1(G37), .A2(n888), .ZN(G395) );
  XNOR2_X1 U984 ( .A(G1986), .B(KEYINPUT41), .ZN(n898) );
  XOR2_X1 U985 ( .A(G1976), .B(G1956), .Z(n890) );
  XNOR2_X1 U986 ( .A(G1971), .B(G1961), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n894) );
  XOR2_X1 U988 ( .A(G1981), .B(G1966), .Z(n892) );
  XNOR2_X1 U989 ( .A(G1996), .B(G1991), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U991 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U992 ( .A(KEYINPUT114), .B(G2474), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(G229) );
  XOR2_X1 U995 ( .A(KEYINPUT113), .B(G2072), .Z(n900) );
  XNOR2_X1 U996 ( .A(G2084), .B(G2078), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(G2100), .Z(n903) );
  XNOR2_X1 U999 ( .A(G2067), .B(G2090), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1001 ( .A(G2096), .B(KEYINPUT43), .Z(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT42), .B(G2678), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(G227) );
  NOR2_X1 U1005 ( .A1(n914), .A2(G401), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT117), .B(n908), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n909), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1010 ( .A1(G395), .A2(n911), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n914), .ZN(G319) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1015 ( .A(G1976), .B(G23), .Z(n916) );
  XOR2_X1 U1016 ( .A(G1971), .B(G22), .Z(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(G24), .B(G1986), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1020 ( .A(KEYINPUT58), .B(n919), .Z(n937) );
  XOR2_X1 U1021 ( .A(G1966), .B(G21), .Z(n930) );
  XNOR2_X1 U1022 ( .A(G20), .B(n920), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(G1341), .B(G19), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(G6), .B(G1981), .ZN(n921) );
  NOR2_X1 U1025 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1027 ( .A(KEYINPUT59), .B(G1348), .Z(n925) );
  XNOR2_X1 U1028 ( .A(G4), .B(n925), .ZN(n926) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1030 ( .A(KEYINPUT60), .B(n928), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n934) );
  XOR2_X1 U1032 ( .A(KEYINPUT126), .B(n931), .Z(n932) );
  XNOR2_X1 U1033 ( .A(G5), .B(n932), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(KEYINPUT127), .B(n935), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1037 ( .A(KEYINPUT61), .B(n938), .Z(n939) );
  NOR2_X1 U1038 ( .A1(G16), .A2(n939), .ZN(n964) );
  XOR2_X1 U1039 ( .A(G2072), .B(G33), .Z(n940) );
  NAND2_X1 U1040 ( .A1(n940), .A2(G28), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G32), .B(n941), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(KEYINPUT124), .B(n942), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n952) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n947) );
  XNOR2_X1 U1045 ( .A(n945), .B(G26), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1047 ( .A(G27), .B(n948), .Z(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(n953), .B(KEYINPUT53), .ZN(n956) );
  XOR2_X1 U1051 ( .A(G2084), .B(KEYINPUT54), .Z(n954) );
  XNOR2_X1 U1052 ( .A(G34), .B(n954), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G35), .B(G2090), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(n959), .ZN(n961) );
  INV_X1 U1057 ( .A(G29), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n962), .A2(G11), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n991) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n989) );
  XOR2_X1 U1062 ( .A(G1348), .B(n965), .Z(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n979) );
  XNOR2_X1 U1064 ( .A(n968), .B(G1956), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(n969), .B(KEYINPUT125), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G166), .B(G1971), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G171), .B(G1961), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n980), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G168), .B(G1966), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n985), .B(KEYINPUT57), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n1024) );
  INV_X1 U1081 ( .A(KEYINPUT55), .ZN(n1020) );
  XOR2_X1 U1082 ( .A(KEYINPUT52), .B(KEYINPUT122), .Z(n1018) );
  XNOR2_X1 U1083 ( .A(KEYINPUT120), .B(KEYINPUT50), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(G2072), .B(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(G164), .B(G2078), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n996), .B(n995), .ZN(n1015) );
  XOR2_X1 U1088 ( .A(G160), .B(G2084), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1003), .B(KEYINPUT51), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(n1010), .B(KEYINPUT118), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT119), .B(n1013), .Z(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(n1016), .B(KEYINPUT121), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1104 ( .A1(n1021), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(n1022), .B(KEYINPUT123), .ZN(n1023) );
  NOR2_X1 U1106 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1107 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

