//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n188), .A2(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(G137), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT65), .B(new_n196), .C1(new_n197), .C2(G137), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n202), .A2(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n207), .A2(new_n208), .A3(new_n200), .A4(new_n204), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n195), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(G134), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n203), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G131), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n188), .A2(new_n190), .A3(new_n214), .A4(G128), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n209), .A2(new_n213), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n210), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(G116), .B(G119), .Z(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT2), .B(G113), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  NOR4_X1   g041(.A1(new_n210), .A2(new_n220), .A3(new_n227), .A4(new_n224), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n226), .A2(new_n228), .B1(new_n225), .B2(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT28), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n206), .A2(new_n209), .ZN(new_n231));
  INV_X1    g045(.A(new_n195), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n209), .A2(new_n213), .A3(new_n219), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n225), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT28), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n238));
  NOR2_X1   g052(.A1(G237), .A2(G953), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G210), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n238), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G101), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n230), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n204), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT65), .B1(new_n211), .B2(new_n196), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n208), .B1(new_n247), .B2(new_n207), .ZN(new_n248));
  INV_X1    g062(.A(new_n209), .ZN(new_n249));
  OAI211_X1 g063(.A(KEYINPUT64), .B(new_n232), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n209), .A2(KEYINPUT64), .A3(new_n219), .A4(new_n213), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(KEYINPUT64), .B(KEYINPUT30), .C1(new_n210), .C2(new_n220), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n224), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n235), .A2(new_n227), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n221), .A2(KEYINPUT66), .A3(new_n225), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n243), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT29), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n244), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  INV_X1    g078(.A(new_n237), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n229), .B2(KEYINPUT28), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT29), .A3(new_n243), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G472), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n256), .A2(new_n259), .A3(new_n243), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT31), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n224), .A2(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n243), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n271), .B(new_n274), .C1(new_n266), .C2(new_n243), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT32), .ZN(new_n276));
  NOR2_X1   g090(.A1(G472), .A2(G902), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n275), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n269), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n269), .B(KEYINPUT68), .C1(new_n278), .C2(new_n279), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(G234), .B2(new_n264), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT23), .B1(new_n216), .B2(G119), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n288), .B(KEYINPUT69), .ZN(new_n289));
  INV_X1    g103(.A(G119), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(G128), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT70), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G119), .B(G128), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT24), .B(G110), .Z(new_n297));
  OAI22_X1  g111(.A1(new_n295), .A2(G110), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(G140), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n301), .B1(new_n305), .B2(G140), .ZN(new_n306));
  INV_X1    g120(.A(G140), .ZN(new_n307));
  AOI211_X1 g121(.A(new_n299), .B(new_n307), .C1(new_n302), .C2(new_n304), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT16), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT16), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n302), .A2(new_n304), .A3(new_n310), .A4(new_n307), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n311), .A2(new_n312), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n309), .A2(G146), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G125), .B(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n187), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n298), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n309), .A2(new_n316), .A3(new_n314), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n187), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n317), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n295), .A2(new_n324), .A3(G110), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n289), .A2(new_n292), .B1(KEYINPUT23), .B2(new_n291), .ZN(new_n326));
  INV_X1    g140(.A(G110), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT71), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n297), .A2(new_n296), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n323), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n322), .A2(new_n317), .B1(new_n296), .B2(new_n297), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n330), .B1(new_n334), .B2(new_n329), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n320), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT22), .B(G137), .Z(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT76), .ZN(new_n338));
  INV_X1    g152(.A(G953), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n339), .A2(G221), .A3(G234), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT73), .B1(new_n307), .B2(G125), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT72), .B(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(new_n307), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n303), .A2(G125), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n347));
  OAI211_X1 g161(.A(KEYINPUT73), .B(G140), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n313), .B1(new_n349), .B2(KEYINPUT16), .ZN(new_n350));
  AOI21_X1  g164(.A(G146), .B1(new_n350), .B2(new_n316), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n310), .B1(new_n345), .B2(new_n348), .ZN(new_n352));
  NOR4_X1   g166(.A1(new_n352), .A2(new_n313), .A3(new_n187), .A4(new_n315), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n331), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n325), .A2(new_n328), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT75), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n332), .ZN(new_n357));
  INV_X1    g171(.A(new_n341), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n320), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n342), .A2(new_n264), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n342), .A2(KEYINPUT25), .A3(new_n264), .A4(new_n359), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n287), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n360), .A2(new_n286), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n284), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G113), .B(G122), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT17), .ZN(new_n372));
  INV_X1    g186(.A(G237), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n339), .A3(G214), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n189), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n239), .B(G214), .C1(KEYINPUT82), .C2(G143), .ZN(new_n377));
  AOI211_X1 g191(.A(new_n372), .B(new_n208), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(new_n208), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n380), .B2(new_n372), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n322), .A3(new_n317), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n345), .A2(G146), .A3(new_n348), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n383), .A2(new_n384), .A3(new_n319), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n383), .B2(new_n319), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n379), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n371), .B1(new_n382), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(G902), .B1(new_n392), .B2(KEYINPUT87), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n382), .A2(new_n371), .A3(new_n391), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT87), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n393), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT86), .B(G475), .Z(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT9), .B(G234), .Z(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n402), .A2(new_n285), .A3(G953), .ZN(new_n403));
  XNOR2_X1  g217(.A(G116), .B(G122), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G116), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT14), .A3(G122), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(G107), .A3(new_n408), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n409), .A2(KEYINPUT88), .ZN(new_n410));
  XOR2_X1   g224(.A(G128), .B(G143), .Z(new_n411));
  OR2_X1    g225(.A1(new_n411), .A2(G134), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(G134), .ZN(new_n413));
  INV_X1    g227(.A(G107), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(new_n404), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(KEYINPUT88), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n404), .B(new_n414), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT13), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n189), .A3(G128), .ZN(new_n420));
  OAI211_X1 g234(.A(G134), .B(new_n420), .C1(new_n411), .C2(new_n419), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n421), .A3(new_n412), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n403), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n417), .A2(new_n422), .A3(new_n403), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G478), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n427), .A2(KEYINPUT15), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n264), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n428), .B1(new_n426), .B2(new_n264), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT84), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n345), .B2(new_n348), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n318), .A2(KEYINPUT19), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n434), .B(new_n187), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n317), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n187), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n380), .B1(new_n440), .B2(KEYINPUT84), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n385), .A2(new_n387), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n439), .A2(new_n441), .B1(new_n442), .B2(new_n390), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n433), .B1(new_n443), .B2(new_n371), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(KEYINPUT84), .ZN(new_n445));
  INV_X1    g259(.A(new_n380), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n445), .A2(new_n317), .A3(new_n446), .A4(new_n438), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n391), .ZN(new_n448));
  INV_X1    g262(.A(new_n371), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(KEYINPUT85), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n394), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n452));
  NOR2_X1   g266(.A1(G475), .A2(G902), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n400), .B(new_n432), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n339), .A2(G952), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(G234), .B2(G237), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XOR2_X1   g273(.A(KEYINPUT21), .B(G898), .Z(new_n460));
  NAND2_X1  g274(.A1(G234), .A2(G237), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(G902), .A3(G953), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT89), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n396), .A2(new_n392), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n398), .B1(new_n466), .B2(new_n393), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n451), .A2(new_n453), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT20), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n463), .A4(new_n432), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT5), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n290), .A3(G116), .ZN(new_n476));
  OAI211_X1 g290(.A(G113), .B(new_n476), .C1(new_n222), .C2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n222), .B2(new_n223), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT3), .B1(new_n370), .B2(G107), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n414), .A3(G104), .ZN(new_n481));
  INV_X1    g295(.A(G101), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n370), .A2(G107), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n479), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n414), .A2(G104), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n370), .A2(G107), .ZN(new_n486));
  OAI21_X1  g300(.A(G101), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n478), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n478), .A2(new_n488), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G122), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT8), .Z(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT81), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n195), .A2(new_n344), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n339), .A2(G224), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n188), .A2(new_n190), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n214), .B1(G143), .B2(new_n187), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n216), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n215), .A3(new_n305), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n497), .A2(KEYINPUT7), .A3(new_n498), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n502), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n505));
  INV_X1    g319(.A(new_n498), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n495), .A2(new_n496), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G101), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT4), .A3(new_n484), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n512), .A3(G101), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n224), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n489), .A2(new_n492), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n493), .B1(new_n489), .B2(new_n490), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n507), .A2(new_n503), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT81), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n508), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n489), .A2(new_n514), .ZN(new_n520));
  INV_X1    g334(.A(new_n492), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(KEYINPUT6), .A3(new_n515), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n504), .B(new_n506), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n525), .A3(new_n521), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n519), .A2(new_n264), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G210), .B1(G237), .B2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n519), .A2(new_n527), .A3(new_n264), .A4(new_n529), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G214), .B1(G237), .B2(G902), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT10), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT78), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT78), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n188), .A2(new_n539), .A3(KEYINPUT1), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(G128), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n499), .A2(new_n216), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n541), .A2(new_n499), .B1(new_n542), .B2(new_n214), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n536), .B1(new_n543), .B2(new_n488), .ZN(new_n544));
  INV_X1    g358(.A(new_n231), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n232), .A2(new_n511), .A3(new_n513), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n484), .A2(new_n487), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT10), .A3(new_n219), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(new_n499), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n488), .B1(new_n550), .B2(new_n215), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n547), .A2(new_n219), .ZN(new_n552));
  OAI211_X1 g366(.A(KEYINPUT12), .B(new_n231), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n488), .A2(new_n501), .A3(new_n215), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n543), .B2(new_n488), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT12), .B1(new_n556), .B2(new_n231), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n549), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G140), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT77), .ZN(new_n560));
  INV_X1    g374(.A(G227), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G953), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n560), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n549), .A2(new_n563), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n231), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT79), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n566), .B1(new_n554), .B2(new_n557), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n549), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n564), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n571), .A3(new_n264), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT79), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n558), .A2(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n578), .B(G469), .C1(new_n579), .C2(G902), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n572), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G221), .B1(new_n402), .B2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT80), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT80), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n535), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n368), .A2(new_n474), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  NAND2_X1  g403(.A1(new_n271), .A2(new_n274), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n243), .B1(new_n230), .B2(new_n237), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n264), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n277), .B1(new_n590), .B2(new_n591), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n366), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n534), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n531), .B2(new_n532), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n463), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n426), .A2(KEYINPUT33), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n426), .A2(KEYINPUT33), .ZN(new_n602));
  OAI211_X1 g416(.A(G478), .B(new_n264), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n426), .A2(new_n264), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n604), .A2(KEYINPUT90), .A3(new_n427), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT90), .B1(new_n604), .B2(new_n427), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n600), .A2(new_n471), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n584), .A2(new_n586), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n597), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT34), .B(G104), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  NOR2_X1   g429(.A1(new_n597), .A2(new_n612), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT91), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n454), .B2(new_n455), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n469), .A2(KEYINPUT91), .A3(new_n470), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n432), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n400), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n620), .A2(new_n600), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  AOI21_X1  g440(.A(new_n358), .B1(new_n357), .B2(new_n320), .ZN(new_n627));
  INV_X1    g441(.A(new_n320), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n628), .B(new_n341), .C1(new_n356), .C2(new_n332), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT25), .B1(new_n630), .B2(new_n264), .ZN(new_n631));
  INV_X1    g445(.A(new_n363), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n286), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n287), .A2(new_n264), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT92), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n357), .B2(new_n320), .ZN(new_n636));
  AOI211_X1 g450(.A(KEYINPUT92), .B(new_n628), .C1(new_n356), .C2(new_n332), .ZN(new_n637));
  OAI22_X1  g451(.A1(new_n636), .A2(new_n637), .B1(KEYINPUT36), .B2(new_n341), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n336), .A2(KEYINPUT92), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n341), .A2(KEYINPUT36), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n357), .A2(new_n635), .A3(new_n320), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n634), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n595), .B1(new_n633), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n587), .A2(new_n645), .A3(new_n474), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT37), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n327), .ZN(G12));
  INV_X1    g462(.A(new_n283), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n594), .A2(KEYINPUT32), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT68), .B1(new_n652), .B2(new_n269), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n633), .A2(new_n644), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n462), .A2(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n459), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n620), .A2(new_n622), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n654), .A2(new_n587), .A3(new_n655), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XNOR2_X1  g475(.A(new_n657), .B(KEYINPUT93), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT39), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n611), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT40), .Z(new_n665));
  INV_X1    g479(.A(new_n652), .ZN(new_n666));
  INV_X1    g480(.A(G472), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n272), .A2(new_n261), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n221), .A2(new_n225), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n257), .B2(new_n258), .ZN(new_n671));
  AOI21_X1  g485(.A(G902), .B1(new_n671), .B2(new_n261), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n667), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n533), .B(KEYINPUT38), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n400), .B1(new_n454), .B2(new_n455), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n621), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n655), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n665), .A2(new_n534), .A3(new_n676), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  AND3_X1   g495(.A1(new_n282), .A2(new_n283), .A3(new_n655), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n677), .A2(new_n607), .A3(new_n657), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT94), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT94), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n677), .A2(new_n607), .A3(new_n685), .A4(new_n657), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n682), .A2(new_n587), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT95), .B(G146), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G48));
  NAND2_X1  g504(.A1(new_n576), .A2(new_n264), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n582), .A3(new_n577), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n282), .A2(new_n366), .A3(new_n283), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n609), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n623), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  AND3_X1   g514(.A1(new_n694), .A2(KEYINPUT96), .A3(new_n599), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT96), .B1(new_n694), .B2(new_n599), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n682), .A2(KEYINPUT97), .A3(new_n474), .A4(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT97), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n474), .A2(new_n282), .A3(new_n283), .A4(new_n655), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n701), .A2(new_n702), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT98), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NAND2_X1  g525(.A1(new_n694), .A2(new_n463), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT99), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n266), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n713), .B(new_n237), .C1(new_n671), .C2(new_n236), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n261), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n271), .B(new_n274), .C1(new_n714), .C2(new_n716), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n717), .A2(new_n277), .B1(new_n592), .B2(G472), .ZN(new_n718));
  INV_X1    g532(.A(new_n365), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n633), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT100), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT100), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n633), .A2(new_n718), .A3(new_n722), .A4(new_n719), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n712), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n678), .A2(new_n535), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(G122), .Z(G24));
  AOI21_X1  g541(.A(KEYINPUT101), .B1(new_n655), .B2(new_n718), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT101), .B(new_n718), .C1(new_n364), .C2(new_n643), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n687), .B(new_n703), .C1(new_n728), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NOR2_X1   g546(.A1(new_n533), .A2(new_n598), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(G469), .B1(new_n579), .B2(G902), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n577), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n582), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n280), .A2(new_n633), .A3(new_n719), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n687), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AND4_X1   g554(.A1(new_n282), .A2(new_n738), .A3(new_n283), .A4(new_n366), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n684), .A2(new_n686), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n740), .A2(KEYINPUT42), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT102), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n208), .ZN(G33));
  NAND2_X1  g560(.A1(new_n741), .A2(new_n659), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  OAI21_X1  g562(.A(G469), .B1(new_n579), .B2(KEYINPUT45), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT103), .Z(new_n750));
  NAND2_X1  g564(.A1(new_n579), .A2(KEYINPUT45), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT104), .Z(new_n752));
  AOI22_X1  g566(.A1(new_n750), .A2(new_n752), .B1(G469), .B2(G902), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT105), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(KEYINPUT105), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n577), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n758), .A2(new_n582), .A3(new_n663), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n471), .A2(new_n607), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n760), .B1(KEYINPUT106), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n362), .A2(new_n363), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n643), .B1(new_n767), .B2(new_n286), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n766), .A2(new_n596), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n734), .B1(new_n769), .B2(KEYINPUT44), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n759), .B(new_n770), .C1(KEYINPUT44), .C2(new_n769), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  NAND2_X1  g586(.A1(new_n758), .A2(new_n582), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n758), .A2(KEYINPUT47), .A3(new_n582), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n366), .A2(new_n734), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n284), .A3(new_n687), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(new_n582), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n367), .A2(new_n598), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(KEYINPUT107), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n675), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n674), .B1(new_n782), .B2(KEYINPUT107), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n692), .A2(new_n577), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT49), .Z(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n761), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n459), .B(new_n766), .C1(new_n723), .C2(new_n721), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n675), .A2(new_n534), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n694), .A3(new_n790), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT50), .Z(new_n792));
  INV_X1    g606(.A(new_n766), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n734), .A2(new_n459), .A3(new_n693), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n793), .B(new_n794), .C1(new_n730), .C2(new_n728), .ZN(new_n795));
  INV_X1    g609(.A(new_n674), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n796), .A2(new_n366), .A3(new_n794), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n471), .A3(new_n608), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n789), .A2(new_n733), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n692), .A2(new_n781), .A3(new_n577), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT118), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n800), .B1(new_n777), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n792), .A2(new_n795), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n775), .A2(new_n776), .A3(new_n801), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n805), .B1(new_n807), .B2(new_n800), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n792), .A2(new_n808), .A3(new_n795), .A4(new_n798), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n793), .A2(new_n739), .A3(new_n794), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT48), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n457), .B1(new_n789), .B2(new_n703), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n797), .A2(new_n677), .A3(new_n607), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT119), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n806), .A2(new_n809), .A3(new_n811), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT120), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT101), .ZN(new_n818));
  INV_X1    g632(.A(new_n718), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n818), .B1(new_n768), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n742), .B1(new_n820), .B2(new_n729), .ZN(new_n821));
  INV_X1    g635(.A(new_n737), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n432), .B(new_n657), .C1(new_n364), .C2(new_n643), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n581), .A2(new_n585), .A3(new_n582), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n585), .B1(new_n581), .B2(new_n582), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n400), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n823), .A2(new_n826), .A3(new_n620), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n821), .A2(new_n822), .B1(new_n827), .B2(new_n654), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n744), .B(new_n747), .C1(new_n828), .C2(new_n734), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n400), .B(new_n621), .C1(new_n454), .C2(new_n455), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n600), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n611), .A2(new_n366), .A3(new_n831), .A4(new_n596), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n646), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT109), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n616), .A2(new_n609), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT109), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n646), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n834), .A2(new_n588), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT110), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n613), .B1(new_n833), .B2(KEYINPUT109), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT110), .A3(new_n588), .A4(new_n837), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n829), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n724), .A2(new_n725), .B1(new_n695), .B2(new_n609), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n709), .A2(new_n699), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT108), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT108), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n709), .A2(new_n844), .A3(new_n847), .A4(new_n699), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n737), .B1(new_n850), .B2(new_n658), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n657), .A2(KEYINPUT112), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n633), .A2(new_n851), .A3(new_n644), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n768), .A2(KEYINPUT113), .A3(new_n852), .A4(new_n851), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n674), .A4(new_n725), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n688), .A2(new_n731), .A3(new_n660), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n843), .A2(new_n849), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT115), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n861), .A2(KEYINPUT115), .A3(new_n862), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n731), .A2(new_n660), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT111), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n857), .A2(KEYINPUT52), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n731), .A2(new_n660), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n866), .A2(new_n688), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n858), .A2(new_n859), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(KEYINPUT114), .A3(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n876), .A2(new_n843), .A3(new_n849), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n863), .B(new_n864), .C1(new_n877), .C2(KEYINPUT53), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n878), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n861), .A2(new_n862), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n845), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n876), .A2(KEYINPUT53), .A3(new_n843), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n861), .A2(KEYINPUT117), .A3(new_n862), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n882), .A2(new_n884), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n878), .A2(KEYINPUT54), .B1(new_n887), .B2(KEYINPUT116), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n817), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(G952), .A2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n788), .B1(new_n889), .B2(new_n890), .ZN(G75));
  AND3_X1   g705(.A1(new_n861), .A2(KEYINPUT117), .A3(new_n862), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT117), .B1(new_n861), .B2(new_n862), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n264), .B1(new_n894), .B2(new_n884), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G210), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n523), .A2(new_n526), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n524), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT55), .Z(new_n901));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(new_n897), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n898), .A2(new_n903), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n339), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  NAND2_X1  g721(.A1(G469), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT122), .Z(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT57), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n882), .A2(new_n884), .A3(new_n886), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n913), .B2(new_n887), .ZN(new_n914));
  INV_X1    g728(.A(new_n576), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT123), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n885), .B1(new_n894), .B2(new_n884), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n885), .A2(new_n882), .A3(new_n884), .A4(new_n886), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n910), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n576), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n895), .A2(new_n752), .A3(new_n750), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n906), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(new_n451), .Z(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n906), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT59), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n601), .B2(new_n602), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n913), .B2(new_n887), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n879), .B2(new_n888), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n601), .A2(new_n602), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n906), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(new_n638), .A2(new_n642), .ZN(new_n936));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n912), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n912), .A2(new_n938), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n924), .B(new_n939), .C1(new_n940), .C2(new_n630), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g756(.A(new_n339), .B1(new_n460), .B2(G224), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n840), .A2(new_n842), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n849), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n339), .ZN(new_n946));
  INV_X1    g760(.A(G898), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n899), .B1(new_n947), .B2(G953), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G69));
  NOR2_X1   g763(.A1(new_n436), .A2(new_n437), .ZN(new_n950));
  XNOR2_X1  g764(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n255), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(G900), .A2(G953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n779), .A2(new_n771), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n866), .A2(new_n688), .A3(new_n869), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n759), .A2(new_n725), .A3(new_n739), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n957), .A2(new_n744), .A3(new_n747), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n953), .B(new_n954), .C1(new_n959), .C2(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n956), .A2(new_n680), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT62), .Z(new_n962));
  INV_X1    g776(.A(new_n664), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n830), .B1(new_n471), .B2(new_n608), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n368), .A2(new_n963), .A3(new_n733), .A4(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n955), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n966), .A2(new_n339), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(new_n953), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n339), .B1(new_n953), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(G900), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n561), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n968), .B(new_n972), .Z(G72));
  OR2_X1    g787(.A1(new_n966), .A2(new_n945), .ZN(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n974), .A2(KEYINPUT127), .A3(new_n976), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n668), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n976), .B1(new_n959), .B2(new_n945), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n260), .A2(new_n243), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n906), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n878), .A2(new_n669), .A3(new_n985), .A4(new_n976), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n981), .A2(new_n984), .A3(new_n986), .ZN(G57));
endmodule


