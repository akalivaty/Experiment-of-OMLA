//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G469), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n190), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n195), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G104), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(G107), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n196), .A2(new_n199), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n195), .A2(G107), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n198), .A2(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(G101), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n210), .A3(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n212), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  OAI21_X1  g030(.A(G128), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n211), .A2(new_n216), .A3(G128), .A4(new_n213), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n206), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT10), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT83), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n196), .A2(new_n199), .A3(new_n224), .A4(new_n201), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n200), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI211_X1 g042(.A(KEYINPUT4), .B(new_n200), .C1(new_n223), .C2(new_n225), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n214), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  INV_X1    g046(.A(new_n215), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT64), .B(G146), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G143), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n231), .A2(new_n232), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n221), .B1(new_n230), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT11), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n241), .B(new_n243), .C1(new_n244), .C2(G137), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G137), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT11), .A4(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n244), .A2(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G131), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n252), .A2(new_n254), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n208), .A2(new_n210), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n215), .B1(new_n260), .B2(new_n212), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n219), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n202), .A2(new_n205), .A3(KEYINPUT84), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT84), .B1(new_n202), .B2(new_n205), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(KEYINPUT72), .B(new_n219), .C1(new_n259), .C2(new_n261), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n264), .A2(new_n267), .A3(KEYINPUT10), .A4(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n239), .A2(KEYINPUT85), .A3(new_n257), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n223), .A2(new_n225), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G101), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(new_n238), .C1(new_n226), .C2(new_n227), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n218), .A2(new_n219), .ZN(new_n275));
  INV_X1    g089(.A(new_n206), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT10), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n269), .A2(new_n274), .A3(new_n257), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n194), .B1(new_n270), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n269), .A2(new_n274), .A3(new_n279), .ZN(new_n284));
  INV_X1    g098(.A(new_n257), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT86), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n277), .B1(new_n267), .B2(new_n262), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n291), .B2(new_n257), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n285), .A3(KEYINPUT12), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n280), .A2(new_n281), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n280), .A2(new_n281), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n288), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n194), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n270), .A2(new_n282), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n288), .B1(new_n299), .B2(new_n294), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n287), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT87), .B(new_n287), .C1(new_n298), .C2(new_n300), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n189), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n283), .A2(new_n294), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n193), .B1(new_n299), .B2(new_n286), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n189), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(G469), .A2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n188), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT88), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n314), .B(new_n188), .C1(new_n305), .C2(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G110), .B(G122), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT8), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n319));
  INV_X1    g133(.A(G113), .ZN(new_n320));
  INV_X1    g134(.A(G116), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G119), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(KEYINPUT70), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G116), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(G119), .ZN(new_n328));
  INV_X1    g142(.A(new_n322), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(KEYINPUT5), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT70), .B(G116), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n322), .B1(new_n331), .B2(G119), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT69), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(new_n320), .ZN(new_n335));
  NAND3_X1  g149(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n335), .A2(new_n336), .B1(new_n334), .B2(new_n320), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n324), .A2(new_n330), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n267), .A2(new_n319), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n329), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n328), .A2(KEYINPUT71), .A3(new_n329), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(KEYINPUT5), .A3(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n344), .A2(new_n324), .B1(new_n337), .B2(new_n332), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n339), .B1(new_n345), .B2(new_n276), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n319), .B1(new_n267), .B2(new_n338), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n318), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT91), .B(G224), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n191), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT7), .ZN(new_n351));
  INV_X1    g165(.A(G125), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n235), .A2(new_n237), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n211), .A2(new_n213), .A3(new_n232), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n351), .B1(new_n355), .B2(KEYINPUT93), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n352), .B(new_n219), .C1(new_n259), .C2(new_n261), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n238), .B2(new_n352), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n356), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT94), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n271), .A2(G101), .ZN(new_n362));
  INV_X1    g176(.A(new_n227), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n337), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n328), .A2(KEYINPUT71), .A3(new_n329), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT71), .B1(new_n328), .B2(new_n329), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n332), .A2(new_n337), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n364), .A2(new_n370), .A3(new_n273), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n344), .A2(new_n324), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n369), .A3(new_n267), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n373), .A3(new_n317), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n348), .A2(new_n359), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n361), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n373), .ZN(new_n379));
  INV_X1    g193(.A(new_n317), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n374), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n358), .B(new_n350), .Z(new_n383));
  AOI21_X1  g197(.A(new_n317), .B1(new_n371), .B2(new_n373), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT89), .B(KEYINPUT6), .Z(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n382), .B(new_n383), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n377), .A2(new_n390), .A3(new_n306), .ZN(new_n391));
  OAI21_X1  g205(.A(G210), .B1(G237), .B2(G902), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT95), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n377), .A2(new_n390), .A3(new_n306), .A4(new_n392), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G214), .B1(G237), .B2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT101), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n331), .B2(G122), .ZN(new_n403));
  AND4_X1   g217(.A1(new_n402), .A2(new_n325), .A3(new_n327), .A4(G122), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT14), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n321), .A2(G122), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(KEYINPUT104), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n325), .A2(new_n327), .A3(G122), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT101), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n331), .A2(new_n402), .A3(G122), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT105), .B1(new_n412), .B2(KEYINPUT14), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n403), .A2(new_n404), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT105), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n408), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT104), .B1(new_n405), .B2(new_n407), .ZN(new_n419));
  OAI21_X1  g233(.A(G107), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G128), .B(G143), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(G134), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT102), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n414), .B2(new_n406), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n412), .A2(KEYINPUT102), .A3(new_n407), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n422), .B1(new_n426), .B2(new_n198), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n187), .A2(new_n429), .A3(G953), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n430), .B(KEYINPUT106), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT13), .ZN(new_n433));
  AOI22_X1  g247(.A1(KEYINPUT103), .A2(new_n433), .B1(new_n258), .B2(G143), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(KEYINPUT103), .B2(new_n433), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G134), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n436), .B(new_n421), .Z(new_n437));
  AND3_X1   g251(.A1(new_n424), .A2(G107), .A3(new_n425), .ZN(new_n438));
  AOI21_X1  g252(.A(G107), .B1(new_n424), .B2(new_n425), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n428), .A2(new_n432), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n432), .B1(new_n428), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n306), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n428), .A2(new_n440), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n431), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n428), .A2(new_n432), .A3(new_n440), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n445), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n306), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G475), .ZN(new_n455));
  NOR2_X1   g269(.A1(G237), .A2(G953), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(G143), .A3(G214), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G143), .B1(new_n456), .B2(G214), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT17), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n460), .A2(new_n461), .A3(new_n253), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n458), .A2(new_n459), .A3(G131), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n456), .A2(G214), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n212), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n253), .B1(new_n465), .B2(new_n457), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n462), .B1(new_n467), .B2(new_n461), .ZN(new_n468));
  INV_X1    g282(.A(G140), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n352), .A2(G140), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n472), .A2(KEYINPUT16), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n470), .A2(KEYINPUT16), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n207), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n472), .B2(KEYINPUT16), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G146), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT99), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT99), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n475), .B2(new_n477), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n468), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n470), .A2(new_n471), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT80), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n234), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(G146), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n466), .A2(KEYINPUT18), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT18), .A2(G131), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n460), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT96), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n487), .A2(new_n488), .B1(new_n460), .B2(new_n491), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT96), .A3(new_n490), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n482), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(G113), .B(G122), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n195), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n482), .A2(new_n498), .A3(new_n501), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n455), .B1(new_n505), .B2(new_n306), .ZN(new_n506));
  NOR2_X1   g320(.A1(G475), .A2(G902), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT100), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n493), .A2(new_n494), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT96), .B1(new_n496), .B2(new_n490), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT19), .B1(new_n485), .B2(new_n486), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT19), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n483), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n511), .B(new_n234), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n463), .A2(new_n466), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n477), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n486), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT80), .B1(new_n470), .B2(new_n471), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n514), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n260), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(new_n511), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n509), .A2(new_n510), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT98), .A3(new_n502), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n504), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT98), .B1(new_n524), .B2(new_n502), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n508), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT20), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n502), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT98), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n525), .A3(new_n504), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT20), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n508), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n506), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT107), .ZN(new_n537));
  INV_X1    g351(.A(G952), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G953), .ZN(new_n539));
  NAND2_X1  g353(.A1(G234), .A2(G237), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT21), .B(G898), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(G902), .A3(G953), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n454), .A2(new_n536), .A3(new_n537), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n454), .A2(new_n536), .A3(new_n545), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT107), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n401), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT81), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT22), .B(G137), .Z(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n477), .A2(new_n487), .ZN(new_n556));
  INV_X1    g370(.A(G119), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G128), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT78), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n258), .A2(G119), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G110), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n558), .A3(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(KEYINPUT23), .B2(new_n561), .ZN(new_n568));
  INV_X1    g382(.A(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n556), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n564), .A2(new_n565), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n478), .B1(new_n569), .B2(new_n568), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n555), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  OAI221_X1 g389(.A(new_n478), .B1(new_n569), .B2(new_n568), .C1(new_n564), .C2(new_n565), .ZN(new_n576));
  INV_X1    g390(.A(new_n555), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n564), .A2(new_n565), .B1(new_n569), .B2(new_n568), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n556), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n551), .B1(new_n580), .B2(G902), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n575), .A2(new_n579), .A3(new_n306), .A4(new_n550), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n581), .A2(new_n582), .B1(KEYINPUT82), .B2(KEYINPUT25), .ZN(new_n583));
  INV_X1    g397(.A(G234), .ZN(new_n584));
  OAI21_X1  g398(.A(G217), .B1(new_n584), .B2(G902), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT77), .Z(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n306), .ZN(new_n587));
  OAI22_X1  g401(.A1(new_n583), .A2(new_n586), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT30), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n245), .A2(new_n250), .A3(new_n251), .ZN(new_n590));
  AOI21_X1  g404(.A(G134), .B1(new_n247), .B2(new_n249), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n244), .A2(G137), .ZN(new_n592));
  OAI21_X1  g406(.A(G131), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n590), .A2(new_n253), .B1(new_n593), .B2(KEYINPUT68), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT68), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(G131), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n264), .A2(new_n594), .A3(new_n596), .A4(new_n268), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n238), .B1(new_n255), .B2(new_n256), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n589), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n590), .A2(new_n253), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n593), .A2(KEYINPUT68), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n600), .A2(new_n262), .A3(new_n596), .A4(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n598), .A2(new_n602), .A3(new_n589), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n370), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n456), .A2(G210), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT27), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT73), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT26), .B(G101), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n370), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n597), .A2(new_n610), .A3(new_n598), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n604), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT31), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n604), .A2(KEYINPUT31), .A3(new_n609), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n611), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n610), .B1(new_n598), .B2(new_n602), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT28), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT74), .B1(new_n617), .B2(KEYINPUT28), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT74), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT28), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n611), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n609), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n616), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT32), .ZN(new_n628));
  NOR2_X1   g442(.A1(G472), .A2(G902), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT75), .Z(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n627), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n614), .A2(new_n615), .B1(new_n624), .B2(new_n625), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT32), .B1(new_n633), .B2(new_n630), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n619), .A2(new_n620), .A3(new_n609), .A4(new_n623), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT29), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI211_X1 g452(.A(KEYINPUT76), .B(new_n609), .C1(new_n604), .C2(new_n611), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT76), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n604), .A2(new_n611), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n625), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n610), .B1(new_n597), .B2(new_n598), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT28), .B1(new_n617), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n620), .A3(new_n623), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n609), .A2(KEYINPUT29), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n306), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n588), .B1(new_n635), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n316), .A2(new_n549), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G101), .ZN(G3));
  OAI21_X1  g466(.A(G472), .B1(new_n633), .B2(G902), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n630), .B2(new_n633), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n588), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n316), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n444), .A2(G902), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT33), .B1(new_n450), .B2(KEYINPUT108), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT33), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n659), .B(new_n660), .C1(new_n448), .C2(new_n449), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n657), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n443), .A2(new_n444), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n536), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n400), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n394), .B2(new_n398), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n664), .A2(new_n545), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n656), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT34), .B(G104), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  NAND3_X1  g484(.A1(new_n379), .A2(new_n380), .A3(new_n386), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT90), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n672), .A2(new_n387), .B1(new_n374), .B2(new_n381), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n673), .B2(new_n383), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n392), .B1(new_n674), .B2(new_n377), .ZN(new_n675));
  AND4_X1   g489(.A1(new_n306), .A2(new_n377), .A3(new_n392), .A4(new_n390), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n400), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n545), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n536), .A2(new_n453), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n656), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT35), .B(G107), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  OR4_X1    g497(.A1(KEYINPUT36), .A2(new_n571), .A3(new_n574), .A4(new_n555), .ZN(new_n684));
  INV_X1    g498(.A(new_n587), .ZN(new_n685));
  OAI22_X1  g499(.A1(new_n571), .A2(new_n574), .B1(KEYINPUT36), .B2(new_n555), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n581), .A2(new_n582), .ZN(new_n688));
  NAND2_X1  g502(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n586), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n654), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n316), .A2(new_n549), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  NAND2_X1  g510(.A1(new_n635), .A2(new_n649), .ZN(new_n697));
  INV_X1    g511(.A(new_n687), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n583), .B2(new_n586), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n544), .A2(G900), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n541), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n679), .A2(new_n702), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n697), .A2(new_n666), .A3(new_n699), .A4(new_n703), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n270), .A2(new_n282), .B1(new_n293), .B2(new_n292), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n193), .B1(new_n705), .B2(new_n288), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT86), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT87), .B1(new_n709), .B2(new_n287), .ZN(new_n710));
  INV_X1    g524(.A(new_n304), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n311), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n314), .B1(new_n714), .B2(new_n188), .ZN(new_n715));
  INV_X1    g529(.A(new_n315), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n704), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  XOR2_X1   g532(.A(new_n399), .B(KEYINPUT38), .Z(new_n719));
  OAI21_X1  g533(.A(new_n625), .B1(new_n617), .B2(new_n644), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n612), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(G902), .B1(new_n721), .B2(KEYINPUT109), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(KEYINPUT109), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G472), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n635), .A2(KEYINPUT110), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT110), .B1(new_n635), .B2(new_n724), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n506), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n528), .A2(KEYINPUT20), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n534), .B1(new_n533), .B2(new_n508), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n453), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n692), .A2(new_n400), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n719), .A2(new_n727), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n701), .B(KEYINPUT39), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n316), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT40), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n736), .A2(KEYINPUT40), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n212), .ZN(G45));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n742));
  INV_X1    g556(.A(new_n657), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT108), .B1(new_n441), .B2(new_n442), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n660), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n450), .A2(KEYINPUT108), .A3(KEYINPUT33), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n663), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n731), .B(new_n701), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n742), .B1(new_n749), .B2(new_n677), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n664), .A2(KEYINPUT111), .A3(new_n666), .A4(new_n701), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n692), .B1(new_n635), .B2(new_n649), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n316), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G146), .ZN(G48));
  NAND2_X1  g569(.A1(new_n299), .A2(new_n286), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n756), .A2(new_n194), .B1(new_n283), .B2(new_n294), .ZN(new_n757));
  OAI21_X1  g571(.A(G469), .B1(new_n757), .B2(G902), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n188), .A3(new_n309), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n667), .A2(new_n650), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT41), .B(G113), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G15));
  NAND3_X1  g577(.A1(new_n680), .A2(new_n650), .A3(new_n760), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT112), .B(G116), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G18));
  NAND2_X1  g580(.A1(new_n548), .A2(new_n546), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n677), .A2(new_n759), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n752), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G119), .ZN(G21));
  INV_X1    g584(.A(new_n653), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n646), .A2(new_n625), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n616), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n772), .B1(new_n774), .B2(new_n631), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n772), .A3(new_n631), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n771), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n677), .A2(new_n732), .ZN(new_n779));
  INV_X1    g593(.A(new_n588), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n759), .A2(new_n678), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G122), .ZN(G24));
  INV_X1    g597(.A(new_n768), .ZN(new_n784));
  AOI211_X1 g598(.A(KEYINPUT113), .B(new_n630), .C1(new_n616), .C2(new_n773), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n699), .B(new_n653), .C1(new_n775), .C2(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n784), .A2(new_n786), .A3(new_n749), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n352), .ZN(G27));
  NAND4_X1  g602(.A1(new_n395), .A2(new_n400), .A3(new_n397), .A4(new_n398), .ZN(new_n789));
  INV_X1    g603(.A(new_n188), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n749), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n301), .A2(new_n189), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n311), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n650), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT42), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n789), .A2(new_n794), .A3(new_n790), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(KEYINPUT42), .A3(new_n650), .A4(new_n792), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G131), .ZN(G33));
  NAND4_X1  g616(.A1(new_n791), .A2(new_n650), .A3(new_n703), .A4(new_n795), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G134), .ZN(G36));
  AND2_X1   g618(.A1(new_n654), .A2(new_n699), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n747), .B2(new_n748), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n662), .A2(KEYINPUT116), .A3(new_n663), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n731), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(KEYINPUT43), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n536), .B(KEYINPUT117), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n662), .A2(new_n663), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n811), .A2(KEYINPUT43), .A3(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT44), .B(new_n805), .C1(new_n810), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n789), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n811), .A2(KEYINPUT43), .A3(new_n812), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(KEYINPUT43), .B2(new_n809), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT44), .B1(new_n818), .B2(new_n805), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n189), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n712), .A2(KEYINPUT114), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n305), .B2(new_n822), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n301), .A2(new_n821), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT115), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n310), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT46), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(KEYINPUT46), .A3(new_n310), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n309), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n820), .A2(new_n188), .A3(new_n834), .A4(new_n735), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  OR4_X1    g650(.A1(new_n697), .A2(new_n789), .A3(new_n780), .A4(new_n749), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT119), .Z(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(KEYINPUT118), .A2(KEYINPUT47), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n833), .A2(new_n309), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT46), .B1(new_n829), .B2(new_n310), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n188), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(KEYINPUT118), .A2(KEYINPUT47), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n844), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n834), .A2(new_n188), .A3(new_n840), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n839), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(new_n469), .ZN(G42));
  NAND2_X1  g663(.A1(new_n538), .A2(new_n191), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n761), .A2(new_n769), .A3(new_n764), .A4(new_n782), .ZN(new_n851));
  INV_X1    g665(.A(new_n786), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n799), .A2(new_n792), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(new_n803), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n731), .A2(new_n453), .A3(new_n702), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n316), .A2(new_n752), .A3(new_n815), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n801), .A2(new_n851), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n664), .B(KEYINPUT120), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n679), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n401), .A2(new_n678), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n316), .A2(new_n859), .A3(new_n655), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n651), .A3(new_n694), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n787), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n794), .A2(new_n790), .A3(new_n699), .A4(new_n702), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n865), .B(new_n779), .C1(new_n725), .C2(new_n726), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n754), .A2(new_n717), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n787), .B1(new_n316), .B2(new_n704), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(KEYINPUT52), .A3(new_n754), .A4(new_n866), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n863), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(KEYINPUT121), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n863), .B(new_n872), .C1(KEYINPUT121), .C2(KEYINPUT53), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT54), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n863), .A2(new_n872), .A3(new_n875), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n875), .B1(new_n863), .B2(new_n872), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n541), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n818), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n758), .A2(new_n309), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n789), .A2(new_n790), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n650), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT48), .Z(new_n890));
  AND2_X1   g704(.A1(new_n887), .A2(new_n884), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n725), .A2(new_n726), .A3(new_n588), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n664), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n778), .A2(new_n780), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n539), .B(new_n893), .C1(new_n896), .C2(new_n784), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n879), .A2(new_n883), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n758), .A2(new_n790), .A3(new_n309), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n845), .A2(new_n847), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n896), .A2(new_n789), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT50), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n719), .A2(new_n665), .A3(new_n760), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n896), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n905), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(KEYINPUT50), .A3(new_n885), .A4(new_n895), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n812), .A2(new_n731), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n891), .A2(new_n892), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n888), .A2(new_n852), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n903), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n903), .A2(new_n914), .A3(KEYINPUT51), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n850), .B1(new_n899), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n886), .B(KEYINPUT49), .Z(new_n921));
  AND4_X1   g735(.A1(new_n188), .A2(new_n811), .A3(new_n400), .A4(new_n812), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n719), .A2(new_n892), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(G75));
  NOR2_X1   g738(.A1(new_n881), .A2(new_n882), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(G210), .A3(G902), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n673), .B(new_n383), .Z(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n926), .B2(new_n927), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n191), .A2(G952), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G51));
  XNOR2_X1  g747(.A(new_n757), .B(KEYINPUT123), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n873), .A2(KEYINPUT53), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n863), .A2(new_n872), .A3(new_n875), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(KEYINPUT54), .A3(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n883), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n310), .B(KEYINPUT57), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n935), .A2(new_n936), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n941), .A2(new_n306), .A3(new_n829), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n932), .B1(new_n940), .B2(new_n942), .ZN(G54));
  NAND4_X1  g757(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n944));
  INV_X1    g758(.A(new_n533), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(new_n947), .A3(new_n932), .ZN(G60));
  NAND2_X1  g762(.A1(G478), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT59), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n658), .B2(new_n661), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n883), .B2(new_n937), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n880), .B1(new_n876), .B2(new_n877), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT54), .B1(new_n935), .B2(new_n936), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n658), .A2(new_n661), .ZN(new_n956));
  AOI211_X1 g770(.A(new_n932), .B(new_n952), .C1(new_n955), .C2(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT60), .Z(new_n959));
  NAND4_X1  g773(.A1(new_n925), .A2(new_n684), .A3(new_n686), .A4(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n959), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n580), .B1(new_n941), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n932), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n960), .A2(new_n962), .A3(KEYINPUT61), .A4(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G66));
  AOI21_X1  g782(.A(new_n191), .B1(new_n543), .B2(new_n349), .ZN(new_n969));
  INV_X1    g783(.A(new_n851), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n862), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n972), .B2(new_n191), .ZN(new_n973));
  INV_X1    g787(.A(G898), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n673), .B1(new_n974), .B2(G953), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  NAND2_X1  g790(.A1(G227), .A2(G900), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n650), .A2(new_n779), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n834), .A2(new_n188), .A3(new_n735), .A4(new_n978), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n754), .A2(new_n801), .A3(new_n870), .A4(new_n803), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n835), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n845), .A2(new_n847), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n838), .ZN(new_n983));
  AOI21_X1  g797(.A(G953), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n191), .A2(G900), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n599), .A2(new_n603), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n512), .A2(new_n514), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(G953), .B(new_n977), .C1(new_n988), .C2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n991), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n984), .B2(new_n987), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n977), .A2(G953), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n859), .A2(new_n650), .A3(new_n815), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(new_n736), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n835), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n835), .A2(KEYINPUT124), .A3(new_n997), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n870), .A2(new_n754), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n740), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1004), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1006), .B(KEYINPUT62), .C1(new_n738), .C2(new_n739), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n848), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(G953), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n994), .B(new_n995), .C1(new_n1009), .C2(new_n993), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n992), .A2(new_n1010), .ZN(G72));
  NAND3_X1  g825(.A1(new_n604), .A2(new_n625), .A3(new_n611), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n835), .A2(new_n979), .A3(new_n980), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1014), .A2(new_n848), .A3(new_n972), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1013), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n981), .A2(new_n983), .A3(new_n971), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1020), .A2(KEYINPUT126), .A3(new_n1017), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1012), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n641), .A2(new_n609), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1002), .A2(new_n1008), .A3(new_n971), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1023), .B1(new_n1024), .B2(new_n1017), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n642), .A2(new_n639), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1018), .B1(new_n1026), .B2(new_n612), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n878), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n963), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n1022), .A2(new_n1025), .A3(new_n1029), .ZN(G57));
endmodule


