

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U549 ( .A1(n694), .A2(n693), .ZN(n699) );
  NAND2_X1 U550 ( .A1(G8), .A2(n727), .ZN(n785) );
  XOR2_X1 U551 ( .A(KEYINPUT74), .B(n574), .Z(n990) );
  XOR2_X1 U552 ( .A(KEYINPUT73), .B(n566), .Z(n516) );
  BUF_X1 U553 ( .A(n689), .Z(n707) );
  NOR2_X1 U554 ( .A1(G1966), .A2(n785), .ZN(n739) );
  NOR2_X1 U555 ( .A1(n528), .A2(n527), .ZN(G160) );
  AND2_X1 U556 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U557 ( .A1(G113), .A2(n873), .ZN(n517) );
  XNOR2_X1 U558 ( .A(n517), .B(KEYINPUT66), .ZN(n520) );
  INV_X1 U559 ( .A(G2104), .ZN(n521) );
  NOR2_X2 U560 ( .A1(G2105), .A2(n521), .ZN(n869) );
  NAND2_X1 U561 ( .A1(G101), .A2(n869), .ZN(n518) );
  XOR2_X1 U562 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U563 ( .A1(n520), .A2(n519), .ZN(n528) );
  NAND2_X1 U564 ( .A1(n521), .A2(G2105), .ZN(n522) );
  XNOR2_X2 U565 ( .A(n522), .B(KEYINPUT65), .ZN(n874) );
  NAND2_X1 U566 ( .A1(G125), .A2(n874), .ZN(n526) );
  XNOR2_X1 U567 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n524) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U569 ( .A(n524), .B(n523), .ZN(n870) );
  NAND2_X1 U570 ( .A1(G137), .A2(n870), .ZN(n525) );
  NAND2_X1 U571 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n632) );
  NAND2_X1 U573 ( .A1(G89), .A2(n632), .ZN(n529) );
  XNOR2_X1 U574 ( .A(n529), .B(KEYINPUT76), .ZN(n530) );
  XNOR2_X1 U575 ( .A(n530), .B(KEYINPUT4), .ZN(n532) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n640) );
  INV_X1 U577 ( .A(G651), .ZN(n534) );
  NOR2_X2 U578 ( .A1(n640), .A2(n534), .ZN(n630) );
  NAND2_X1 U579 ( .A1(G76), .A2(n630), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U581 ( .A(n533), .B(KEYINPUT5), .ZN(n540) );
  NOR2_X2 U582 ( .A1(G651), .A2(n640), .ZN(n647) );
  NAND2_X1 U583 ( .A1(G51), .A2(n647), .ZN(n537) );
  NOR2_X1 U584 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n535), .Z(n646) );
  NAND2_X1 U586 ( .A1(G63), .A2(n646), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT6), .B(n538), .Z(n539) );
  NAND2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U590 ( .A(n541), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U591 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U592 ( .A1(G102), .A2(n869), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G138), .A2(n870), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U595 ( .A1(G126), .A2(n874), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G114), .A2(n873), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U598 ( .A1(n547), .A2(n546), .ZN(G164) );
  NAND2_X1 U599 ( .A1(G64), .A2(n646), .ZN(n548) );
  XNOR2_X1 U600 ( .A(n548), .B(KEYINPUT68), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G52), .A2(n647), .ZN(n549) );
  XOR2_X1 U602 ( .A(KEYINPUT69), .B(n549), .Z(n550) );
  NAND2_X1 U603 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U604 ( .A1(G90), .A2(n632), .ZN(n553) );
  NAND2_X1 U605 ( .A1(G77), .A2(n630), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U608 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U609 ( .A(KEYINPUT70), .B(n557), .ZN(G171) );
  INV_X1 U610 ( .A(G171), .ZN(G301) );
  NAND2_X1 U611 ( .A1(G85), .A2(n632), .ZN(n559) );
  NAND2_X1 U612 ( .A1(G72), .A2(n630), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U614 ( .A1(G47), .A2(n647), .ZN(n561) );
  NAND2_X1 U615 ( .A1(G60), .A2(n646), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U617 ( .A1(n563), .A2(n562), .ZN(G290) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G860), .ZN(n596) );
  NAND2_X1 U620 ( .A1(G81), .A2(n632), .ZN(n564) );
  XNOR2_X1 U621 ( .A(n564), .B(KEYINPUT72), .ZN(n565) );
  XNOR2_X1 U622 ( .A(KEYINPUT12), .B(n565), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n630), .A2(G68), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n516), .ZN(n568) );
  XNOR2_X1 U625 ( .A(n568), .B(KEYINPUT13), .ZN(n570) );
  NAND2_X1 U626 ( .A1(G43), .A2(n647), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n646), .A2(G56), .ZN(n571) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n571), .Z(n572) );
  NOR2_X1 U630 ( .A1(n573), .A2(n572), .ZN(n574) );
  OR2_X1 U631 ( .A1(n596), .A2(n990), .ZN(G153) );
  INV_X1 U632 ( .A(G57), .ZN(G237) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  NAND2_X1 U635 ( .A1(G91), .A2(n632), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G78), .A2(n630), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G53), .A2(n647), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G65), .A2(n646), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n700) );
  INV_X1 U642 ( .A(n700), .ZN(G299) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U644 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n821) );
  NAND2_X1 U646 ( .A1(n821), .A2(G567), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT71), .ZN(n583) );
  XNOR2_X1 U648 ( .A(KEYINPUT11), .B(n583), .ZN(G234) );
  NAND2_X1 U649 ( .A1(G301), .A2(G868), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G92), .A2(n632), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G66), .A2(n646), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G79), .A2(n630), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G54), .A2(n647), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT75), .B(n588), .Z(n589) );
  NOR2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U658 ( .A(KEYINPUT15), .B(n591), .ZN(n972) );
  INV_X1 U659 ( .A(G868), .ZN(n658) );
  NAND2_X1 U660 ( .A1(n972), .A2(n658), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(G284) );
  NOR2_X1 U662 ( .A1(G286), .A2(n658), .ZN(n595) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n596), .A2(G559), .ZN(n597) );
  INV_X1 U666 ( .A(n972), .ZN(n620) );
  NAND2_X1 U667 ( .A1(n597), .A2(n620), .ZN(n598) );
  XNOR2_X1 U668 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(n990), .A2(G868), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G868), .A2(n620), .ZN(n599) );
  NOR2_X1 U671 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n601), .A2(n600), .ZN(G282) );
  XOR2_X1 U673 ( .A(G2100), .B(KEYINPUT78), .Z(n611) );
  NAND2_X1 U674 ( .A1(G111), .A2(n873), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G99), .A2(n869), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n874), .A2(G123), .ZN(n604) );
  XNOR2_X1 U678 ( .A(n604), .B(KEYINPUT18), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G135), .A2(n870), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U681 ( .A(KEYINPUT77), .B(n607), .Z(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n929) );
  XNOR2_X1 U683 ( .A(G2096), .B(n929), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U685 ( .A1(G55), .A2(n647), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n612), .B(KEYINPUT80), .ZN(n619) );
  NAND2_X1 U687 ( .A1(G80), .A2(n630), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G67), .A2(n646), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G93), .A2(n632), .ZN(n615) );
  XNOR2_X1 U691 ( .A(KEYINPUT79), .B(n615), .ZN(n616) );
  NOR2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n659) );
  NAND2_X1 U694 ( .A1(G559), .A2(n620), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n621), .B(n990), .ZN(n656) );
  NOR2_X1 U696 ( .A1(n656), .A2(G860), .ZN(n622) );
  XOR2_X1 U697 ( .A(n659), .B(n622), .Z(G145) );
  NAND2_X1 U698 ( .A1(G88), .A2(n632), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G75), .A2(n630), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n646), .A2(G62), .ZN(n625) );
  XOR2_X1 U702 ( .A(KEYINPUT84), .B(n625), .Z(n626) );
  NOR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n647), .A2(G50), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(G303) );
  INV_X1 U706 ( .A(G303), .ZN(G166) );
  NAND2_X1 U707 ( .A1(G73), .A2(n630), .ZN(n631) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n631), .Z(n637) );
  NAND2_X1 U709 ( .A1(G86), .A2(n632), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G61), .A2(n646), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U712 ( .A(KEYINPUT83), .B(n635), .Z(n636) );
  NOR2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n647), .A2(G48), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G87), .A2(n640), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n641), .B(KEYINPUT82), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n642) );
  XOR2_X1 U719 ( .A(KEYINPUT81), .B(n642), .Z(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n647), .A2(G49), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(G288) );
  XNOR2_X1 U724 ( .A(G166), .B(G305), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(n659), .ZN(n651) );
  XOR2_X1 U726 ( .A(n651), .B(KEYINPUT19), .Z(n653) );
  XNOR2_X1 U727 ( .A(n700), .B(KEYINPUT85), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n655), .B(G288), .ZN(n895) );
  XOR2_X1 U731 ( .A(n895), .B(n656), .Z(n657) );
  NOR2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n661) );
  NOR2_X1 U733 ( .A1(G868), .A2(n659), .ZN(n660) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XOR2_X1 U736 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U742 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U743 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U744 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U745 ( .A1(G96), .A2(n669), .ZN(n827) );
  NAND2_X1 U746 ( .A1(n827), .A2(G2106), .ZN(n673) );
  NAND2_X1 U747 ( .A1(G69), .A2(G120), .ZN(n670) );
  NOR2_X1 U748 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U749 ( .A1(G108), .A2(n671), .ZN(n828) );
  NAND2_X1 U750 ( .A1(n828), .A2(G567), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n829) );
  NAND2_X1 U752 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U753 ( .A1(n829), .A2(n674), .ZN(n675) );
  XOR2_X1 U754 ( .A(KEYINPUT87), .B(n675), .Z(n826) );
  NAND2_X1 U755 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U756 ( .A1(G2067), .A2(n972), .ZN(n677) );
  XNOR2_X1 U757 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n684) );
  NAND2_X1 U758 ( .A1(G1996), .A2(n684), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n677), .A2(n676), .ZN(n680) );
  NOR2_X1 U760 ( .A1(G1384), .A2(G164), .ZN(n678) );
  XNOR2_X1 U761 ( .A(n678), .B(KEYINPUT64), .ZN(n755) );
  INV_X1 U762 ( .A(n755), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n756) );
  NOR2_X1 U764 ( .A1(n679), .A2(n756), .ZN(n689) );
  NAND2_X1 U765 ( .A1(n680), .A2(n707), .ZN(n683) );
  NOR2_X1 U766 ( .A1(G1996), .A2(n684), .ZN(n681) );
  NOR2_X1 U767 ( .A1(n990), .A2(n681), .ZN(n682) );
  NAND2_X1 U768 ( .A1(n683), .A2(n682), .ZN(n688) );
  NAND2_X1 U769 ( .A1(G1348), .A2(n972), .ZN(n983) );
  NAND2_X1 U770 ( .A1(n983), .A2(n684), .ZN(n685) );
  NOR2_X1 U771 ( .A1(G1341), .A2(n685), .ZN(n686) );
  NOR2_X1 U772 ( .A1(n707), .A2(n686), .ZN(n687) );
  NOR2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n694) );
  INV_X1 U774 ( .A(n689), .ZN(n727) );
  NAND2_X1 U775 ( .A1(G1348), .A2(n727), .ZN(n691) );
  NAND2_X1 U776 ( .A1(G2067), .A2(n707), .ZN(n690) );
  NAND2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n692), .A2(n972), .ZN(n693) );
  NAND2_X1 U779 ( .A1(n707), .A2(G2072), .ZN(n695) );
  XNOR2_X1 U780 ( .A(n695), .B(KEYINPUT27), .ZN(n697) );
  INV_X1 U781 ( .A(G1956), .ZN(n943) );
  NOR2_X1 U782 ( .A1(n943), .A2(n707), .ZN(n696) );
  NOR2_X1 U783 ( .A1(n697), .A2(n696), .ZN(n701) );
  NAND2_X1 U784 ( .A1(n701), .A2(n700), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n704) );
  NOR2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U787 ( .A(n702), .B(KEYINPUT28), .Z(n703) );
  NAND2_X1 U788 ( .A1(n704), .A2(n703), .ZN(n706) );
  XOR2_X1 U789 ( .A(KEYINPUT29), .B(KEYINPUT97), .Z(n705) );
  XNOR2_X1 U790 ( .A(n706), .B(n705), .ZN(n712) );
  XNOR2_X1 U791 ( .A(KEYINPUT94), .B(G1961), .ZN(n952) );
  NOR2_X1 U792 ( .A1(n707), .A2(n952), .ZN(n710) );
  XNOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .ZN(n708) );
  XNOR2_X1 U794 ( .A(n708), .B(KEYINPUT95), .ZN(n1001) );
  NOR2_X1 U795 ( .A1(n1001), .A2(n727), .ZN(n709) );
  NOR2_X1 U796 ( .A1(n710), .A2(n709), .ZN(n719) );
  NOR2_X1 U797 ( .A1(G301), .A2(n719), .ZN(n711) );
  NOR2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n724) );
  NOR2_X1 U799 ( .A1(G2084), .A2(n727), .ZN(n736) );
  NOR2_X1 U800 ( .A1(n739), .A2(n736), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n713), .A2(G8), .ZN(n714) );
  OR2_X1 U802 ( .A1(n714), .A2(KEYINPUT30), .ZN(n716) );
  NAND2_X1 U803 ( .A1(n714), .A2(KEYINPUT30), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U805 ( .A(n717), .B(KEYINPUT98), .ZN(n718) );
  NOR2_X1 U806 ( .A1(G168), .A2(n718), .ZN(n721) );
  AND2_X1 U807 ( .A1(n719), .A2(G301), .ZN(n720) );
  NOR2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U809 ( .A(n722), .B(KEYINPUT31), .ZN(n723) );
  NOR2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U811 ( .A(n725), .B(KEYINPUT99), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n737), .A2(G286), .ZN(n726) );
  XNOR2_X1 U813 ( .A(n726), .B(KEYINPUT100), .ZN(n733) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n785), .ZN(n729) );
  NOR2_X1 U815 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U816 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U817 ( .A(KEYINPUT101), .B(n730), .Z(n731) );
  NAND2_X1 U818 ( .A1(n731), .A2(G303), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U820 ( .A1(n734), .A2(G8), .ZN(n735) );
  XNOR2_X1 U821 ( .A(n735), .B(KEYINPUT32), .ZN(n743) );
  NAND2_X1 U822 ( .A1(G8), .A2(n736), .ZN(n741) );
  INV_X1 U823 ( .A(n737), .ZN(n738) );
  NOR2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U826 ( .A1(n743), .A2(n742), .ZN(n779) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n749), .A2(n744), .ZN(n976) );
  INV_X1 U830 ( .A(KEYINPUT33), .ZN(n745) );
  AND2_X1 U831 ( .A1(n976), .A2(n745), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n779), .A2(n746), .ZN(n754) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n975) );
  INV_X1 U834 ( .A(n975), .ZN(n747) );
  NOR2_X1 U835 ( .A1(n747), .A2(n785), .ZN(n748) );
  NOR2_X1 U836 ( .A1(KEYINPUT33), .A2(n748), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n785), .A2(n750), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n776) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n969) );
  NOR2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n816) );
  XOR2_X1 U843 ( .A(KEYINPUT90), .B(G1991), .Z(n1002) );
  NAND2_X1 U844 ( .A1(G95), .A2(n869), .ZN(n758) );
  NAND2_X1 U845 ( .A1(G131), .A2(n870), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n762) );
  NAND2_X1 U847 ( .A1(G107), .A2(n873), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G119), .A2(n874), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n881) );
  NOR2_X1 U851 ( .A1(n1002), .A2(n881), .ZN(n763) );
  XNOR2_X1 U852 ( .A(n763), .B(KEYINPUT91), .ZN(n773) );
  XOR2_X1 U853 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n765) );
  NAND2_X1 U854 ( .A1(G105), .A2(n869), .ZN(n764) );
  XNOR2_X1 U855 ( .A(n765), .B(n764), .ZN(n769) );
  NAND2_X1 U856 ( .A1(G117), .A2(n873), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G129), .A2(n874), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n870), .A2(G141), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n885) );
  NAND2_X1 U862 ( .A1(G1996), .A2(n885), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n928) );
  NAND2_X1 U864 ( .A1(n816), .A2(n928), .ZN(n805) );
  XNOR2_X1 U865 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U866 ( .A1(n816), .A2(n982), .ZN(n774) );
  AND2_X1 U867 ( .A1(n805), .A2(n774), .ZN(n787) );
  AND2_X1 U868 ( .A1(n969), .A2(n787), .ZN(n775) );
  NAND2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n791) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U871 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n781) );
  AND2_X1 U873 ( .A1(n785), .A2(n787), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n789) );
  NOR2_X1 U875 ( .A1(G1981), .A2(G305), .ZN(n782) );
  XNOR2_X1 U876 ( .A(n782), .B(KEYINPUT93), .ZN(n783) );
  XNOR2_X1 U877 ( .A(KEYINPUT24), .B(n783), .ZN(n784) );
  NOR2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n803) );
  XNOR2_X1 U882 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  NAND2_X1 U883 ( .A1(G104), .A2(n869), .ZN(n793) );
  NAND2_X1 U884 ( .A1(G140), .A2(n870), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U886 ( .A(KEYINPUT34), .B(n794), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n873), .A2(G116), .ZN(n795) );
  XNOR2_X1 U888 ( .A(n795), .B(KEYINPUT88), .ZN(n797) );
  NAND2_X1 U889 ( .A1(G128), .A2(n874), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U891 ( .A(KEYINPUT35), .B(n798), .ZN(n799) );
  XNOR2_X1 U892 ( .A(KEYINPUT89), .B(n799), .ZN(n800) );
  NOR2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U894 ( .A(KEYINPUT36), .B(n802), .ZN(n890) );
  NOR2_X1 U895 ( .A1(n813), .A2(n890), .ZN(n932) );
  NAND2_X1 U896 ( .A1(n816), .A2(n932), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n803), .A2(n811), .ZN(n804) );
  XNOR2_X1 U898 ( .A(n804), .B(KEYINPUT102), .ZN(n819) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n885), .ZN(n920) );
  INV_X1 U900 ( .A(n805), .ZN(n808) );
  AND2_X1 U901 ( .A1(n1002), .A2(n881), .ZN(n927) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n927), .A2(n806), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n920), .A2(n809), .ZN(n810) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n810), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n813), .A2(n890), .ZN(n936) );
  NAND2_X1 U909 ( .A1(n814), .A2(n936), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U911 ( .A(KEYINPUT103), .B(n817), .Z(n818) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U913 ( .A(n820), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n821), .ZN(G217) );
  NAND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n822) );
  XNOR2_X1 U916 ( .A(KEYINPUT105), .B(n822), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(G661), .ZN(n824) );
  XNOR2_X1 U918 ( .A(KEYINPUT106), .B(n824), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  INV_X1 U927 ( .A(n829), .ZN(G319) );
  XOR2_X1 U928 ( .A(KEYINPUT110), .B(G1976), .Z(n831) );
  XNOR2_X1 U929 ( .A(G1961), .B(G1971), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U931 ( .A(n832), .B(KEYINPUT41), .Z(n834) );
  XNOR2_X1 U932 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U934 ( .A(G1981), .B(G1956), .Z(n836) );
  XNOR2_X1 U935 ( .A(G1986), .B(G1966), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U937 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U938 ( .A(KEYINPUT109), .B(G2474), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U940 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2678), .B(KEYINPUT43), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U943 ( .A(KEYINPUT42), .B(G2090), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2100), .B(G2096), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n850) );
  XOR2_X1 U949 ( .A(G2078), .B(G2084), .Z(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(G227) );
  NAND2_X1 U951 ( .A1(n874), .A2(G124), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U953 ( .A1(G136), .A2(n870), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G112), .A2(n873), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G100), .A2(n869), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(KEYINPUT111), .B(n856), .Z(n857) );
  NOR2_X1 U959 ( .A1(n858), .A2(n857), .ZN(G162) );
  XNOR2_X1 U960 ( .A(G160), .B(G164), .ZN(n867) );
  NAND2_X1 U961 ( .A1(G118), .A2(n873), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G130), .A2(n874), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G106), .A2(n869), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G142), .A2(n870), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U967 ( .A(KEYINPUT45), .B(n863), .Z(n864) );
  NOR2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n929), .B(n868), .ZN(n889) );
  NAND2_X1 U971 ( .A1(G103), .A2(n869), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G139), .A2(n870), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U974 ( .A1(G115), .A2(n873), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G127), .A2(n874), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(KEYINPUT112), .B(n877), .Z(n878) );
  XNOR2_X1 U978 ( .A(KEYINPUT47), .B(n878), .ZN(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n915) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n883) );
  XNOR2_X1 U981 ( .A(n881), .B(KEYINPUT113), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n915), .B(n884), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n885), .B(G162), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U987 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U988 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U989 ( .A(G286), .B(KEYINPUT114), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n972), .B(G301), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n990), .B(n895), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U994 ( .A1(G37), .A2(n898), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2443), .B(G2427), .Z(n900) );
  XNOR2_X1 U996 ( .A(G2438), .B(G2454), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(G2435), .Z(n903) );
  XNOR2_X1 U999 ( .A(G1348), .B(G1341), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1001 ( .A(G2430), .B(G2446), .Z(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT104), .B(G2451), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(n908) );
  NAND2_X1 U1005 ( .A1(G14), .A2(n908), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n914), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n914), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G2072), .B(n915), .Z(n917) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT50), .ZN(n925) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT117), .B(n921), .Z(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n922) );
  XNOR2_X1 U1023 ( .A(n923), .B(n922), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n938) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(KEYINPUT115), .B(n934), .Z(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  XOR2_X1 U1034 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n1015) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n1015), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n941), .A2(G29), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT119), .B(n942), .ZN(n1026) );
  XNOR2_X1 U1038 ( .A(G20), .B(n943), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(G1341), .B(G19), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(G1981), .B(G6), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1043 ( .A(KEYINPUT59), .B(G1348), .Z(n948) );
  XNOR2_X1 U1044 ( .A(G4), .B(n948), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT60), .B(n951), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n952), .B(G5), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G21), .B(G1966), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n966) );
  XNOR2_X1 U1051 ( .A(G1986), .B(G24), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G1971), .B(G22), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT124), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT125), .B(n960), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1058 ( .A(KEYINPUT126), .B(n963), .Z(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n964), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT61), .B(n967), .Z(n968) );
  NOR2_X1 U1062 ( .A1(G16), .A2(n968), .ZN(n1023) );
  XOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .Z(n997) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(n971), .B(KEYINPUT57), .ZN(n994) );
  XNOR2_X1 U1067 ( .A(G1961), .B(G301), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n972), .A2(G1348), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n989) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n979) );
  INV_X1 U1071 ( .A(G1971), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(G166), .A2(n977), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1074 ( .A(KEYINPUT122), .B(n980), .Z(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1077 ( .A(G1956), .B(G299), .Z(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT121), .B(n985), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G1341), .B(n990), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(KEYINPUT123), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1020) );
  XNOR2_X1 U1086 ( .A(G2067), .B(G26), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G33), .B(G2072), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1008) );
  XOR2_X1 U1089 ( .A(G1996), .B(G32), .Z(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(G28), .ZN(n1006) );
  XOR2_X1 U1091 ( .A(n1001), .B(G27), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(n1002), .B(G25), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1009), .B(KEYINPUT53), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(G2084), .B(G34), .Z(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT54), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G35), .B(G2090), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(n1016), .B(n1015), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(G29), .A2(n1017), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT120), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(G11), .A2(n1021), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(n1024), .B(KEYINPUT127), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1027), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

