//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT13), .B1(new_n187), .B2(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(new_n190), .A2(KEYINPUT91), .ZN(new_n191));
  INV_X1    g005(.A(new_n189), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n190), .A2(KEYINPUT91), .B1(KEYINPUT13), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G134), .ZN(new_n195));
  XOR2_X1   g009(.A(G116), .B(G122), .Z(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G107), .ZN(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G122), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G128), .B(G143), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n195), .A2(new_n205), .A3(KEYINPUT92), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n203), .B1(new_n191), .B2(new_n193), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(new_n204), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n200), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n212), .A2(KEYINPUT93), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n202), .B(new_n203), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT14), .A3(G122), .ZN(new_n216));
  OAI211_X1 g030(.A(G107), .B(new_n216), .C1(new_n196), .C2(KEYINPUT14), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(KEYINPUT93), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n214), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT9), .B(G234), .ZN(new_n221));
  INV_X1    g035(.A(G217), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(new_n222), .A3(G953), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT94), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n219), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(new_n206), .B2(new_n210), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT94), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n223), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n220), .A2(new_n224), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G478), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(KEYINPUT15), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n235), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT20), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n241));
  INV_X1    g055(.A(G140), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G125), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n243), .A2(KEYINPUT72), .A3(KEYINPUT16), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G125), .B(G140), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT72), .B1(new_n246), .B2(KEYINPUT16), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n243), .A2(KEYINPUT16), .ZN(new_n248));
  OAI211_X1 g062(.A(G146), .B(new_n245), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(new_n252), .C1(new_n246), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G953), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n256), .A2(new_n258), .A3(G214), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n187), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT68), .B(G953), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n262), .A2(G143), .A3(G214), .A4(new_n259), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n261), .B2(new_n263), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n249), .B(new_n254), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n261), .A2(new_n263), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT18), .A3(G131), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n246), .B(new_n252), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT18), .A2(G131), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n261), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G113), .B(G122), .ZN(new_n275));
  INV_X1    g089(.A(G104), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT17), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n268), .A2(KEYINPUT17), .A3(G131), .ZN(new_n281));
  INV_X1    g095(.A(G125), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G140), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n243), .A2(new_n283), .A3(KEYINPUT16), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n248), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n252), .B1(new_n286), .B2(new_n244), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n281), .A2(new_n287), .A3(new_n249), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n277), .B(new_n273), .C1(new_n280), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n279), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(G475), .A2(G902), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n241), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n268), .A2(G131), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT17), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(new_n287), .A3(new_n249), .A4(new_n281), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n277), .B1(new_n298), .B2(new_n273), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n232), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n240), .A2(new_n292), .B1(new_n300), .B2(G475), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n290), .A2(new_n291), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT89), .ZN(new_n303));
  INV_X1    g117(.A(new_n291), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n279), .B2(new_n289), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n241), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(KEYINPUT20), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n301), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n301), .B2(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n239), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT3), .B1(new_n276), .B2(G107), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n199), .A3(G104), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n276), .A2(G107), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT77), .A3(G101), .ZN(new_n317));
  INV_X1    g131(.A(G101), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n312), .A2(new_n314), .A3(new_n318), .A4(new_n315), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(KEYINPUT4), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT2), .B(G113), .Z(new_n322));
  XNOR2_X1  g136(.A(G116), .B(G119), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G116), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n215), .A2(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n321), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n322), .A2(new_n323), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n329), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(KEYINPUT66), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n316), .A2(KEYINPUT77), .A3(new_n335), .A4(G101), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n320), .A2(new_n331), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G113), .B1(new_n326), .B2(KEYINPUT5), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n332), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n276), .A2(G107), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n199), .A2(G104), .ZN(new_n344));
  OAI21_X1  g158(.A(G101), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n319), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT84), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n330), .B1(new_n340), .B2(new_n339), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n319), .A2(new_n345), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n337), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G110), .B(G122), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n337), .A2(new_n347), .A3(new_n353), .A4(new_n351), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n252), .A2(G143), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n187), .A2(G146), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT0), .A2(G128), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(KEYINPUT0), .A2(G128), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G143), .B(G146), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n361), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(G125), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n358), .A2(new_n359), .A3(new_n369), .A4(G128), .ZN(new_n370));
  INV_X1    g184(.A(G128), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n358), .B2(KEYINPUT1), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n372), .B2(new_n365), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n367), .B(new_n368), .C1(G125), .C2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n364), .A2(KEYINPUT85), .A3(G125), .A4(new_n366), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n255), .A2(G224), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n352), .A2(new_n379), .A3(new_n354), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n357), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(KEYINPUT7), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n374), .A2(KEYINPUT7), .A3(new_n377), .A4(new_n375), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n338), .A2(KEYINPUT86), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n338), .A2(KEYINPUT86), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n385), .A2(new_n340), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n349), .B1(new_n387), .B2(new_n330), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n353), .B(KEYINPUT8), .Z(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n346), .B2(new_n348), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n383), .A2(new_n384), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(G902), .B1(new_n391), .B2(new_n356), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G210), .B1(G237), .B2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n381), .A2(new_n392), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n397), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G214), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n262), .ZN(new_n404));
  NAND2_X1  g218(.A1(G234), .A2(G237), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n404), .A2(G902), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT21), .B(G898), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n405), .A2(G952), .A3(new_n255), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n403), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n399), .A2(new_n401), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n311), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT22), .B(G137), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT74), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT75), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(G119), .B(G128), .Z(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT24), .B(G110), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT23), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n325), .B2(G128), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n371), .A2(KEYINPUT23), .A3(G119), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n425), .B(new_n426), .C1(G119), .C2(new_n371), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G110), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT71), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n430), .A3(G110), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n423), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n287), .A2(new_n249), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n421), .A2(new_n422), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n427), .B2(G110), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n246), .A2(new_n252), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n249), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT73), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT73), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(new_n441), .A3(new_n438), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n420), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n439), .A2(new_n418), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n414), .B1(new_n445), .B2(G902), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n443), .A2(KEYINPUT25), .A3(new_n232), .A4(new_n444), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n222), .B1(G234), .B2(new_n232), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n445), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n331), .A2(new_n334), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G137), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G134), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n203), .A2(G137), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n264), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT64), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT67), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT11), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n203), .B2(G137), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(KEYINPUT11), .A3(G134), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n264), .A4(new_n460), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n462), .A2(new_n463), .A3(new_n373), .A4(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n461), .A2(KEYINPUT64), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT64), .ZN(new_n470));
  AOI211_X1 g284(.A(new_n470), .B(new_n264), .C1(new_n459), .C2(new_n460), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n373), .B(new_n467), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(new_n466), .A3(new_n460), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G131), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n467), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n364), .A2(new_n366), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n468), .A2(new_n473), .A3(KEYINPUT30), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n472), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT65), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n483), .B(KEYINPUT30), .C1(new_n478), .C2(new_n472), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n457), .B(new_n479), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT70), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n262), .A2(G210), .A3(new_n259), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT26), .B(G101), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n489), .B2(new_n490), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n468), .A2(new_n473), .A3(new_n456), .A4(new_n478), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n485), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT31), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n485), .A2(KEYINPUT31), .A3(new_n494), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n457), .B2(new_n480), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n457), .A2(new_n480), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n495), .A2(new_n501), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n494), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n509));
  NOR2_X1   g323(.A1(G472), .A2(G902), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n506), .B1(new_n498), .B2(new_n499), .ZN(new_n512));
  INV_X1    g326(.A(new_n510), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT32), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G472), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n485), .A2(new_n495), .ZN(new_n517));
  INV_X1    g331(.A(new_n494), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT29), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n504), .A2(new_n505), .A3(new_n494), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n502), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n468), .A2(new_n473), .A3(new_n478), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n457), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n495), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n523), .B1(new_n526), .B2(KEYINPUT28), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n518), .A2(new_n520), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n516), .B1(new_n522), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n455), .B1(new_n515), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n370), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT78), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT78), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n358), .A2(new_n538), .A3(KEYINPUT1), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(G128), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n540), .B2(new_n360), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n534), .B1(new_n541), .B2(new_n346), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n320), .A2(new_n477), .A3(new_n336), .ZN(new_n543));
  INV_X1    g357(.A(new_n476), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n349), .A2(KEYINPUT10), .A3(new_n373), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G140), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT76), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n262), .A2(G227), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n548), .B(new_n549), .Z(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT82), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n546), .A2(KEYINPUT82), .A3(new_n550), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n476), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n546), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n369), .B1(G143), .B2(new_n252), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n371), .B1(new_n559), .B2(new_n538), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n365), .B1(new_n560), .B2(new_n537), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n349), .B1(new_n561), .B2(new_n535), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n346), .B(new_n370), .C1(new_n365), .C2(new_n372), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n544), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT81), .B1(new_n564), .B2(KEYINPUT12), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n540), .A2(new_n360), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n346), .B1(new_n566), .B2(new_n370), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n349), .A2(new_n373), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n476), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT81), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT12), .B(new_n476), .C1(new_n567), .C2(new_n568), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT80), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n562), .A2(new_n563), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT80), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT12), .A4(new_n476), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n558), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n557), .B(G469), .C1(new_n580), .C2(new_n550), .ZN(new_n581));
  INV_X1    g395(.A(G469), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n551), .B1(new_n573), .B2(new_n579), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n550), .B1(new_n556), .B2(new_n546), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n582), .B(new_n232), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n582), .A2(new_n232), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n581), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(G221), .B1(new_n221), .B2(G902), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n588), .A2(KEYINPUT83), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT83), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n413), .A2(new_n532), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  INV_X1    g408(.A(new_n449), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n446), .B2(new_n447), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n453), .ZN(new_n597));
  OAI21_X1  g411(.A(G472), .B1(new_n512), .B2(G902), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n598), .A2(KEYINPUT95), .B1(new_n510), .B2(new_n508), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n600), .B(G472), .C1(new_n512), .C2(G902), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n592), .A2(new_n597), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n403), .B1(new_n396), .B2(new_n398), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n408), .A2(new_n410), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n292), .A2(new_n240), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n300), .A2(G475), .ZN(new_n609));
  INV_X1    g423(.A(new_n306), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT20), .B1(new_n305), .B2(new_n241), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT90), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n301), .A2(new_n307), .A3(new_n308), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n231), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n227), .B2(new_n223), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n223), .B(KEYINPUT96), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n220), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(KEYINPUT97), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n220), .B2(new_n620), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n618), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n234), .A2(G902), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n617), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n233), .A2(new_n234), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT98), .B1(new_n615), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n613), .A3(new_n632), .A4(new_n614), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n603), .A2(new_n607), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND2_X1  g451(.A1(new_n236), .A2(new_n238), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n307), .A3(new_n301), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n606), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n603), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G107), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND2_X1  g458(.A1(new_n598), .A2(KEYINPUT95), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n508), .A2(new_n510), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n601), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n420), .A2(KEYINPUT36), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n440), .A3(new_n442), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n440), .A2(new_n442), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(KEYINPUT36), .B2(new_n420), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n452), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n596), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT100), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n588), .A2(new_n589), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT83), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n638), .B1(new_n613), .B2(new_n614), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n399), .A2(new_n401), .A3(new_n411), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n588), .A2(KEYINPUT83), .A3(new_n589), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n653), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n599), .A2(new_n662), .A3(new_n663), .A4(new_n601), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n654), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT101), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(G12));
  AOI21_X1  g482(.A(new_n653), .B1(new_n515), .B2(new_n531), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n669), .A2(new_n592), .A3(new_n604), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n409), .B1(new_n406), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n639), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  NAND2_X1  g489(.A1(new_n399), .A2(new_n401), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT38), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n615), .A2(new_n239), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n402), .A2(new_n678), .A3(new_n653), .A4(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n672), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n592), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n684));
  INV_X1    g498(.A(new_n517), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n518), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n232), .B1(new_n526), .B2(new_n494), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n515), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n680), .A2(new_n683), .A3(new_n684), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT102), .B(G143), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G45));
  AOI21_X1  g506(.A(new_n530), .B1(new_n511), .B2(new_n514), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n693), .A2(new_n590), .A3(new_n591), .A4(new_n653), .ZN(new_n694));
  INV_X1    g508(.A(new_n672), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n631), .A2(new_n613), .A3(new_n614), .A4(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n694), .A2(KEYINPUT103), .A3(new_n604), .A4(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n669), .A2(new_n592), .A3(new_n604), .A4(new_n697), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NOR2_X1   g517(.A1(new_n583), .A2(new_n584), .ZN(new_n704));
  OAI21_X1  g518(.A(G469), .B1(new_n704), .B2(G902), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n589), .A3(new_n585), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n634), .A2(new_n532), .A3(new_n607), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT41), .B(G113), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT104), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n708), .B(new_n710), .ZN(G15));
  NAND3_X1  g525(.A1(new_n532), .A2(new_n640), .A3(new_n707), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  NOR2_X1   g527(.A1(new_n606), .A2(new_n706), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n669), .A2(new_n658), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  NAND2_X1  g530(.A1(new_n598), .A2(KEYINPUT106), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n718), .B(G472), .C1(new_n512), .C2(G902), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n720));
  INV_X1    g534(.A(new_n527), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n498), .A2(new_n499), .B1(new_n721), .B2(new_n518), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n720), .B1(new_n722), .B2(new_n513), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n500), .B1(new_n494), .B2(new_n527), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(KEYINPUT105), .A3(new_n510), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n717), .A2(new_n719), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n596), .A2(new_n728), .A3(new_n453), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n728), .B1(new_n596), .B2(new_n453), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n727), .A2(new_n732), .A3(new_n679), .A4(new_n714), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NOR3_X1   g548(.A1(new_n726), .A2(new_n653), .A3(new_n696), .ZN(new_n735));
  INV_X1    g549(.A(new_n604), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n706), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND2_X1  g553(.A1(new_n655), .A2(KEYINPUT108), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n588), .A2(new_n741), .A3(new_n589), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n403), .B1(new_n399), .B2(new_n401), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n740), .A2(new_n743), .A3(KEYINPUT109), .A4(new_n742), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT107), .B1(new_n450), .B2(new_n454), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n729), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n511), .A2(KEYINPUT110), .A3(new_n514), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n530), .B1(new_n515), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n748), .A2(new_n754), .A3(new_n697), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n515), .A2(new_n531), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n597), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n746), .B2(new_n747), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n755), .A2(KEYINPUT42), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  AND3_X1   g575(.A1(new_n381), .A2(new_n392), .A3(new_n394), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n394), .B1(new_n381), .B2(new_n392), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT87), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n402), .B1(new_n764), .B2(new_n400), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n741), .B1(new_n588), .B2(new_n589), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT109), .B1(new_n767), .B2(new_n742), .ZN(new_n768));
  INV_X1    g582(.A(new_n747), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n532), .B(new_n673), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n758), .A2(KEYINPUT111), .A3(new_n673), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  OAI21_X1  g589(.A(new_n557), .B1(new_n580), .B2(new_n550), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n582), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n587), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n586), .B1(new_n778), .B2(new_n779), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n585), .B1(new_n784), .B2(KEYINPUT46), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n589), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n681), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(KEYINPUT112), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n787), .B2(new_n681), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n615), .A2(KEYINPUT43), .A3(new_n631), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT43), .B1(new_n615), .B2(new_n631), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n647), .B(new_n662), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n743), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n792), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n458), .ZN(G39));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n786), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT47), .B(new_n589), .C1(new_n783), .C2(new_n785), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n756), .A2(new_n597), .A3(new_n765), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n697), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  NOR2_X1   g623(.A1(new_n309), .A2(new_n310), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n750), .A2(new_n810), .A3(new_n629), .ZN(new_n811));
  INV_X1    g625(.A(new_n589), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n705), .A2(new_n585), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n812), .B(new_n403), .C1(new_n813), .C2(KEYINPUT49), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n811), .B(new_n814), .C1(KEYINPUT49), .C2(new_n813), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(new_n689), .A3(new_n678), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n705), .A2(new_n812), .A3(new_n585), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n804), .A2(new_n805), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT43), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n810), .B2(new_n629), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n410), .B1(new_n820), .B2(new_n793), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n750), .A2(new_n726), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n821), .A2(new_n822), .A3(new_n743), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n678), .A2(new_n402), .A3(new_n706), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n821), .A3(new_n822), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT50), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n825), .A2(new_n821), .A3(new_n828), .A4(new_n822), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n743), .A2(new_n707), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n410), .B(new_n830), .C1(new_n820), .C2(new_n793), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n726), .A2(new_n653), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n689), .A2(new_n830), .A3(new_n455), .A4(new_n410), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n810), .A2(new_n631), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n824), .A2(new_n827), .A3(new_n829), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n831), .A2(new_n754), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT48), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n833), .A2(new_n634), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n821), .A2(new_n822), .A3(new_n737), .ZN(new_n845));
  AND4_X1   g659(.A1(G952), .A2(new_n844), .A3(new_n255), .A4(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n842), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n843), .B1(new_n842), .B2(new_n846), .ZN(new_n848));
  OAI22_X1  g662(.A1(new_n839), .A2(new_n840), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND4_X1   g663(.A1(KEYINPUT51), .A2(new_n827), .A3(new_n829), .A4(new_n835), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n818), .A2(KEYINPUT116), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n804), .A2(new_n852), .A3(new_n805), .A4(new_n817), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n853), .A3(new_n823), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n850), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n855), .B1(new_n850), .B2(new_n854), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n670), .A2(new_n673), .B1(new_n735), .B2(new_n737), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n662), .A2(new_n655), .A3(new_n672), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n615), .A2(new_n239), .A3(new_n736), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n689), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n702), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n702), .A2(new_n860), .A3(new_n867), .A4(new_n863), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n708), .A2(new_n733), .A3(new_n712), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n311), .B(new_n659), .C1(new_n615), .C2(new_n631), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n593), .B(new_n715), .C1(new_n602), .C2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n872), .A3(new_n665), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n638), .A2(new_n612), .A3(new_n672), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n874), .A2(KEYINPUT113), .A3(new_n743), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT113), .B1(new_n874), .B2(new_n743), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n735), .A2(new_n748), .B1(new_n877), .B2(new_n694), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n873), .A2(new_n774), .A3(new_n760), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n869), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(KEYINPUT53), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n864), .A2(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n868), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n879), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT54), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n755), .A2(KEYINPUT42), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n758), .A2(new_n759), .ZN(new_n888));
  AND4_X1   g702(.A1(KEYINPUT111), .A2(new_n748), .A3(new_n532), .A4(new_n673), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT111), .B1(new_n758), .B2(new_n673), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n708), .A2(new_n733), .A3(new_n712), .ZN(new_n892));
  INV_X1    g706(.A(new_n872), .ZN(new_n893));
  INV_X1    g707(.A(new_n665), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n878), .A4(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(KEYINPUT53), .A3(new_n868), .A4(new_n866), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n884), .B1(new_n883), .B2(new_n879), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n859), .A2(new_n886), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT119), .ZN(new_n902));
  OR2_X1    g716(.A1(G952), .A2(G953), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(KEYINPUT119), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n816), .B1(new_n904), .B2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n262), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n232), .B1(new_n897), .B2(new_n898), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n909), .B2(G210), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n357), .A2(new_n380), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n378), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n908), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n913), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n915), .A2(KEYINPUT120), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(KEYINPUT120), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G51));
  AOI211_X1 g732(.A(new_n232), .B(new_n780), .C1(new_n897), .C2(new_n898), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n586), .B(KEYINPUT57), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n897), .A2(new_n899), .A3(new_n898), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n704), .B(KEYINPUT121), .Z(new_n924));
  AOI21_X1  g738(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT122), .B1(new_n925), .B2(new_n907), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  INV_X1    g741(.A(new_n924), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n882), .A2(new_n868), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT53), .B1(new_n929), .B2(new_n896), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n869), .A2(new_n879), .A3(new_n884), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT54), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n900), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n928), .B1(new_n933), .B2(new_n920), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n927), .B(new_n908), .C1(new_n934), .C2(new_n919), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n926), .A2(new_n935), .ZN(G54));
  NAND2_X1  g750(.A1(KEYINPUT58), .A2(G475), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT123), .Z(new_n938));
  AND2_X1   g752(.A1(new_n909), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n908), .B1(new_n939), .B2(new_n290), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n290), .B2(new_n939), .ZN(G60));
  AND2_X1   g755(.A1(new_n617), .A2(new_n625), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n886), .A2(new_n900), .ZN(new_n943));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT59), .Z(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n933), .A2(new_n942), .A3(new_n946), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n907), .ZN(G63));
  NAND2_X1  g763(.A1(new_n897), .A2(new_n898), .ZN(new_n950));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n907), .B1(new_n953), .B2(new_n445), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT61), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n649), .A2(new_n651), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n950), .A2(new_n957), .A3(new_n952), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n954), .B(new_n958), .C1(new_n955), .C2(KEYINPUT61), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G66));
  INV_X1    g776(.A(G224), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n407), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n873), .B2(new_n404), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n911), .B1(G898), .B2(new_n262), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G69));
  OAI21_X1  g781(.A(new_n479), .B1(new_n482), .B2(new_n484), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT125), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n251), .B1(new_n246), .B2(new_n253), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n404), .A2(G900), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n808), .B1(new_n792), .B2(new_n800), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n702), .A2(new_n860), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n754), .A2(new_n862), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n792), .B2(new_n975), .ZN(new_n976));
  OR3_X1    g790(.A1(new_n973), .A2(new_n976), .A3(new_n891), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n971), .B(new_n972), .C1(new_n977), .C2(new_n404), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n658), .B1(new_n810), .B2(new_n629), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n532), .A3(new_n743), .ZN(new_n980));
  OAI221_X1 g794(.A(new_n808), .B1(new_n682), .B2(new_n980), .C1(new_n792), .C2(new_n800), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n974), .A2(new_n690), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n985), .A2(new_n262), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n978), .B1(new_n986), .B2(new_n971), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n988), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n978), .B(new_n990), .C1(new_n986), .C2(new_n971), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT126), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n873), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n985), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n686), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n881), .A2(new_n885), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n519), .A2(new_n496), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n994), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n999), .B(new_n908), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n685), .A2(new_n518), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n996), .B1(new_n977), .B2(new_n997), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1003), .A2(new_n1009), .ZN(G57));
endmodule


