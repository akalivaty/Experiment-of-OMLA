

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U547 ( .A(n711), .Z(n511) );
  AND2_X1 U548 ( .A1(n530), .A2(n745), .ZN(n510) );
  NOR2_X2 U549 ( .A1(G164), .A2(G1384), .ZN(n710) );
  AND2_X2 U550 ( .A1(n540), .A2(n539), .ZN(n888) );
  XNOR2_X1 U551 ( .A(n529), .B(KEYINPUT65), .ZN(n540) );
  NOR2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n535) );
  XNOR2_X1 U553 ( .A(n527), .B(n526), .ZN(n695) );
  NOR2_X1 U554 ( .A1(n605), .A2(n850), .ZN(n606) );
  NOR2_X1 U555 ( .A1(n544), .A2(n543), .ZN(G164) );
  NOR2_X2 U556 ( .A1(G651), .A2(n574), .ZN(n792) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(n535), .Z(n711) );
  XNOR2_X1 U558 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U559 ( .A(n673), .B(KEYINPUT31), .ZN(n674) );
  INV_X1 U560 ( .A(KEYINPUT98), .ZN(n521) );
  AND2_X1 U561 ( .A1(n520), .A2(G8), .ZN(n519) );
  NAND2_X1 U562 ( .A1(n522), .A2(n521), .ZN(n520) );
  INV_X1 U563 ( .A(n682), .ZN(n522) );
  AND2_X2 U564 ( .A1(n525), .A2(n710), .ZN(n664) );
  INV_X1 U565 ( .A(n709), .ZN(n525) );
  XNOR2_X1 U566 ( .A(n524), .B(KEYINPUT32), .ZN(n690) );
  INV_X1 U567 ( .A(KEYINPUT23), .ZN(n596) );
  NOR2_X1 U568 ( .A1(n621), .A2(n971), .ZN(n633) );
  NAND2_X1 U569 ( .A1(n664), .A2(G2072), .ZN(n646) );
  NAND2_X1 U570 ( .A1(n518), .A2(n521), .ZN(n517) );
  INV_X1 U571 ( .A(n683), .ZN(n518) );
  INV_X1 U572 ( .A(KEYINPUT101), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n528), .A2(n962), .ZN(n527) );
  INV_X1 U574 ( .A(G2104), .ZN(n529) );
  XNOR2_X1 U575 ( .A(n597), .B(n596), .ZN(n600) );
  AND2_X1 U576 ( .A1(n523), .A2(n519), .ZN(n512) );
  AND2_X1 U577 ( .A1(n682), .A2(KEYINPUT98), .ZN(n513) );
  XOR2_X1 U578 ( .A(KEYINPUT90), .B(n741), .Z(n514) );
  AND2_X1 U579 ( .A1(n978), .A2(n698), .ZN(n515) );
  AND2_X1 U580 ( .A1(n738), .A2(n514), .ZN(n516) );
  NAND2_X1 U581 ( .A1(n512), .A2(n517), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n683), .A2(n513), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n701), .A2(n694), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n531), .A2(n534), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n532), .A2(n515), .ZN(n531) );
  OR2_X1 U586 ( .A1(n696), .A2(KEYINPUT33), .ZN(n532) );
  OR2_X1 U587 ( .A1(n707), .A2(n706), .ZN(n533) );
  AND2_X1 U588 ( .A1(n708), .A2(n533), .ZN(n534) );
  INV_X1 U589 ( .A(KEYINPUT94), .ZN(n631) );
  INV_X1 U590 ( .A(KEYINPUT96), .ZN(n673) );
  INV_X1 U591 ( .A(KEYINPUT92), .ZN(n665) );
  INV_X1 U592 ( .A(KEYINPUT71), .ZN(n609) );
  XNOR2_X1 U593 ( .A(n609), .B(KEYINPUT12), .ZN(n610) );
  XNOR2_X1 U594 ( .A(n611), .B(n610), .ZN(n613) );
  XNOR2_X1 U595 ( .A(n549), .B(KEYINPUT64), .ZN(n796) );
  INV_X1 U596 ( .A(KEYINPUT13), .ZN(n614) );
  XNOR2_X1 U597 ( .A(n615), .B(n614), .ZN(n618) );
  NAND2_X1 U598 ( .A1(n711), .A2(G138), .ZN(n537) );
  INV_X1 U599 ( .A(G2105), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n888), .A2(G102), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(KEYINPUT88), .ZN(n544) );
  NOR2_X2 U603 ( .A1(n540), .A2(n539), .ZN(n891) );
  NAND2_X1 U604 ( .A1(G126), .A2(n891), .ZN(n542) );
  AND2_X1 U605 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NAND2_X1 U606 ( .A1(G114), .A2(n892), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  INV_X1 U608 ( .A(G651), .ZN(n548) );
  NOR2_X1 U609 ( .A1(G543), .A2(n548), .ZN(n545) );
  XOR2_X1 U610 ( .A(KEYINPUT1), .B(n545), .Z(n795) );
  NAND2_X1 U611 ( .A1(G64), .A2(n795), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT0), .B(G543), .Z(n574) );
  NAND2_X1 U613 ( .A1(G52), .A2(n792), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n555) );
  NOR2_X1 U615 ( .A1(n574), .A2(n548), .ZN(n791) );
  NAND2_X1 U616 ( .A1(G77), .A2(n791), .ZN(n551) );
  NOR2_X1 U617 ( .A1(G543), .A2(G651), .ZN(n549) );
  NAND2_X1 U618 ( .A1(G90), .A2(n796), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(KEYINPUT69), .B(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT9), .B(n553), .ZN(n554) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(G171) );
  NAND2_X1 U623 ( .A1(G89), .A2(n796), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U625 ( .A1(G76), .A2(n791), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(KEYINPUT5), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G63), .A2(n795), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G51), .A2(n792), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(n562), .Z(n563) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G75), .A2(n791), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G62), .A2(n795), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G88), .A2(n796), .ZN(n568) );
  XNOR2_X1 U639 ( .A(KEYINPUT81), .B(n568), .ZN(n569) );
  NOR2_X1 U640 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n792), .A2(G50), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(G303) );
  NAND2_X1 U643 ( .A1(G74), .A2(G651), .ZN(n573) );
  XNOR2_X1 U644 ( .A(n573), .B(KEYINPUT80), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n574), .A2(G87), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U647 ( .A1(n795), .A2(n577), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G49), .A2(n792), .ZN(n578) );
  XOR2_X1 U649 ( .A(KEYINPUT79), .B(n578), .Z(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(G288) );
  NAND2_X1 U651 ( .A1(n795), .A2(G61), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G86), .A2(n796), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n791), .A2(G73), .ZN(n583) );
  XOR2_X1 U655 ( .A(KEYINPUT2), .B(n583), .Z(n584) );
  NOR2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n792), .A2(G48), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U659 ( .A1(n791), .A2(G72), .ZN(n588) );
  XOR2_X1 U660 ( .A(KEYINPUT67), .B(n588), .Z(n590) );
  NAND2_X1 U661 ( .A1(G85), .A2(n796), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U663 ( .A(KEYINPUT68), .B(n591), .Z(n595) );
  NAND2_X1 U664 ( .A1(G60), .A2(n795), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G47), .A2(n792), .ZN(n592) );
  AND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(G290) );
  NAND2_X1 U668 ( .A1(G101), .A2(n888), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G113), .A2(n892), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT66), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n767) );
  NAND2_X1 U672 ( .A1(G137), .A2(n511), .ZN(n602) );
  NAND2_X1 U673 ( .A1(G125), .A2(n891), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n766) );
  INV_X1 U675 ( .A(G40), .ZN(n603) );
  OR2_X1 U676 ( .A1(n766), .A2(n603), .ZN(n604) );
  OR2_X1 U677 ( .A1(n767), .A2(n604), .ZN(n709) );
  INV_X1 U678 ( .A(n664), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G8), .A2(n605), .ZN(n706) );
  INV_X1 U680 ( .A(G1996), .ZN(n850) );
  XOR2_X1 U681 ( .A(n606), .B(KEYINPUT26), .Z(n608) );
  NAND2_X1 U682 ( .A1(n605), .A2(G1341), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n621) );
  NAND2_X1 U684 ( .A1(n796), .A2(G81), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G68), .A2(n791), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G56), .A2(n795), .ZN(n616) );
  XOR2_X1 U688 ( .A(KEYINPUT14), .B(n616), .Z(n617) );
  NOR2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n792), .A2(G43), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n971) );
  NAND2_X1 U692 ( .A1(G66), .A2(n795), .ZN(n628) );
  NAND2_X1 U693 ( .A1(G79), .A2(n791), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G92), .A2(n796), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n792), .A2(G54), .ZN(n624) );
  XOR2_X1 U697 ( .A(KEYINPUT74), .B(n624), .Z(n625) );
  NOR2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U700 ( .A(n629), .B(KEYINPUT15), .ZN(n630) );
  XOR2_X2 U701 ( .A(KEYINPUT75), .B(n630), .Z(n964) );
  NOR2_X1 U702 ( .A1(n633), .A2(n964), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n639) );
  NAND2_X1 U704 ( .A1(n633), .A2(n964), .ZN(n637) );
  NOR2_X1 U705 ( .A1(n664), .A2(G1348), .ZN(n635) );
  NOR2_X1 U706 ( .A1(G2067), .A2(n605), .ZN(n634) );
  NOR2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n651) );
  NAND2_X1 U710 ( .A1(G65), .A2(n795), .ZN(n641) );
  NAND2_X1 U711 ( .A1(G53), .A2(n792), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U713 ( .A1(G78), .A2(n791), .ZN(n643) );
  NAND2_X1 U714 ( .A1(G91), .A2(n796), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n773) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(n646), .Z(n647) );
  XNOR2_X1 U718 ( .A(KEYINPUT93), .B(n647), .ZN(n649) );
  INV_X1 U719 ( .A(G1956), .ZN(n849) );
  NOR2_X1 U720 ( .A1(n664), .A2(n849), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n773), .A2(n652), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n773), .A2(n652), .ZN(n653) );
  XOR2_X1 U725 ( .A(n653), .B(KEYINPUT28), .Z(n654) );
  NAND2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n657) );
  XNOR2_X1 U727 ( .A(KEYINPUT95), .B(KEYINPUT29), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(n661) );
  INV_X1 U729 ( .A(G1961), .ZN(n970) );
  NAND2_X1 U730 ( .A1(n605), .A2(n970), .ZN(n659) );
  XNOR2_X1 U731 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NAND2_X1 U732 ( .A1(n664), .A2(n943), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n670) );
  NAND2_X1 U734 ( .A1(n670), .A2(G171), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n677) );
  NOR2_X1 U736 ( .A1(G2084), .A2(n605), .ZN(n684) );
  INV_X1 U737 ( .A(G8), .ZN(n662) );
  OR2_X1 U738 ( .A1(n662), .A2(G1966), .ZN(n663) );
  NOR2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n666), .B(n665), .ZN(n685) );
  NAND2_X1 U741 ( .A1(n685), .A2(G8), .ZN(n667) );
  NOR2_X1 U742 ( .A1(n684), .A2(n667), .ZN(n668) );
  XOR2_X1 U743 ( .A(n668), .B(KEYINPUT30), .Z(n669) );
  NOR2_X1 U744 ( .A1(G168), .A2(n669), .ZN(n672) );
  NOR2_X1 U745 ( .A1(G171), .A2(n670), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n686) );
  NAND2_X1 U748 ( .A1(n686), .A2(G286), .ZN(n683) );
  NOR2_X1 U749 ( .A1(G1971), .A2(n706), .ZN(n678) );
  XOR2_X1 U750 ( .A(KEYINPUT97), .B(n678), .Z(n680) );
  NOR2_X1 U751 ( .A1(G2090), .A2(n605), .ZN(n679) );
  NOR2_X1 U752 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U753 ( .A1(n681), .A2(G303), .ZN(n682) );
  NAND2_X1 U754 ( .A1(G8), .A2(n684), .ZN(n688) );
  AND2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n701) );
  NOR2_X1 U758 ( .A1(G288), .A2(G1976), .ZN(n691) );
  XNOR2_X1 U759 ( .A(n691), .B(KEYINPUT99), .ZN(n974) );
  NOR2_X1 U760 ( .A1(G1971), .A2(G303), .ZN(n692) );
  XOR2_X1 U761 ( .A(n692), .B(KEYINPUT100), .Z(n693) );
  AND2_X1 U762 ( .A1(n974), .A2(n693), .ZN(n694) );
  NAND2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n962) );
  NOR2_X1 U764 ( .A1(n706), .A2(n695), .ZN(n696) );
  XOR2_X1 U765 ( .A(G1981), .B(G305), .Z(n978) );
  NOR2_X1 U766 ( .A1(n706), .A2(n974), .ZN(n697) );
  NAND2_X1 U767 ( .A1(KEYINPUT33), .A2(n697), .ZN(n698) );
  NOR2_X1 U768 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U769 ( .A1(G8), .A2(n699), .ZN(n700) );
  XNOR2_X1 U770 ( .A(n700), .B(KEYINPUT102), .ZN(n702) );
  NAND2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n703), .A2(n706), .ZN(n708) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XNOR2_X1 U774 ( .A(n704), .B(KEYINPUT91), .ZN(n705) );
  XNOR2_X1 U775 ( .A(n705), .B(KEYINPUT24), .ZN(n707) );
  NOR2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n752) );
  NAND2_X1 U777 ( .A1(G140), .A2(n511), .ZN(n713) );
  NAND2_X1 U778 ( .A1(G104), .A2(n888), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U780 ( .A(KEYINPUT34), .B(n714), .ZN(n719) );
  NAND2_X1 U781 ( .A1(G128), .A2(n891), .ZN(n716) );
  NAND2_X1 U782 ( .A1(G116), .A2(n892), .ZN(n715) );
  NAND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U784 ( .A(KEYINPUT35), .B(n717), .Z(n718) );
  NOR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U786 ( .A(KEYINPUT36), .B(n720), .Z(n899) );
  XOR2_X1 U787 ( .A(G2067), .B(KEYINPUT37), .Z(n748) );
  AND2_X1 U788 ( .A1(n899), .A2(n748), .ZN(n917) );
  NAND2_X1 U789 ( .A1(n752), .A2(n917), .ZN(n745) );
  XNOR2_X1 U790 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U791 ( .A1(n982), .A2(n752), .ZN(n738) );
  NAND2_X1 U792 ( .A1(G131), .A2(n511), .ZN(n722) );
  NAND2_X1 U793 ( .A1(G95), .A2(n888), .ZN(n721) );
  NAND2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U795 ( .A1(G119), .A2(n891), .ZN(n723) );
  XNOR2_X1 U796 ( .A(KEYINPUT89), .B(n723), .ZN(n724) );
  NOR2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U798 ( .A1(n892), .A2(G107), .ZN(n726) );
  NAND2_X1 U799 ( .A1(n727), .A2(n726), .ZN(n882) );
  AND2_X1 U800 ( .A1(n882), .A2(G1991), .ZN(n736) );
  NAND2_X1 U801 ( .A1(G141), .A2(n511), .ZN(n729) );
  NAND2_X1 U802 ( .A1(G117), .A2(n892), .ZN(n728) );
  NAND2_X1 U803 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n888), .A2(G105), .ZN(n730) );
  XOR2_X1 U805 ( .A(KEYINPUT38), .B(n730), .Z(n731) );
  NOR2_X1 U806 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U807 ( .A1(n891), .A2(G129), .ZN(n733) );
  NAND2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n883) );
  AND2_X1 U809 ( .A1(n883), .A2(G1996), .ZN(n735) );
  NOR2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n914) );
  INV_X1 U811 ( .A(n752), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n914), .A2(n737), .ZN(n741) );
  NAND2_X1 U813 ( .A1(n510), .A2(n516), .ZN(n755) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n883), .ZN(n932) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n882), .ZN(n919) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n739) );
  NOR2_X1 U817 ( .A1(n919), .A2(n739), .ZN(n740) );
  NOR2_X1 U818 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U819 ( .A1(n932), .A2(n742), .ZN(n744) );
  XOR2_X1 U820 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n743) );
  XNOR2_X1 U821 ( .A(n744), .B(n743), .ZN(n746) );
  NAND2_X1 U822 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U823 ( .A(n747), .B(KEYINPUT104), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n748), .A2(n899), .ZN(n749) );
  XNOR2_X1 U825 ( .A(n749), .B(KEYINPUT105), .ZN(n929) );
  NAND2_X1 U826 ( .A1(n750), .A2(n929), .ZN(n751) );
  XNOR2_X1 U827 ( .A(KEYINPUT106), .B(n751), .ZN(n753) );
  NAND2_X1 U828 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U829 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U830 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U831 ( .A(G2443), .B(G2446), .Z(n758) );
  XNOR2_X1 U832 ( .A(G2427), .B(G2451), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n758), .B(n757), .ZN(n764) );
  XOR2_X1 U834 ( .A(G2430), .B(G2454), .Z(n760) );
  XNOR2_X1 U835 ( .A(G1348), .B(G1341), .ZN(n759) );
  XNOR2_X1 U836 ( .A(n760), .B(n759), .ZN(n762) );
  XOR2_X1 U837 ( .A(G2435), .B(G2438), .Z(n761) );
  XNOR2_X1 U838 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U839 ( .A(n764), .B(n763), .Z(n765) );
  AND2_X1 U840 ( .A1(G14), .A2(n765), .ZN(G401) );
  AND2_X1 U841 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  INV_X1 U843 ( .A(G57), .ZN(G237) );
  NOR2_X1 U844 ( .A1(n767), .A2(n766), .ZN(G160) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n768) );
  XOR2_X1 U846 ( .A(n768), .B(KEYINPUT10), .Z(n1024) );
  NAND2_X1 U847 ( .A1(n1024), .A2(G567), .ZN(n769) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(n769), .Z(G234) );
  INV_X1 U849 ( .A(G860), .ZN(n776) );
  OR2_X1 U850 ( .A1(n971), .A2(n776), .ZN(G153) );
  XOR2_X1 U851 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U852 ( .A1(G868), .A2(G301), .ZN(n770) );
  XOR2_X1 U853 ( .A(KEYINPUT73), .B(n770), .Z(n772) );
  OR2_X1 U854 ( .A1(n964), .A2(G868), .ZN(n771) );
  NAND2_X1 U855 ( .A1(n772), .A2(n771), .ZN(G284) );
  INV_X1 U856 ( .A(n773), .ZN(G299) );
  INV_X1 U857 ( .A(G868), .ZN(n802) );
  NOR2_X1 U858 ( .A1(G286), .A2(n802), .ZN(n775) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(G297) );
  NAND2_X1 U861 ( .A1(n776), .A2(G559), .ZN(n777) );
  NAND2_X1 U862 ( .A1(n777), .A2(n964), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U864 ( .A1(G868), .A2(n971), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n964), .A2(G868), .ZN(n779) );
  NOR2_X1 U866 ( .A1(G559), .A2(n779), .ZN(n780) );
  NOR2_X1 U867 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U868 ( .A1(G135), .A2(n511), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G111), .A2(n892), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n788) );
  NAND2_X1 U871 ( .A1(G123), .A2(n891), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT18), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n888), .A2(G99), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n918) );
  XNOR2_X1 U876 ( .A(n918), .B(G2096), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n789), .B(KEYINPUT76), .ZN(n790) );
  INV_X1 U878 ( .A(G2100), .ZN(n840) );
  NAND2_X1 U879 ( .A1(n790), .A2(n840), .ZN(G156) );
  INV_X1 U880 ( .A(G303), .ZN(G166) );
  NAND2_X1 U881 ( .A1(G80), .A2(n791), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G55), .A2(n792), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n800) );
  NAND2_X1 U884 ( .A1(n795), .A2(G67), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G93), .A2(n796), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n801), .B(KEYINPUT77), .ZN(n1019) );
  NAND2_X1 U889 ( .A1(n802), .A2(n1019), .ZN(n803) );
  XNOR2_X1 U890 ( .A(n803), .B(KEYINPUT82), .ZN(n812) );
  XNOR2_X1 U891 ( .A(G288), .B(KEYINPUT19), .ZN(n805) );
  XOR2_X1 U892 ( .A(G299), .B(G166), .Z(n804) );
  XNOR2_X1 U893 ( .A(n805), .B(n804), .ZN(n808) );
  XNOR2_X1 U894 ( .A(G290), .B(G305), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n806), .B(n1019), .ZN(n807) );
  XNOR2_X1 U896 ( .A(n808), .B(n807), .ZN(n905) );
  NAND2_X1 U897 ( .A1(G559), .A2(n964), .ZN(n809) );
  XNOR2_X1 U898 ( .A(n971), .B(n809), .ZN(n1018) );
  XOR2_X1 U899 ( .A(n905), .B(n1018), .Z(n810) );
  NAND2_X1 U900 ( .A1(G868), .A2(n810), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2084), .A2(G2078), .ZN(n813) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U904 ( .A1(G2090), .A2(n814), .ZN(n815) );
  XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n815), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n816), .A2(G2072), .ZN(n817) );
  XOR2_X1 U907 ( .A(KEYINPUT83), .B(n817), .Z(G158) );
  XNOR2_X1 U908 ( .A(KEYINPUT84), .B(G44), .ZN(n818) );
  XNOR2_X1 U909 ( .A(n818), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U910 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NAND2_X1 U911 ( .A1(G69), .A2(G120), .ZN(n819) );
  NOR2_X1 U912 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U913 ( .A1(G108), .A2(n820), .ZN(n1022) );
  NAND2_X1 U914 ( .A1(n1022), .A2(G567), .ZN(n827) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n821), .Z(n822) );
  NOR2_X1 U917 ( .A1(G218), .A2(n822), .ZN(n823) );
  XOR2_X1 U918 ( .A(KEYINPUT85), .B(n823), .Z(n824) );
  NAND2_X1 U919 ( .A1(G96), .A2(n824), .ZN(n825) );
  XNOR2_X1 U920 ( .A(KEYINPUT86), .B(n825), .ZN(n1023) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n1023), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n834) );
  NAND2_X1 U923 ( .A1(G661), .A2(G483), .ZN(n828) );
  XOR2_X1 U924 ( .A(KEYINPUT87), .B(n828), .Z(n829) );
  NOR2_X1 U925 ( .A1(n834), .A2(n829), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U927 ( .A1(n1024), .A2(G2106), .ZN(n830) );
  XOR2_X1 U928 ( .A(KEYINPUT107), .B(n830), .Z(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U930 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U932 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U933 ( .A(n834), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT42), .B(G2678), .Z(n836) );
  XNOR2_X1 U935 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U937 ( .A(n837), .B(G2096), .Z(n839) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2072), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n844) );
  XNOR2_X1 U940 ( .A(KEYINPUT108), .B(n840), .ZN(n842) );
  XNOR2_X1 U941 ( .A(G2090), .B(KEYINPUT109), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2084), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U946 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1991), .B(G1986), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n854) );
  XNOR2_X1 U949 ( .A(G1981), .B(n849), .ZN(n852) );
  XOR2_X1 U950 ( .A(n850), .B(G1966), .Z(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n854), .B(n853), .Z(n856) );
  XOR2_X1 U953 ( .A(n970), .B(G1976), .Z(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U955 ( .A(G1971), .B(G2474), .Z(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G100), .A2(n888), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G112), .A2(n892), .ZN(n859) );
  NAND2_X1 U959 ( .A1(n860), .A2(n859), .ZN(n867) );
  NAND2_X1 U960 ( .A1(G124), .A2(n891), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n861), .B(KEYINPUT112), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G136), .A2(n511), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(KEYINPUT113), .B(n865), .Z(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G130), .A2(n891), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G118), .A2(n892), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G142), .A2(n511), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G106), .A2(n888), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n872), .Z(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n918), .B(n875), .ZN(n887) );
  XOR2_X1 U976 ( .A(KEYINPUT117), .B(KEYINPUT48), .Z(n877) );
  XNOR2_X1 U977 ( .A(G160), .B(KEYINPUT46), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U979 ( .A(n878), .B(KEYINPUT114), .Z(n880) );
  XNOR2_X1 U980 ( .A(G164), .B(KEYINPUT116), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U982 ( .A(n881), .B(G162), .Z(n885) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n901) );
  NAND2_X1 U986 ( .A1(G139), .A2(n511), .ZN(n890) );
  NAND2_X1 U987 ( .A1(G103), .A2(n888), .ZN(n889) );
  NAND2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U989 ( .A1(G127), .A2(n891), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G115), .A2(n892), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(KEYINPUT115), .B(n898), .Z(n923) );
  XOR2_X1 U995 ( .A(n923), .B(n899), .Z(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U997 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U998 ( .A(KEYINPUT118), .B(G286), .Z(n904) );
  XNOR2_X1 U999 ( .A(G171), .B(n964), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n907) );
  XOR2_X1 U1001 ( .A(n971), .B(n905), .Z(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n908), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n910), .ZN(n911) );
  AND2_X1 U1007 ( .A1(G319), .A2(n911), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(G225) );
  XNOR2_X1 U1010 ( .A(KEYINPUT119), .B(G225), .ZN(G308) );
  XNOR2_X1 U1012 ( .A(G160), .B(G2084), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(KEYINPUT120), .B(n922), .ZN(n928) );
  XOR2_X1 U1018 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1021 ( .A(KEYINPUT50), .B(n926), .Z(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n936) );
  XNOR2_X1 U1024 ( .A(G2090), .B(G162), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(n931), .B(KEYINPUT121), .ZN(n933) );
  NOR2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(KEYINPUT51), .B(n934), .ZN(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n937), .ZN(n938) );
  INV_X1 U1030 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1031 ( .A1(n938), .A2(n957), .ZN(n939) );
  NAND2_X1 U1032 ( .A1(n939), .A2(G29), .ZN(n1016) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(G33), .B(G2072), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n949) );
  XOR2_X1 U1036 ( .A(G25), .B(G1991), .Z(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(G28), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(n943), .B(G27), .ZN(n945) );
  XOR2_X1 U1039 ( .A(G1996), .B(G32), .Z(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n950), .B(KEYINPUT53), .ZN(n953) );
  XOR2_X1 U1044 ( .A(G2084), .B(KEYINPUT54), .Z(n951) );
  XNOR2_X1 U1045 ( .A(G34), .B(n951), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G35), .B(G2090), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(n957), .B(n956), .ZN(n958) );
  NOR2_X1 U1050 ( .A1(G29), .A2(n958), .ZN(n959) );
  XOR2_X1 U1051 ( .A(KEYINPUT122), .B(n959), .Z(n960) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n960), .ZN(n1014) );
  INV_X1 U1053 ( .A(G16), .ZN(n1010) );
  XOR2_X1 U1054 ( .A(n1010), .B(KEYINPUT56), .Z(n986) );
  XOR2_X1 U1055 ( .A(G303), .B(G1971), .Z(n969) );
  XOR2_X1 U1056 ( .A(G299), .B(G1956), .Z(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(KEYINPUT124), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(n964), .B(G1348), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT123), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(G171), .B(n970), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n971), .B(G1341), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n984) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1070 ( .A(KEYINPUT57), .B(n980), .Z(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n1012) );
  XOR2_X1 U1074 ( .A(G1348), .B(KEYINPUT59), .Z(n987) );
  XNOR2_X1 U1075 ( .A(G4), .B(n987), .ZN(n994) );
  XOR2_X1 U1076 ( .A(G1341), .B(G19), .Z(n989) );
  XOR2_X1 U1077 ( .A(G1956), .B(G20), .Z(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(G6), .B(G1981), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(KEYINPUT125), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1083 ( .A(KEYINPUT60), .B(n995), .Z(n997) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G21), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT126), .B(n998), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(G1961), .B(G5), .Z(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1007) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(G1986), .B(G24), .Z(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1017), .Z(G311) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(G860), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(n1019), .B(KEYINPUT78), .Z(n1020) );
  XNOR2_X1 U1105 ( .A(n1021), .B(n1020), .ZN(G145) );
  INV_X1 U1106 ( .A(G120), .ZN(G236) );
  INV_X1 U1107 ( .A(G96), .ZN(G221) );
  INV_X1 U1108 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(G325) );
  INV_X1 U1110 ( .A(G325), .ZN(G261) );
  INV_X1 U1111 ( .A(G108), .ZN(G238) );
  INV_X1 U1112 ( .A(n1024), .ZN(G223) );
endmodule

