//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n596, new_n599, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n452), .B2(G2106), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G113), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n467), .B2(new_n464), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(G113), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n468), .B(new_n470), .C1(new_n462), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g052(.A1(G124), .A2(new_n477), .B1(new_n463), .B2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n478), .A2(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n476), .C1(new_n460), .C2(new_n461), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(new_n476), .A3(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT71), .B1(new_n462), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n485), .A2(new_n476), .A3(G138), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n484), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n477), .B2(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n503), .B1(new_n500), .B2(G543), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(G166));
  NAND2_X1  g091(.A1(new_n501), .A2(new_n503), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n500), .A2(G543), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n517), .A2(G89), .A3(new_n512), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(KEYINPUT73), .A3(new_n521), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n504), .A2(new_n526), .B1(new_n510), .B2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n504), .A2(G64), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n506), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n504), .A2(G90), .A3(new_n512), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n510), .A2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n530), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g113(.A1(new_n533), .A2(new_n536), .A3(new_n530), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n506), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n510), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n513), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND3_X1  g128(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n510), .A2(new_n556), .A3(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n504), .A2(G91), .A3(new_n512), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n558), .B(new_n559), .C1(new_n506), .C2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G166), .ZN(G303));
  INV_X1    g137(.A(new_n513), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G87), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n510), .A2(G49), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  AOI22_X1  g142(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n506), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n510), .A2(G48), .ZN(new_n570));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n513), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n569), .A2(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n563), .A2(G85), .B1(G47), .B2(new_n510), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n506), .B2(new_n575), .ZN(G290));
  INV_X1    g151(.A(G868), .ZN(new_n577));
  NOR2_X1   g152(.A1(G301), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g153(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G92), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n513), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n504), .A2(G92), .A3(new_n512), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n510), .A2(G54), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n506), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n578), .B1(new_n591), .B2(new_n577), .ZN(G321));
  XNOR2_X1  g167(.A(G321), .B(KEYINPUT78), .ZN(G284));
  OR3_X1    g168(.A1(G168), .A2(KEYINPUT79), .A3(new_n577), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT79), .B1(G168), .B2(new_n577), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n594), .B(new_n595), .C1(G868), .C2(new_n596), .ZN(G297));
  OAI211_X1 g172(.A(new_n594), .B(new_n595), .C1(G868), .C2(new_n596), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G860), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g176(.A1(new_n591), .A2(new_n599), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n488), .A2(new_n465), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n463), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n477), .A2(G123), .ZN(new_n611));
  OR2_X1    g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n612), .B(G2104), .C1(G111), .C2(new_n476), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT81), .B(G2096), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G2438), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G2427), .ZN(new_n621));
  INV_X1    g196(.A(G2427), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G2438), .ZN(new_n623));
  INV_X1    g198(.A(G2430), .ZN(new_n624));
  AND3_X1   g199(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n621), .B2(new_n623), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n621), .A2(new_n623), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G2430), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(new_n618), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n627), .A2(new_n631), .A3(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g211(.A1(new_n634), .A2(new_n627), .A3(new_n631), .A4(KEYINPUT14), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n639), .A3(new_n637), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n641), .A2(KEYINPUT82), .A3(new_n643), .A4(new_n644), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n641), .A2(new_n644), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(new_n642), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(KEYINPUT83), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT84), .Z(new_n670));
  OR2_X1    g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n684), .B(new_n683), .S(new_n676), .Z(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OR3_X1    g262(.A1(new_n682), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n682), .B2(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n691), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n693), .A3(new_n689), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n692), .A2(new_n696), .A3(new_n694), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G21), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G168), .B2(new_n702), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G1966), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT25), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G139), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n488), .A2(new_n476), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT91), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(new_n476), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n717), .B2(G33), .ZN(new_n719));
  INV_X1    g294(.A(G2072), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n702), .A2(G19), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n547), .B2(new_n702), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n719), .A2(new_n720), .B1(G1341), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n717), .A2(G35), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G162), .B2(new_n717), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT29), .Z(new_n726));
  INV_X1    g301(.A(G2090), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n702), .A2(G5), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G171), .B2(new_n702), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT94), .B(G1961), .Z(new_n730));
  OAI221_X1 g305(.A(new_n723), .B1(new_n726), .B2(new_n727), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n705), .B(new_n731), .C1(new_n729), .C2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n717), .A2(G32), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT26), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n488), .A2(G2105), .ZN(new_n737));
  INV_X1    g312(.A(G129), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n465), .A2(G105), .ZN(new_n740));
  INV_X1    g315(.A(G141), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n710), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n733), .B1(new_n743), .B2(new_n717), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT27), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1996), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT31), .B(G11), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT93), .B(G28), .Z(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(KEYINPUT30), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n748), .B2(KEYINPUT30), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n614), .B2(new_n717), .ZN(new_n752));
  AND2_X1   g327(.A1(KEYINPUT24), .A2(G34), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n717), .B1(KEYINPUT24), .B2(G34), .ZN(new_n754));
  OAI22_X1  g329(.A1(G160), .A2(new_n717), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n752), .B1(G2084), .B2(new_n755), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n756), .B1(G1341), .B2(new_n722), .C1(G2084), .C2(new_n755), .ZN(new_n757));
  NAND2_X1  g332(.A1(G164), .A2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G27), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n717), .A2(G26), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT28), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n488), .A2(G140), .A3(new_n476), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n488), .A2(G128), .A3(G2105), .ZN(new_n765));
  OR2_X1    g340(.A1(G104), .A2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n766), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n763), .B1(new_n769), .B2(new_n717), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2067), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n759), .A2(new_n760), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n757), .A2(new_n761), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n732), .A2(new_n746), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n719), .A2(new_n720), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT92), .Z(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G1966), .B2(new_n704), .ZN(new_n778));
  NOR2_X1   g353(.A1(G4), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n591), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT90), .B(G1348), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n726), .A2(new_n727), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT95), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n702), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n778), .A2(new_n782), .A3(new_n784), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n463), .A2(G131), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n477), .A2(G119), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n476), .A2(G107), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT85), .Z(new_n795));
  MUX2_X1   g370(.A(G25), .B(new_n795), .S(G29), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT35), .B(G1991), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G24), .B(G290), .S(G16), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1986), .ZN(new_n801));
  AND2_X1   g376(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n702), .A2(G23), .ZN(new_n804));
  INV_X1    g379(.A(G288), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n702), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT87), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n702), .A2(G22), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G166), .B2(new_n702), .ZN(new_n811));
  INV_X1    g386(.A(G1971), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G6), .A2(G16), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n569), .A2(new_n572), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G16), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT32), .B(G1981), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n809), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n803), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT89), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n775), .A2(new_n789), .A3(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  NAND3_X1  g404(.A1(new_n504), .A2(G93), .A3(new_n512), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n510), .A2(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n504), .A2(G67), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G651), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n833), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n506), .B1(new_n834), .B2(new_n835), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT96), .B1(new_n840), .B2(new_n832), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n547), .A3(new_n841), .ZN(new_n842));
  OAI221_X1 g417(.A(KEYINPUT96), .B1(new_n840), .B2(new_n832), .C1(new_n543), .C2(new_n546), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT38), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n591), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n848), .A2(new_n849), .A3(G860), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n833), .A2(new_n837), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  NAND2_X1  g429(.A1(new_n477), .A2(G130), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n476), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G142), .B2(new_n463), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n607), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n794), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n492), .A2(new_n496), .A3(new_n768), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n768), .B1(new_n492), .B2(new_n496), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n739), .A2(new_n742), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n497), .A2(new_n769), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n743), .B1(new_n868), .B2(new_n863), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n862), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n864), .B2(new_n865), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n743), .A3(new_n863), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT97), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n716), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT98), .B1(new_n867), .B2(new_n869), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT99), .B1(new_n878), .B2(new_n715), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n880));
  AOI211_X1 g455(.A(new_n880), .B(new_n716), .C1(new_n875), .C2(new_n877), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n861), .B(new_n874), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n474), .B(new_n614), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(G162), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n874), .B1(new_n879), .B2(new_n881), .ZN(new_n887));
  INV_X1    g462(.A(new_n861), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n882), .A2(KEYINPUT100), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n876), .B1(new_n871), .B2(new_n872), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n715), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n880), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n878), .A2(KEYINPUT99), .A3(new_n715), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n861), .B1(new_n900), .B2(new_n874), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n887), .A2(new_n903), .A3(new_n888), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n884), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n902), .A2(new_n905), .A3(KEYINPUT101), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n885), .B1(new_n894), .B2(new_n901), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n889), .A2(KEYINPUT100), .A3(new_n882), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n893), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g487(.A(G290), .B(new_n815), .ZN(new_n913));
  XNOR2_X1  g488(.A(G166), .B(G288), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n582), .A2(new_n583), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n559), .B1(new_n560), .B2(new_n506), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n504), .A2(G66), .ZN(new_n922));
  NAND2_X1  g497(.A1(G79), .A2(G543), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n924), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n919), .A2(new_n921), .A3(new_n925), .A4(new_n558), .ZN(new_n926));
  OAI21_X1  g501(.A(G299), .B1(new_n587), .B2(new_n584), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT41), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT102), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n602), .B(new_n844), .ZN(new_n938));
  MUX2_X1   g513(.A(new_n932), .B(new_n937), .S(new_n938), .Z(new_n939));
  NOR2_X1   g514(.A1(new_n916), .A2(new_n917), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n918), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n940), .B2(new_n939), .ZN(new_n942));
  MUX2_X1   g517(.A(new_n851), .B(new_n942), .S(G868), .Z(G295));
  MUX2_X1   g518(.A(new_n851), .B(new_n942), .S(G868), .Z(G331));
  XOR2_X1   g519(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  INV_X1    g521(.A(new_n533), .ZN(new_n947));
  INV_X1    g522(.A(new_n536), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT74), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(G286), .A3(new_n537), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G286), .B1(new_n949), .B2(new_n537), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n844), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(G168), .B1(new_n538), .B2(new_n539), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n954), .A2(new_n843), .A3(new_n842), .A4(new_n950), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n953), .A2(new_n955), .B1(new_n929), .B2(new_n931), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(KEYINPUT105), .A3(new_n955), .ZN(new_n957));
  INV_X1    g532(.A(new_n844), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n954), .A4(new_n950), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n956), .B1(new_n961), .B2(new_n933), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n915), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n913), .B(new_n914), .Z(new_n964));
  AOI21_X1  g539(.A(new_n928), .B1(new_n957), .B2(new_n960), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(new_n956), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n946), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n965), .A2(new_n964), .A3(new_n956), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n931), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT106), .A4(new_n930), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n929), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n957), .A2(new_n972), .A3(new_n960), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n934), .A2(new_n953), .A3(new_n936), .A4(new_n955), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n915), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR4_X1   g550(.A1(new_n968), .A2(new_n975), .A3(KEYINPUT43), .A4(G37), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n945), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n975), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n946), .B1(new_n963), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT107), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n963), .A2(new_n966), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n981), .B2(KEYINPUT43), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n977), .B1(new_n980), .B2(new_n982), .ZN(G397));
  AOI21_X1  g558(.A(G1384), .B1(new_n492), .B2(new_n496), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n474), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(G1996), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n743), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT108), .ZN(new_n991));
  INV_X1    g566(.A(new_n988), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n768), .B(G2067), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT109), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n866), .A2(G1996), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n991), .B(new_n995), .C1(new_n988), .C2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n794), .B(new_n798), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(G290), .B(G1986), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n992), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n1004));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(G166), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT113), .B(G8), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(new_n987), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n497), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n985), .A2(KEYINPUT110), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1012), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n987), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT111), .B(G2090), .Z(new_n1025));
  AOI22_X1  g600(.A1(new_n812), .A2(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1010), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1020), .A2(new_n812), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1029), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1008), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1007), .A2(KEYINPUT112), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1007), .A2(KEYINPUT112), .ZN(new_n1034));
  NOR4_X1   g609(.A1(new_n1026), .A2(new_n1033), .A3(new_n1034), .A4(new_n1005), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n805), .A2(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1009), .B1(new_n987), .B2(new_n984), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1038), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1038), .ZN(new_n1045));
  INV_X1    g620(.A(G1981), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT114), .B1(new_n815), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NOR4_X1   g623(.A1(new_n569), .A2(new_n572), .A3(new_n1048), .A4(G1981), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1047), .A2(new_n1049), .B1(new_n1046), .B2(new_n815), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1045), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n815), .A2(new_n1046), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1048), .B1(G305), .B2(G1981), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1049), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT49), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1044), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1032), .A2(new_n1036), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT124), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1032), .A2(new_n1036), .A3(new_n1061), .A4(new_n1058), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n1064));
  INV_X1    g639(.A(G1348), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n987), .A2(new_n984), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1067), .A2(G2067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n591), .B1(new_n1069), .B2(KEYINPUT60), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1066), .A2(new_n1068), .B1(new_n589), .B2(new_n590), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1064), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n591), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1064), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1073), .B(new_n1074), .C1(new_n591), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1996), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1012), .A2(new_n1018), .A3(new_n1079), .A4(new_n1019), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT58), .B(G1341), .Z(new_n1082));
  AOI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(new_n1067), .B2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1012), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(KEYINPUT118), .A3(new_n1079), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n547), .ZN(new_n1087));
  NAND2_X1  g662(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1012), .A2(new_n1018), .A3(new_n1019), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1956), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n921), .B2(KEYINPUT117), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G299), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n921), .B(new_n558), .C1(KEYINPUT117), .C2(KEYINPUT57), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT61), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1097), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n1098), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1086), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n547), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1078), .A2(new_n1089), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1100), .B1(new_n1098), .B2(new_n1071), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1113));
  INV_X1    g688(.A(G1966), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1023), .ZN(new_n1116));
  INV_X1    g691(.A(G2084), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n987), .A4(new_n1021), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1009), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1112), .B1(new_n1119), .B2(G286), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT121), .B1(new_n1121), .B2(G8), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1022), .A2(G2084), .A3(new_n1023), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1966), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT121), .B(G8), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(G286), .A2(new_n1010), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1120), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1024), .A2(G1961), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1020), .B2(G2078), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G301), .B(KEYINPUT54), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n466), .B(KEYINPUT122), .Z(new_n1134));
  OR2_X1    g709(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1135));
  NAND2_X1  g710(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1130), .B(new_n986), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  AND4_X1   g712(.A1(new_n473), .A2(new_n1134), .A3(new_n1016), .A4(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1133), .B1(new_n1011), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1012), .A2(KEYINPUT53), .A3(new_n760), .A4(new_n1016), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1129), .A2(new_n1131), .A3(new_n1140), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1132), .A2(new_n1139), .B1(new_n1141), .B2(new_n1133), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1126), .A2(new_n1112), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1119), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1128), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1111), .A2(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1141), .A2(G171), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1128), .A2(new_n1144), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1128), .B2(new_n1144), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1063), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G288), .A2(G1976), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1038), .B1(new_n1056), .B2(KEYINPUT49), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1045), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1008), .B1(new_n1026), .B2(new_n1005), .ZN(new_n1159));
  AOI211_X1 g734(.A(G286), .B(new_n1009), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1058), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(KEYINPUT63), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1035), .B1(new_n1032), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1058), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT116), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT116), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1162), .B(new_n1169), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1002), .B1(new_n1152), .B2(new_n1171), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n988), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT46), .B1(new_n988), .B2(G1996), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n993), .A2(new_n866), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1173), .A2(new_n1174), .B1(new_n992), .B2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT47), .ZN(new_n1177));
  OR3_X1    g752(.A1(new_n997), .A2(new_n795), .A3(new_n798), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n768), .A2(G2067), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n988), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n988), .A2(G1986), .A3(G290), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT48), .Z(new_n1182));
  AOI211_X1 g757(.A(new_n1177), .B(new_n1180), .C1(new_n999), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1172), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n671), .A2(G319), .A3(new_n672), .ZN(new_n1187));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g763(.A1(new_n671), .A2(KEYINPUT125), .A3(G319), .A4(new_n672), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n657), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g768(.A(new_n656), .ZN(new_n1195));
  AOI21_X1  g769(.A(KEYINPUT83), .B1(new_n649), .B2(new_n652), .ZN(new_n1196));
  OAI211_X1 g770(.A(KEYINPUT126), .B(new_n1191), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n1194), .A2(new_n700), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g772(.A(new_n967), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n963), .A2(new_n946), .A3(new_n978), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n1186), .B1(new_n911), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g776(.A(KEYINPUT101), .B1(new_n902), .B2(new_n905), .ZN(new_n1203));
  NAND4_X1  g777(.A1(new_n909), .A2(new_n907), .A3(new_n884), .A4(new_n904), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n892), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1197), .A2(new_n700), .ZN(new_n1206));
  AOI21_X1  g780(.A(KEYINPUT126), .B1(new_n657), .B2(new_n1191), .ZN(new_n1207));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1208), .B1(new_n967), .B2(new_n976), .ZN(new_n1209));
  NOR3_X1   g783(.A1(new_n1205), .A2(new_n1209), .A3(KEYINPUT127), .ZN(new_n1210));
  NOR2_X1   g784(.A1(new_n1202), .A2(new_n1210), .ZN(G308));
  NAND2_X1  g785(.A1(new_n911), .A2(new_n1201), .ZN(G225));
endmodule


