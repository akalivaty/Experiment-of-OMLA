//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT67), .B(G77), .Z(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n210), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g0023(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n213), .B1(KEYINPUT1), .B2(new_n223), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT68), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G68), .Z(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  XNOR2_X1  g0044(.A(KEYINPUT8), .B(G58), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n208), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n246), .A2(new_n248), .B1(G150), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(new_n208), .B2(new_n201), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n254), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n207), .B2(G20), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n258), .A2(new_n260), .B1(new_n259), .B2(new_n257), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n255), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT9), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT74), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI211_X1 g0071(.A(G1), .B(G13), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(G274), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G226), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n214), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G1698), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n280), .A2(new_n282), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G222), .ZN(new_n290));
  INV_X1    g0090(.A(G223), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G1698), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n284), .B1(new_n289), .B2(new_n290), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n253), .B1(G33), .B2(G41), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n279), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT9), .B(new_n255), .C1(new_n263), .C2(new_n264), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(G190), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT10), .B1(new_n269), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n267), .B(KEYINPUT74), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(new_n301), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n265), .B1(new_n296), .B2(G169), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n296), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G58), .ZN(new_n314));
  INV_X1    g0114(.A(G68), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G58), .A2(G68), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G159), .ZN(new_n319));
  INV_X1    g0119(.A(new_n249), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n292), .B2(G20), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n283), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n325), .B2(G68), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n254), .B1(new_n326), .B2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT76), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT76), .B1(new_n280), .B2(new_n282), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT7), .B1(new_n331), .B2(new_n208), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n292), .A2(new_n322), .A3(G20), .ZN(new_n333));
  OAI21_X1  g0133(.A(G68), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n321), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT77), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT76), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n281), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT76), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n208), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n333), .B1(new_n343), .B2(new_n322), .ZN(new_n344));
  OAI211_X1 g0144(.A(KEYINPUT77), .B(new_n336), .C1(new_n344), .C2(new_n315), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n328), .B1(new_n337), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT78), .ZN(new_n348));
  INV_X1    g0148(.A(new_n258), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n207), .A2(G20), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n246), .A2(new_n350), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n349), .A2(new_n351), .B1(new_n256), .B2(new_n246), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n347), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n336), .B1(new_n344), .B2(new_n315), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT77), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n327), .B1(new_n357), .B2(new_n345), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT78), .B1(new_n358), .B2(new_n352), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT79), .ZN(new_n360));
  INV_X1    g0160(.A(G232), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n275), .B1(new_n277), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n292), .A2(G226), .A3(G1698), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n363), .B(new_n364), .C1(new_n291), .C2(new_n289), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n365), .B2(new_n295), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n360), .B1(new_n366), .B2(new_n309), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(G169), .B2(new_n366), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n360), .A3(new_n309), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n354), .A2(new_n359), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT18), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n354), .A2(new_n359), .A3(new_n373), .A4(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n357), .A2(new_n345), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n352), .B1(new_n375), .B2(new_n328), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n366), .A2(G190), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n297), .B2(new_n366), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT17), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT17), .ZN(new_n381));
  NOR4_X1   g0181(.A1(new_n358), .A2(new_n381), .A3(new_n378), .A4(new_n352), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n372), .A2(new_n374), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G97), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n280), .A2(new_n282), .A3(G232), .A4(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n386), .C1(new_n289), .C2(new_n278), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n295), .ZN(new_n388));
  INV_X1    g0188(.A(G238), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n275), .B1(new_n277), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n295), .B2(new_n387), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(KEYINPUT75), .A3(KEYINPUT13), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(G169), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT14), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT14), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n398), .A2(new_n402), .A3(G169), .A4(new_n399), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n393), .A2(G179), .A3(new_n397), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n257), .A2(new_n315), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT12), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n249), .A2(G50), .B1(G20), .B2(new_n315), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n202), .B2(new_n247), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n258), .A2(G68), .A3(new_n350), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT11), .B1(new_n409), .B2(new_n254), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n392), .B2(KEYINPUT13), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n417), .B2(new_n397), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n398), .A2(G200), .A3(new_n399), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g0221(.A(KEYINPUT71), .B(G107), .Z(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n283), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n423), .B1(new_n289), .B2(new_n361), .C1(new_n389), .C2(new_n293), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n295), .ZN(new_n425));
  INV_X1    g0225(.A(new_n275), .ZN(new_n426));
  INV_X1    g0226(.A(new_n277), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(G244), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G179), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n425), .A2(new_n428), .ZN(new_n431));
  INV_X1    g0231(.A(new_n254), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT15), .B(G87), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  INV_X1    g0234(.A(G87), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n248), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n246), .A2(new_n249), .B1(new_n214), .B2(G20), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n432), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n258), .A2(G77), .A3(new_n350), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n214), .B2(new_n256), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n431), .A2(G169), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n430), .B1(new_n446), .B2(KEYINPUT73), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n443), .A2(new_n445), .ZN(new_n448));
  AOI21_X1  g0248(.A(G169), .B1(new_n425), .B2(new_n428), .ZN(new_n449));
  OR3_X1    g0249(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT73), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n431), .A2(G190), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n443), .A2(new_n445), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(G200), .B2(new_n429), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n447), .A2(new_n450), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n313), .A2(new_n384), .A3(new_n421), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT85), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n280), .A2(new_n282), .A3(G264), .A4(G1698), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT82), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n292), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n280), .A2(new_n282), .A3(G257), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT69), .B(G1698), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n463), .A2(new_n464), .B1(G303), .B2(new_n283), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n272), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n273), .A2(G1), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n295), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G270), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n468), .A2(new_n272), .A3(G274), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(G200), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n207), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n256), .A2(new_n474), .A3(new_n253), .A4(new_n252), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G116), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n257), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  INV_X1    g0281(.A(G97), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n481), .B(new_n208), .C1(G33), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(G20), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n254), .A2(KEYINPUT83), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT83), .B1(new_n254), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(KEYINPUT20), .B(new_n483), .C1(new_n485), .C2(new_n486), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n480), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n473), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT84), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n466), .A2(new_n472), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G190), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT84), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n473), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n491), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n466), .A2(new_n472), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT21), .A4(G169), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n466), .B2(new_n472), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n491), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n466), .A2(new_n472), .A3(new_n309), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n457), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT85), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT6), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n513), .A2(new_n482), .A3(G107), .ZN(new_n514));
  XNOR2_X1  g0314(.A(G97), .B(G107), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n516), .A2(new_n208), .B1(new_n202), .B2(new_n320), .ZN(new_n517));
  XNOR2_X1  g0317(.A(KEYINPUT71), .B(G107), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n323), .B2(new_n324), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n254), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n256), .A2(G97), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n476), .B2(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n292), .A2(new_n464), .A3(KEYINPUT4), .A4(G244), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n481), .A3(new_n525), .ZN(new_n526));
  AND4_X1   g0326(.A1(new_n280), .A2(new_n282), .A3(new_n286), .A4(new_n288), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT4), .B1(new_n527), .B2(G244), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n295), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n468), .A2(new_n467), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n530), .A2(G257), .A3(new_n272), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n529), .A2(new_n309), .A3(new_n471), .A4(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n471), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n289), .B2(new_n216), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(new_n481), .A3(new_n524), .A4(new_n525), .ZN(new_n537));
  AOI211_X1 g0337(.A(new_n534), .B(new_n531), .C1(new_n537), .C2(new_n295), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n523), .B(new_n533), .C1(new_n538), .C2(G169), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n531), .B1(new_n537), .B2(new_n295), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n540), .A2(KEYINPUT80), .A3(new_n471), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT80), .B1(new_n540), .B2(new_n471), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n541), .A2(new_n542), .A3(new_n297), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n538), .A2(KEYINPUT81), .A3(G190), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n529), .A2(G190), .A3(new_n471), .A4(new_n532), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT81), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n523), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n539), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT23), .B1(new_n422), .B2(new_n208), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n435), .A2(G20), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n292), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT86), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n208), .A2(KEYINPUT23), .A3(G107), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(G116), .B2(new_n248), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT24), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT22), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT87), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n559), .A2(KEYINPUT86), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n292), .A2(KEYINPUT87), .A3(new_n552), .A4(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n557), .A2(new_n558), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n563), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT24), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n254), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n530), .A2(G264), .A3(new_n272), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n471), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n292), .A2(G257), .A3(G1698), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G294), .ZN(new_n573));
  INV_X1    g0373(.A(G250), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(new_n289), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n571), .B1(new_n295), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n416), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G200), .B2(new_n576), .ZN(new_n578));
  INV_X1    g0378(.A(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT25), .B1(new_n257), .B2(new_n579), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(new_n579), .B2(new_n475), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n569), .A2(new_n578), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n576), .A2(new_n309), .ZN(new_n586));
  INV_X1    g0386(.A(new_n571), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n575), .A2(new_n295), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(G169), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n432), .B1(new_n564), .B2(new_n567), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n586), .B(new_n591), .C1(new_n592), .C2(new_n583), .ZN(new_n593));
  NOR2_X1   g0393(.A1(G87), .A2(G97), .ZN(new_n594));
  NAND3_X1  g0394(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n518), .A2(new_n594), .B1(new_n208), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n247), .B2(new_n482), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n315), .A2(G20), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n280), .A3(new_n282), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n254), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n257), .B1(new_n434), .B2(new_n439), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n440), .A2(new_n476), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n467), .A2(new_n574), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n272), .ZN(new_n607));
  INV_X1    g0407(.A(new_n467), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n272), .A2(G274), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(G1698), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G116), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n611), .B(new_n612), .C1(new_n289), .C2(new_n389), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n295), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n604), .A2(new_n605), .B1(new_n614), .B2(new_n309), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n295), .ZN(new_n616));
  INV_X1    g0416(.A(new_n610), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n590), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n297), .B1(new_n616), .B2(new_n617), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n618), .A2(new_n416), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n476), .A2(G87), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(new_n624), .A3(new_n604), .A4(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n585), .A2(new_n593), .A3(new_n620), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n550), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n456), .A2(new_n512), .A3(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n539), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n602), .A2(new_n603), .A3(new_n625), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT88), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n602), .A2(KEYINPUT88), .A3(new_n603), .A4(new_n625), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n621), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n624), .B1(new_n635), .B2(KEYINPUT89), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT89), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n637), .B(new_n621), .C1(new_n633), .C2(new_n634), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n630), .B(new_n620), .C1(new_n636), .C2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n639), .A2(KEYINPUT90), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT90), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n626), .A2(new_n620), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n643), .A2(new_n640), .A3(new_n539), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n636), .A2(new_n638), .ZN(new_n646));
  INV_X1    g0446(.A(new_n620), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR3_X1    g0448(.A1(new_n541), .A2(new_n542), .A3(new_n297), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n630), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n509), .A2(new_n593), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n648), .A2(new_n651), .A3(new_n585), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n620), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n456), .B1(new_n645), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n370), .B1(new_n358), .B2(new_n352), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT18), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n370), .B(new_n373), .C1(new_n358), .C2(new_n352), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n447), .A2(new_n450), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n420), .B1(new_n414), .B2(new_n405), .ZN(new_n661));
  INV_X1    g0461(.A(new_n383), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n657), .B(new_n658), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n311), .B1(new_n663), .B2(new_n307), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n655), .A2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(G13), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n666), .A2(G1), .A3(G20), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT91), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT92), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n671));
  INV_X1    g0471(.A(G213), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(G343), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n512), .B1(new_n491), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n674), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n507), .A2(new_n499), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n593), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n676), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n676), .B1(new_n592), .B2(new_n583), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(new_n593), .A3(new_n585), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n507), .A2(new_n674), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT93), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n685), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n674), .B(KEYINPUT94), .Z(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n681), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n211), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n518), .A2(new_n478), .A3(new_n594), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n225), .B2(new_n696), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT95), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n690), .B1(new_n645), .B2(new_n654), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n585), .B(new_n620), .C1(new_n636), .C2(new_n638), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n509), .B2(new_n593), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n647), .B1(new_n707), .B2(new_n651), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n640), .B1(new_n643), .B2(new_n539), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n639), .B2(new_n640), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n676), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G330), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n512), .A2(new_n628), .A3(new_n690), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n540), .A2(new_n576), .A3(new_n614), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n494), .A2(G179), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT30), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n589), .A2(new_n618), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n505), .A3(new_n720), .A4(new_n540), .ZN(new_n721));
  NOR4_X1   g0521(.A1(new_n494), .A2(new_n576), .A3(new_n614), .A4(G179), .ZN(new_n722));
  INV_X1    g0522(.A(new_n538), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n718), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n690), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n718), .A2(new_n721), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n722), .A2(new_n723), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT31), .B1(new_n729), .B2(new_n676), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n714), .B1(new_n715), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n713), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n702), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(new_n678), .A2(G330), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT97), .Z(new_n736));
  NOR2_X1   g0536(.A1(new_n666), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n207), .B1(new_n737), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n736), .B(new_n679), .C1(new_n695), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n695), .A2(new_n739), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT98), .Z(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n253), .B1(G20), .B2(new_n590), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n208), .A2(G179), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G190), .A2(G200), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT100), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT100), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G329), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n208), .A2(new_n309), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n747), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n283), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n754), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(new_n416), .A3(G200), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(G322), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n746), .A2(new_n416), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n762), .A2(G303), .B1(new_n764), .B2(G283), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n753), .A2(new_n760), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n754), .A2(G200), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT99), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n416), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n416), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n208), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n769), .A2(G326), .B1(G294), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT102), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n768), .A2(G190), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n766), .B(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n771), .A2(new_n482), .ZN(new_n779));
  INV_X1    g0579(.A(new_n759), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n780), .A2(new_n314), .B1(new_n215), .B2(new_n755), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n779), .B(new_n781), .C1(new_n769), .C2(G50), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n752), .A2(G159), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT32), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n783), .A2(KEYINPUT32), .B1(G68), .B2(new_n775), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n292), .B1(new_n761), .B2(new_n435), .C1(new_n579), .C2(new_n763), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT101), .Z(new_n787));
  NAND4_X1  g0587(.A1(new_n782), .A2(new_n784), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n745), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n744), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n694), .A2(new_n283), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n478), .B2(new_n694), .ZN(new_n795));
  INV_X1    g0595(.A(new_n331), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n694), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G45), .B2(new_n226), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n243), .A2(new_n273), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n743), .B(new_n789), .C1(new_n793), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n792), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n678), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n740), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  INV_X1    g0605(.A(new_n430), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT73), .B1(new_n448), .B2(new_n449), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n674), .A2(new_n448), .ZN(new_n808));
  AND4_X1   g0608(.A1(new_n450), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n808), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n454), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n703), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n811), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n690), .B(new_n813), .C1(new_n645), .C2(new_n654), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n732), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n741), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n744), .A2(new_n790), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n742), .B1(G77), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G283), .A2(new_n775), .B1(new_n769), .B2(G303), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n763), .A2(new_n435), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n823), .B(new_n779), .C1(G107), .C2(new_n762), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n752), .A2(G311), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n283), .B1(new_n755), .B2(new_n478), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G294), .B2(new_n759), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n755), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n759), .A2(G143), .B1(G159), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n769), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  INV_X1    g0633(.A(new_n775), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n830), .B1(new_n831), .B2(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n763), .A2(new_n315), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n796), .B1(new_n259), .B2(new_n761), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n838), .B(new_n839), .C1(G58), .C2(new_n772), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n837), .B(new_n840), .C1(new_n841), .C2(new_n751), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n835), .A2(new_n836), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n828), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n821), .B1(new_n844), .B2(new_n744), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n813), .B2(new_n791), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n818), .A2(new_n846), .ZN(G384));
  NOR2_X1   g0647(.A1(new_n737), .A2(new_n207), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n318), .B1(new_n319), .B2(new_n320), .C1(new_n344), .C2(new_n315), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n432), .B1(new_n849), .B2(new_n335), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n352), .B1(new_n850), .B2(new_n375), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n670), .A2(new_n673), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n384), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n347), .A2(new_n353), .A3(new_n379), .ZN(new_n855));
  INV_X1    g0655(.A(new_n370), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n851), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT37), .B1(new_n857), .B2(new_n853), .ZN(new_n858));
  INV_X1    g0658(.A(new_n852), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n354), .A2(new_n359), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT37), .B1(new_n376), .B2(new_n379), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n371), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT104), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n854), .A2(KEYINPUT104), .A3(KEYINPUT38), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n855), .A2(new_n381), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n376), .A2(KEYINPUT17), .A3(new_n379), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n657), .A2(new_n868), .A3(new_n869), .A4(new_n658), .ZN(new_n870));
  INV_X1    g0670(.A(new_n860), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n656), .A2(new_n855), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(new_n860), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n371), .A2(new_n860), .A3(new_n861), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n866), .A2(new_n867), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n676), .A2(new_n414), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n415), .A2(new_n420), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n420), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n414), .B(new_n676), .C1(new_n405), .C2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n811), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n724), .A2(new_n725), .A3(new_n674), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n730), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n715), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT40), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n885), .A2(new_n888), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n863), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n854), .B2(new_n863), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n893), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n456), .A2(new_n888), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n714), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT39), .B1(new_n877), .B2(new_n878), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n866), .A2(new_n867), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT39), .B1(new_n895), .B2(new_n896), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n415), .A2(new_n676), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n882), .A2(new_n884), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n659), .A2(new_n676), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n909), .B1(new_n814), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n854), .A2(new_n863), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n878), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n864), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n657), .A2(new_n658), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n912), .A2(new_n915), .B1(new_n916), .B2(new_n852), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n705), .A2(new_n712), .A3(new_n456), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n664), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n848), .B1(new_n901), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n921), .B2(new_n901), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n215), .A2(new_n225), .A3(new_n316), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n259), .B2(G68), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n925), .A2(new_n207), .A3(G13), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT103), .Z(new_n927));
  INV_X1    g0727(.A(KEYINPUT36), .ZN(new_n928));
  INV_X1    g0728(.A(new_n516), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n478), .B(new_n224), .C1(new_n929), .C2(KEYINPUT35), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(KEYINPUT35), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n927), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n923), .A2(new_n933), .ZN(G367));
  NAND3_X1  g0734(.A1(new_n676), .A2(new_n633), .A3(new_n634), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n648), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n620), .B2(new_n935), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(new_n802), .ZN(new_n938));
  INV_X1    g0738(.A(new_n797), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n236), .ZN(new_n940));
  INV_X1    g0740(.A(new_n440), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n793), .B1(new_n941), .B2(new_n211), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n742), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(G143), .A2(new_n769), .B1(new_n775), .B2(G159), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n215), .A2(new_n763), .B1(new_n314), .B2(new_n761), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G68), .B2(new_n772), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n292), .B1(new_n755), .B2(new_n259), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G150), .B2(new_n759), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n752), .A2(G137), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n944), .A2(new_n946), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(G303), .ZN(new_n951));
  INV_X1    g0751(.A(G283), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n780), .A2(new_n951), .B1(new_n755), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n763), .A2(new_n482), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n771), .A2(new_n518), .ZN(new_n955));
  NOR4_X1   g0755(.A1(new_n953), .A2(new_n796), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(G294), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n956), .B1(new_n957), .B2(new_n834), .C1(new_n756), .C2(new_n831), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n762), .A2(KEYINPUT46), .A3(G116), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT46), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n761), .B2(new_n478), .ZN(new_n961));
  INV_X1    g0761(.A(G317), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n959), .B(new_n961), .C1(new_n751), .C2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n950), .B1(new_n958), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT47), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n943), .B1(new_n965), .B2(new_n744), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n938), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n651), .B1(new_n548), .B2(new_n690), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n690), .A2(new_n539), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n692), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n968), .B1(new_n692), .B2(new_n971), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n692), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n689), .A2(new_n691), .A3(new_n971), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n972), .A2(new_n973), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(new_n686), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n686), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n685), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n679), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n688), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n733), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n695), .B(KEYINPUT41), .Z(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n739), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n971), .A2(new_n685), .A3(new_n688), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT42), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n593), .B1(new_n649), .B2(new_n650), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(new_n630), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n992), .A2(new_n993), .B1(new_n690), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n937), .B(KEYINPUT43), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n996), .A2(KEYINPUT105), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT105), .B1(new_n996), .B2(new_n997), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT106), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n686), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n971), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT106), .B1(new_n1004), .B2(new_n971), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n967), .B1(new_n989), .B2(new_n1011), .ZN(G387));
  XNOR2_X1  g0812(.A(new_n983), .B(new_n688), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n733), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n733), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n985), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(new_n1016), .A3(new_n695), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n794), .A2(new_n697), .B1(new_n579), .B2(new_n694), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n233), .A2(G45), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT107), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n246), .A2(new_n259), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n698), .B(new_n273), .C1(new_n315), .C2(new_n202), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n797), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1018), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n743), .B1(new_n1025), .B2(new_n793), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n685), .B2(new_n802), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n780), .A2(new_n259), .B1(new_n755), .B2(new_n315), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n215), .A2(new_n761), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1028), .A2(new_n331), .A3(new_n1029), .A4(new_n954), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G159), .A2(new_n769), .B1(new_n775), .B2(new_n246), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n440), .A2(new_n772), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n752), .A2(G150), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n752), .A2(G326), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n796), .B1(G116), .B2(new_n764), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n771), .A2(new_n952), .B1(new_n761), .B2(new_n957), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n769), .A2(G322), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n759), .A2(G317), .B1(G303), .B2(new_n829), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n834), .C2(new_n756), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1035), .B(new_n1036), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1027), .B1(new_n744), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1013), .B2(new_n739), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1017), .A2(new_n1049), .ZN(G393));
  OAI221_X1 g0850(.A(new_n793), .B1(new_n482), .B2(new_n211), .C1(new_n939), .C2(new_n240), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n742), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n971), .A2(new_n802), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n769), .A2(G317), .B1(G311), .B2(new_n759), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  OAI221_X1 g0855(.A(new_n283), .B1(new_n755), .B2(new_n957), .C1(new_n579), .C2(new_n763), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n771), .A2(new_n478), .B1(new_n761), .B2(new_n952), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n752), .C2(G322), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1055), .B(new_n1058), .C1(new_n951), .C2(new_n834), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT110), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n769), .A2(G150), .B1(G159), .B2(new_n759), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT51), .Z(new_n1063));
  NAND2_X1  g0863(.A1(new_n775), .A2(G50), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n771), .A2(new_n202), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n823), .B(new_n1065), .C1(G68), .C2(new_n762), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n796), .B1(new_n245), .B2(new_n755), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G143), .B2(new_n752), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1061), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1052), .B(new_n1053), .C1(new_n744), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n979), .A2(new_n980), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n985), .A2(new_n1015), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n696), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n979), .A2(KEYINPUT108), .A3(new_n980), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n978), .A2(KEYINPUT108), .A3(new_n686), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1014), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1072), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT109), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT109), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1076), .A2(new_n1083), .A3(new_n1078), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n739), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1080), .A2(new_n1085), .ZN(G390));
  AOI21_X1  g0886(.A(new_n743), .B1(new_n245), .B2(new_n819), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n761), .A2(new_n833), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT53), .ZN(new_n1089));
  INV_X1    g0889(.A(G128), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n831), .B2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT54), .B(G143), .Z(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT111), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n752), .A2(G125), .B1(new_n829), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n772), .A2(G159), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n764), .A2(G50), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n283), .B1(new_n759), .B2(G132), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1091), .B(new_n1098), .C1(G137), .C2(new_n775), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT112), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G283), .A2(new_n769), .B1(new_n775), .B2(new_n422), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n838), .B(new_n1065), .C1(G87), .C2(new_n762), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n752), .A2(G294), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n283), .B1(new_n780), .B2(new_n478), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G97), .B2(new_n829), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(KEYINPUT112), .B2(new_n1099), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1087), .B1(new_n745), .B2(new_n1108), .C1(new_n905), .C2(new_n791), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT113), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n653), .A2(new_n620), .A3(new_n710), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n674), .A3(new_n813), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n911), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n906), .B1(new_n1113), .B2(new_n908), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n880), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n912), .A2(new_n906), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n905), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n714), .B1(new_n715), .B2(new_n887), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(new_n885), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n732), .A2(new_n813), .A3(new_n908), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1115), .B(new_n1121), .C1(new_n905), .C2(new_n1116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(new_n738), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1110), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n456), .A2(new_n1118), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n919), .A2(new_n664), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1121), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n908), .B1(new_n1118), .B2(new_n813), .ZN(new_n1129));
  OR3_X1    g0929(.A1(new_n1128), .A2(new_n1113), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n814), .A2(new_n911), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n908), .B1(new_n732), .B2(new_n813), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n1119), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1127), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1123), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1120), .A2(new_n1122), .A3(new_n1134), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n695), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1125), .A2(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(new_n1127), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n912), .A2(new_n915), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n916), .A2(new_n852), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n906), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n903), .B2(new_n904), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n714), .B1(new_n897), .B2(new_n890), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT117), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n859), .A2(new_n265), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT116), .Z(new_n1150));
  NAND2_X1  g0950(.A1(new_n313), .A2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1150), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n307), .A2(new_n312), .A3(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1152), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1148), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1152), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1151), .A2(new_n1154), .A3(new_n1152), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(KEYINPUT117), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1147), .A2(new_n1163), .A3(new_n892), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1147), .B2(new_n892), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1146), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1165), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n889), .B1(new_n914), .B2(new_n864), .ZN(new_n1169));
  OAI21_X1  g0969(.A(G330), .B1(new_n1169), .B2(KEYINPUT40), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n893), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1147), .A2(new_n1163), .A3(new_n892), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n918), .A3(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1140), .A2(new_n1137), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT118), .B1(new_n1174), .B2(KEYINPUT57), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n696), .B1(new_n1174), .B2(KEYINPUT57), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT118), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1175), .A2(new_n1176), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1163), .A2(new_n790), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n741), .B1(G50), .B2(new_n820), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n796), .A2(G41), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n941), .B2(new_n755), .C1(new_n952), .C2(new_n751), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n831), .A2(new_n478), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n834), .A2(new_n482), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G107), .A2(new_n759), .B1(new_n772), .B2(G68), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n764), .A2(G58), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n215), .C2(new_n761), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n259), .B1(G33), .B2(G41), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1194), .B(new_n1195), .C1(new_n1186), .C2(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n752), .A2(G124), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n270), .B(new_n271), .C1(new_n763), .C2(new_n319), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n769), .A2(G125), .B1(G150), .B2(new_n772), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT115), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1093), .A2(new_n762), .B1(G128), .B2(new_n759), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT114), .Z(new_n1203));
  AOI22_X1  g1003(.A1(new_n775), .A2(G132), .B1(G137), .B2(new_n829), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1198), .B(new_n1199), .C1(new_n1205), .C2(KEYINPUT59), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1197), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1185), .B1(new_n1209), .B2(new_n744), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1184), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1178), .B2(new_n739), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1183), .A2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT119), .ZN(G375));
  NAND3_X1  g1015(.A1(new_n1130), .A2(new_n1127), .A3(new_n1133), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1135), .A2(new_n988), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n738), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n909), .A2(new_n790), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n742), .B1(G68), .B2(new_n820), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G116), .A2(new_n775), .B1(new_n769), .B2(G294), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n283), .B1(new_n755), .B2(new_n518), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n202), .A2(new_n763), .B1(new_n761), .B2(new_n482), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(G283), .C2(new_n759), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n752), .A2(G303), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1221), .A2(new_n1032), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n775), .A2(new_n1093), .B1(G137), .B2(new_n759), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n841), .B2(new_n831), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT120), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n796), .B1(new_n833), .B2(new_n755), .C1(new_n751), .C2(new_n1090), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1191), .B1(new_n319), .B2(new_n761), .C1(new_n259), .C2(new_n771), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1226), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1220), .B1(new_n1233), .B2(new_n744), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1218), .B1(new_n1219), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1217), .A2(new_n1235), .ZN(G381));
  INV_X1    g1036(.A(KEYINPUT119), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1214), .B(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G393), .A2(G396), .ZN(new_n1240));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(G387), .A2(G390), .A3(new_n1242), .A4(G381), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n1239), .A3(new_n1243), .ZN(G407));
  NAND2_X1  g1044(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(new_n1245), .C2(G343), .ZN(G409));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n672), .A2(G343), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1174), .A2(new_n988), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT121), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n738), .B1(new_n1178), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1167), .A2(new_n1173), .A3(KEYINPUT121), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1212), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT122), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1249), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI211_X1 g1055(.A(KEYINPUT122), .B(new_n1212), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1239), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1183), .A2(G378), .A3(new_n1213), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1248), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  OR3_X1    g1060(.A1(new_n1216), .A2(KEYINPUT123), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT123), .B1(new_n1216), .B2(new_n1260), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1216), .A2(new_n1260), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1134), .A2(new_n696), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1235), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT124), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G384), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(G384), .A2(new_n1267), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1266), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1265), .A2(KEYINPUT124), .A3(new_n1241), .A4(new_n1235), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1248), .A2(G2897), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1273), .B(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1247), .B1(new_n1259), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1248), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1249), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1164), .A2(new_n1146), .A3(new_n1166), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n918), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1250), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n739), .A3(new_n1252), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1211), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1280), .B1(new_n1285), .B2(KEYINPUT122), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G378), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1183), .A2(G378), .A3(new_n1213), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1279), .B(new_n1273), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .A3(new_n1279), .A4(new_n1273), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(KEYINPUT126), .B(new_n1247), .C1(new_n1259), .C2(new_n1275), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1278), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n804), .B1(new_n1017), .B2(new_n1049), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1240), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1011), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n986), .A2(new_n988), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n738), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1301), .A2(new_n1303), .B1(new_n938), .B2(new_n966), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1304), .A2(G390), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(G387), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1300), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(G390), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(G387), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1299), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(KEYINPUT127), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1297), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1308), .A2(new_n1247), .A3(new_n1311), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1315), .B(KEYINPUT125), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1259), .A2(new_n1275), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1259), .A2(KEYINPUT63), .A3(new_n1273), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1290), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1314), .A2(new_n1321), .ZN(G405));
  AOI21_X1  g1122(.A(new_n1239), .B1(new_n1183), .B2(new_n1213), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1245), .A2(new_n1273), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1273), .B1(new_n1245), .B2(new_n1324), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1312), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1273), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(G375), .A2(G378), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(new_n1323), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1331), .A2(new_n1311), .A3(new_n1308), .A4(new_n1325), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1328), .A2(new_n1332), .ZN(G402));
endmodule


