//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n209), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n209), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  INV_X1    g0021(.A(new_n201), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n221), .B(new_n227), .C1(KEYINPUT1), .C2(new_n216), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n218), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n225), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  OAI22_X1  g0051(.A1(new_n248), .A2(new_n250), .B1(new_n207), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT15), .B(G87), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n207), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n247), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(KEYINPUT72), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(KEYINPUT72), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G77), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n247), .B1(new_n206), .B2(G20), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(G77), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G107), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G238), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n267), .B1(new_n268), .B2(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n272), .A2(KEYINPUT69), .A3(new_n225), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  AND2_X1   g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n206), .A2(new_n282), .B1(new_n275), .B2(new_n276), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n275), .B2(new_n276), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n283), .A2(G244), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n264), .B(new_n291), .C1(G179), .C2(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(G200), .ZN(new_n293));
  INV_X1    g0093(.A(new_n263), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n257), .B2(new_n258), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n279), .A2(G190), .A3(new_n288), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n260), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n202), .ZN(new_n299));
  INV_X1    g0099(.A(new_n262), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n202), .ZN(new_n301));
  INV_X1    g0101(.A(new_n247), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT70), .A2(G58), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT8), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(new_n207), .A3(G33), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n249), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n285), .A2(new_n287), .ZN(new_n309));
  INV_X1    g0109(.A(G226), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n275), .A2(new_n276), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n286), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n265), .A2(G222), .A3(new_n266), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT67), .B(G223), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n314), .B1(new_n251), .B2(new_n265), .C1(new_n269), .C2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT68), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT69), .B1(new_n272), .B2(new_n225), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n275), .A2(new_n274), .A3(new_n276), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n316), .B2(new_n317), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n313), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n308), .B1(new_n324), .B2(new_n290), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n325), .A2(KEYINPUT71), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT71), .B1(new_n325), .B2(new_n327), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n292), .B(new_n297), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  OAI211_X1 g0132(.A(G232), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n265), .A2(new_n335), .A3(G232), .A4(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(G226), .B(new_n266), .C1(new_n331), .C2(new_n332), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G97), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n321), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n309), .B1(new_n270), .B2(new_n312), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT13), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n343), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n340), .B1(new_n336), .B2(new_n334), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n345), .B(new_n346), .C1(new_n347), .C2(new_n321), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(G169), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT79), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n344), .A2(new_n348), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT14), .B1(new_n354), .B2(new_n290), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n349), .A2(KEYINPUT79), .A3(new_n350), .A4(G169), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(G179), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n353), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G68), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n298), .A2(KEYINPUT78), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT12), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT78), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n260), .B2(G68), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n363), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n364), .A2(new_n365), .B1(G68), .B2(new_n262), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n249), .A2(G50), .B1(G20), .B2(new_n359), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n251), .B2(new_n254), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n247), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT76), .B(KEYINPUT11), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n247), .A3(new_n370), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(KEYINPUT77), .A3(new_n373), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n366), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n358), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n378), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n349), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n354), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT82), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  INV_X1    g0189(.A(G223), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n266), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n310), .A2(G1698), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n392), .C1(new_n331), .C2(new_n332), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n321), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G232), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n309), .B1(new_n395), .B2(new_n312), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n388), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n389), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n278), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n283), .A2(G232), .B1(new_n285), .B2(new_n287), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(KEYINPUT82), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(G169), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(G179), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT83), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n399), .A2(KEYINPUT82), .A3(new_n400), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT82), .B1(new_n399), .B2(new_n400), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n290), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT83), .ZN(new_n409));
  INV_X1    g0209(.A(new_n404), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT3), .ZN(new_n414));
  INV_X1    g0214(.A(G33), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(KEYINPUT3), .A2(G33), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n207), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n416), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n417), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n359), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G58), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n359), .ZN(new_n424));
  OAI21_X1  g0224(.A(G20), .B1(new_n424), .B2(new_n201), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n249), .A2(G159), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n413), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n247), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n331), .A2(new_n332), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT7), .B1(new_n430), .B2(new_n207), .ZN(new_n431));
  INV_X1    g0231(.A(new_n421), .ZN(new_n432));
  OAI21_X1  g0232(.A(G68), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n433), .A2(KEYINPUT16), .A3(new_n426), .A4(new_n425), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT80), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n422), .A2(new_n427), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(KEYINPUT80), .A3(KEYINPUT16), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n429), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n304), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n260), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n262), .B2(new_n440), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT81), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT18), .B1(new_n412), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n428), .A2(new_n247), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n434), .A2(new_n435), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT80), .B1(new_n437), .B2(KEYINPUT16), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n442), .B(KEYINPUT81), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n411), .A4(new_n405), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n383), .B1(new_n406), .B2(new_n407), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n399), .A2(new_n381), .A3(new_n400), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(new_n457), .A3(new_n451), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n445), .A2(KEYINPUT17), .A3(new_n457), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n446), .A2(new_n454), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT9), .ZN(new_n463));
  OAI211_X1 g0263(.A(KEYINPUT73), .B(new_n463), .C1(new_n301), .C2(new_n307), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n308), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n464), .B(new_n467), .C1(new_n323), .C2(new_n383), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT74), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n323), .A2(G190), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT10), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(KEYINPUT10), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n470), .A2(KEYINPUT10), .ZN(new_n474));
  INV_X1    g0274(.A(new_n471), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n468), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NOR4_X1   g0277(.A1(new_n330), .A2(new_n387), .A3(new_n462), .A4(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT94), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G250), .A2(G1698), .ZN(new_n480));
  INV_X1    g0280(.A(G257), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(G1698), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(new_n265), .B1(G33), .B2(G294), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n479), .B1(new_n483), .B2(new_n321), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(G1698), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(G250), .B2(G1698), .ZN(new_n486));
  INV_X1    g0286(.A(G294), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n486), .A2(new_n430), .B1(new_n415), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n278), .A3(KEYINPUT94), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT5), .B(G41), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n281), .A2(G1), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n491), .B1(new_n275), .B2(new_n276), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n206), .A2(G45), .ZN(new_n493));
  OR2_X1    g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n492), .A2(G264), .B1(new_n496), .B2(new_n285), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n484), .A2(new_n489), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT95), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT95), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n484), .A2(new_n497), .A3(new_n489), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n290), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n488), .A2(new_n278), .B1(new_n492), .B2(G264), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(new_n285), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n326), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n265), .A2(new_n207), .A3(G87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT22), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT22), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n265), .A2(new_n509), .A3(new_n207), .A4(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n415), .A2(new_n512), .A3(G20), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n207), .A2(G107), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n514), .A2(KEYINPUT23), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(KEYINPUT23), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT24), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n511), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n302), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G13), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(G1), .ZN(new_n524));
  OR2_X1    g0324(.A1(KEYINPUT93), .A2(KEYINPUT25), .ZN(new_n525));
  NAND2_X1  g0325(.A1(KEYINPUT93), .A2(KEYINPUT25), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n514), .A2(new_n524), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n514), .A2(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n206), .A2(G33), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n260), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n247), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI221_X1 g0332(.A(new_n527), .B1(new_n528), .B2(new_n526), .C1(new_n532), .C2(new_n268), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n502), .A2(new_n506), .B1(new_n522), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n499), .A2(new_n381), .A3(new_n501), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n505), .A2(new_n383), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n519), .A2(new_n521), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n533), .B1(new_n539), .B2(new_n247), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT96), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n538), .A2(KEYINPUT96), .A3(new_n540), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n535), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G264), .A2(G1698), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n481), .B2(G1698), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n265), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(KEYINPUT91), .A2(G303), .ZN(new_n549));
  NOR2_X1   g0349(.A1(KEYINPUT91), .A2(G303), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n416), .B(new_n417), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT92), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n548), .A2(KEYINPUT92), .A3(new_n551), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n278), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n495), .ZN(new_n557));
  NOR2_X1   g0357(.A1(KEYINPUT5), .A2(G41), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n491), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n311), .ZN(new_n560));
  INV_X1    g0360(.A(G270), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n504), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n298), .A2(new_n512), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n531), .A2(G116), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G283), .ZN(new_n567));
  AND2_X1   g0367(.A1(KEYINPUT85), .A2(G97), .ZN(new_n568));
  NOR2_X1   g0368(.A1(KEYINPUT85), .A2(G97), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n207), .B(new_n567), .C1(new_n570), .C2(G33), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n246), .A2(new_n225), .B1(G20), .B2(new_n512), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT20), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OR2_X1    g0373(.A1(KEYINPUT85), .A2(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(KEYINPUT85), .A2(G97), .ZN(new_n575));
  AOI21_X1  g0375(.A(G33), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n567), .A2(new_n207), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT20), .B(new_n572), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n565), .B(new_n566), .C1(new_n573), .C2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n564), .A2(new_n580), .A3(G169), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n321), .B1(new_n552), .B2(new_n553), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n326), .B(new_n562), .C1(new_n584), .C2(new_n555), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n580), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n566), .A2(new_n565), .ZN(new_n587));
  INV_X1    g0387(.A(new_n573), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n578), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n556), .A2(G190), .A3(new_n563), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n562), .B1(new_n584), .B2(new_n555), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n589), .B(new_n590), .C1(new_n383), .C2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n564), .A2(new_n580), .A3(KEYINPUT21), .A4(G169), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n583), .A2(new_n586), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(G244), .B(new_n266), .C1(new_n331), .C2(new_n332), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n567), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n278), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n504), .B1(new_n560), .B2(new_n481), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(G190), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n249), .A2(G77), .ZN(new_n605));
  OR2_X1    g0405(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n606));
  NAND2_X1  g0406(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n607));
  AOI21_X1  g0407(.A(G107), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n574), .A2(new_n575), .ZN(new_n609));
  AND2_X1   g0409(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n610));
  NOR2_X1   g0410(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g0412(.A(G97), .B(G107), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n608), .A2(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n605), .B1(new_n614), .B2(new_n207), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n268), .B1(new_n420), .B2(new_n421), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n247), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n260), .A2(G97), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n531), .B2(G97), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n604), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n602), .A2(KEYINPUT86), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT86), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n504), .B(new_n622), .C1(new_n560), .C2(new_n481), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n601), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT87), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n383), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n601), .A2(new_n621), .A3(KEYINPUT87), .A4(new_n623), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(G244), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n629));
  OAI211_X1 g0429(.A(G238), .B(new_n266), .C1(new_n331), .C2(new_n332), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n630), .C1(new_n415), .C2(new_n512), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n278), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n272), .A2(new_n225), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n493), .A2(G250), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT88), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n311), .A2(new_n636), .A3(G250), .A4(new_n493), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n635), .A2(new_n637), .B1(new_n491), .B2(new_n285), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n632), .A2(new_n638), .A3(G190), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT90), .ZN(new_n640));
  INV_X1    g0440(.A(new_n253), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(new_n260), .ZN(new_n642));
  INV_X1    g0442(.A(G87), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n530), .A2(new_n643), .A3(new_n247), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT19), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n207), .B1(new_n339), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n574), .A2(new_n268), .A3(new_n575), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n643), .A2(KEYINPUT89), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G87), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n646), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n265), .A2(new_n207), .A3(G68), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n645), .B1(new_n570), .B2(new_n254), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n642), .B(new_n644), .C1(new_n655), .C2(new_n247), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n632), .A2(new_n638), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G200), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT90), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n632), .A2(new_n638), .A3(new_n659), .A4(G190), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n640), .A2(new_n656), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n642), .B1(new_n655), .B2(new_n247), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n531), .A2(new_n641), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n657), .A2(new_n290), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n632), .A2(new_n638), .A3(new_n326), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n326), .A2(new_n601), .A3(new_n621), .A4(new_n623), .ZN(new_n669));
  INV_X1    g0469(.A(new_n619), .ZN(new_n670));
  AND2_X1   g0470(.A1(G97), .A2(G107), .ZN(new_n671));
  NOR2_X1   g0471(.A1(G97), .A2(G107), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n606), .B(new_n607), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n268), .B1(new_n610), .B2(new_n611), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n570), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G20), .ZN(new_n676));
  OAI21_X1  g0476(.A(G107), .B1(new_n431), .B2(new_n432), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(new_n605), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n670), .B1(new_n678), .B2(new_n247), .ZN(new_n679));
  AOI21_X1  g0479(.A(G169), .B1(new_n601), .B2(new_n603), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n669), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NOR4_X1   g0481(.A1(new_n594), .A2(new_n628), .A3(new_n668), .A4(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n478), .A2(new_n545), .A3(new_n682), .ZN(G372));
  NOR3_X1   g0483(.A1(new_n628), .A2(new_n668), .A3(new_n681), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n586), .A2(new_n593), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n534), .A2(new_n583), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT96), .B1(new_n538), .B2(new_n540), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n538), .A2(KEYINPUT96), .A3(new_n540), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n684), .B(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n667), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT26), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n669), .A2(new_n679), .A3(new_n680), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n668), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n681), .A2(KEYINPUT26), .A3(new_n667), .A4(new_n661), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n478), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n328), .A2(new_n329), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n446), .A2(new_n454), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n379), .A2(new_n292), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n386), .A2(new_n460), .A3(new_n461), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n477), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n697), .A2(new_n704), .ZN(G369));
  NAND2_X1  g0505(.A1(new_n524), .A2(new_n207), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT97), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT27), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n524), .A2(KEYINPUT97), .A3(new_n207), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT98), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT98), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n708), .A2(new_n713), .A3(new_n709), .A4(new_n710), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G213), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n708), .A2(new_n710), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(KEYINPUT27), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n718), .A3(G343), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n545), .B1(new_n540), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n534), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n719), .A2(new_n589), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n594), .B2(KEYINPUT99), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(KEYINPUT99), .B2(new_n594), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n685), .A2(new_n583), .A3(new_n722), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n719), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n685), .B2(new_n583), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n545), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n535), .B2(new_n719), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n729), .A2(new_n734), .ZN(G399));
  NOR3_X1   g0535(.A1(new_n647), .A2(new_n651), .A3(G116), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT100), .ZN(new_n737));
  INV_X1    g0537(.A(new_n219), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G41), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(G1), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n223), .B2(new_n740), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n543), .A2(new_n544), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n682), .A2(new_n744), .A3(new_n534), .A4(new_n719), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n601), .A2(KEYINPUT30), .A3(new_n603), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n503), .A2(new_n632), .A3(new_n638), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT101), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n503), .A2(new_n632), .A3(new_n638), .A4(KEYINPUT101), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n585), .A2(new_n746), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT102), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n750), .A2(G179), .A3(new_n591), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(KEYINPUT102), .A3(new_n749), .A4(new_n746), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n602), .B1(new_n278), .B2(new_n600), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n585), .A2(new_n749), .A3(new_n757), .A4(new_n750), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(G179), .B1(new_n503), .B2(new_n504), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n624), .A2(new_n564), .A3(new_n761), .A4(new_n657), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(KEYINPUT31), .B(new_n730), .C1(new_n756), .C2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n730), .B1(new_n756), .B2(new_n763), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n745), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n768), .A2(G330), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n730), .B1(new_n689), .B2(new_n695), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT103), .B(KEYINPUT29), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT103), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n773), .B2(KEYINPUT29), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n769), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n743), .B1(new_n775), .B2(G1), .ZN(G364));
  NOR2_X1   g0576(.A1(new_n523), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n206), .B1(new_n777), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n739), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n219), .A2(new_n265), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(G116), .B2(new_n219), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n738), .A2(new_n265), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n281), .B2(new_n224), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n244), .A2(G45), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n225), .B1(G20), .B2(new_n290), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n780), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n207), .A2(G190), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n326), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n265), .B1(new_n798), .B2(new_n251), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n326), .A2(G200), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT105), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n796), .A2(KEYINPUT104), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n796), .A2(KEYINPUT104), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n268), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n207), .A2(new_n381), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n797), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n799), .B(new_n805), .C1(G58), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G179), .A2(G200), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n207), .B1(new_n810), .B2(G190), .ZN(new_n811));
  INV_X1    g0611(.A(G97), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n381), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n202), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n814), .A2(G190), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n813), .B(new_n817), .C1(G68), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n801), .A2(new_n806), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n651), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n809), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n802), .A2(new_n803), .A3(new_n810), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G159), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT32), .ZN(new_n827));
  INV_X1    g0627(.A(new_n804), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(G283), .B1(G329), .B2(new_n825), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT106), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  INV_X1    g0631(.A(G322), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n430), .B1(new_n798), .B2(new_n831), .C1(new_n832), .C2(new_n807), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n821), .B2(G303), .ZN(new_n834));
  INV_X1    g0634(.A(G317), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(KEYINPUT33), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(KEYINPUT33), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n818), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n811), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(G294), .B1(G326), .B2(new_n815), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n834), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n823), .A2(new_n827), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n795), .B1(new_n842), .B2(new_n792), .ZN(new_n843));
  INV_X1    g0643(.A(new_n726), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n791), .B(KEYINPUT107), .Z(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(G330), .ZN(new_n847));
  INV_X1    g0647(.A(new_n780), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n726), .B2(new_n727), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(G396));
  INV_X1    g0650(.A(new_n769), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT109), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n264), .A2(new_n730), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT109), .B1(new_n295), .B2(new_n719), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n297), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n292), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n292), .A2(new_n730), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n770), .B(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n780), .B1(new_n851), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n851), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n792), .A2(new_n789), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n848), .B1(new_n251), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n792), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n813), .B1(new_n815), .B2(G303), .ZN(new_n866));
  INV_X1    g0666(.A(G283), .ZN(new_n867));
  INV_X1    g0667(.A(new_n818), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n804), .A2(new_n643), .B1(new_n820), .B2(new_n268), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n824), .A2(new_n831), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n430), .B1(new_n798), .B2(new_n512), .C1(new_n487), .C2(new_n807), .ZN(new_n872));
  NOR4_X1   g0672(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n798), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G143), .A2(new_n808), .B1(new_n874), .B2(G159), .ZN(new_n875));
  INV_X1    g0675(.A(G150), .ZN(new_n876));
  INV_X1    g0676(.A(G137), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n875), .B1(new_n868), .B2(new_n876), .C1(new_n877), .C2(new_n816), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT34), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  INV_X1    g0681(.A(G132), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n265), .B1(new_n423), .B2(new_n811), .C1(new_n824), .C2(new_n882), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n804), .A2(new_n359), .B1(new_n820), .B2(new_n202), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT108), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n873), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n864), .B1(new_n865), .B2(new_n887), .C1(new_n859), .C2(new_n790), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n862), .A2(new_n888), .ZN(G384));
  OR2_X1    g0689(.A1(new_n675), .A2(KEYINPUT35), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n675), .A2(KEYINPUT35), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(G116), .A3(new_n226), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT36), .Z(new_n893));
  OR3_X1    g0693(.A1(new_n223), .A2(new_n251), .A3(new_n424), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n202), .A2(G68), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n206), .B(G13), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n378), .A2(new_n730), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n379), .A2(new_n386), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n378), .B(new_n730), .C1(new_n358), .C2(new_n385), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n768), .A2(new_n859), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT111), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n715), .A2(new_n718), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n442), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n439), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n462), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n439), .A2(new_n906), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n458), .B(new_n907), .C1(new_n412), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n452), .A2(new_n411), .A3(new_n405), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n905), .B1(new_n439), .B2(new_n444), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n913), .A2(new_n914), .A3(new_n458), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT111), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n768), .A2(new_n923), .A3(new_n901), .A4(new_n859), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n903), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n915), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n462), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n458), .B(new_n915), .C1(new_n412), .C2(new_n445), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT37), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n916), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n919), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n926), .B1(new_n934), .B2(new_n921), .ZN(new_n935));
  INV_X1    g0735(.A(new_n902), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n478), .A2(new_n768), .ZN(new_n939));
  OAI21_X1  g0739(.A(G330), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT110), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n699), .A2(new_n905), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n730), .B(new_n858), .C1(new_n689), .C2(new_n695), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n292), .A2(new_n730), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n901), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n917), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n909), .B2(new_n917), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n942), .B(new_n943), .C1(new_n946), .C2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT39), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT38), .B1(new_n929), .B2(new_n932), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n951), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n920), .A2(KEYINPUT39), .A3(new_n921), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n379), .A2(new_n730), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n696), .A2(new_n719), .A3(new_n859), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n958), .A2(new_n857), .B1(new_n899), .B2(new_n900), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n922), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n942), .B1(new_n960), .B2(new_n943), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n772), .A2(new_n478), .A3(new_n774), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n704), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n962), .B(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n941), .A2(new_n965), .B1(new_n206), .B2(new_n777), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n941), .A2(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n897), .B1(new_n966), .B2(new_n967), .ZN(G367));
  INV_X1    g0768(.A(new_n628), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n969), .B(new_n692), .C1(new_n679), .C2(new_n719), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n692), .B2(new_n719), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n733), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n535), .A2(new_n969), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n730), .B1(new_n974), .B2(new_n692), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n972), .B2(KEYINPUT42), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n719), .A2(new_n656), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT112), .Z(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n667), .B2(new_n661), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n667), .B2(new_n978), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n973), .A2(new_n976), .B1(KEYINPUT43), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n721), .A2(new_n728), .A3(new_n971), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n739), .B(KEYINPUT41), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n734), .A2(new_n971), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n734), .A2(new_n971), .ZN(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n988), .A2(new_n729), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n729), .B1(new_n988), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n732), .B1(new_n721), .B2(new_n731), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(new_n728), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n775), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n992), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n986), .B1(new_n997), .B2(new_n775), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n985), .B1(new_n998), .B2(new_n779), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n793), .B1(new_n219), .B2(new_n253), .C1(new_n785), .C2(new_n236), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(new_n780), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n265), .B1(new_n798), .B2(new_n202), .C1(new_n876), .C2(new_n807), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n821), .B2(G58), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n828), .A2(G77), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n877), .C2(new_n824), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n811), .A2(new_n359), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n815), .B2(G143), .ZN(new_n1007));
  INV_X1    g0807(.A(G159), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n868), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n811), .A2(new_n268), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT114), .B(G311), .Z(new_n1011));
  NOR2_X1   g0811(.A1(new_n816), .A2(new_n1011), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G294), .C2(new_n818), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n820), .B2(new_n512), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n821), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n549), .A2(new_n550), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n430), .B1(new_n807), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G283), .B2(new_n874), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n835), .B2(new_n824), .C1(new_n570), .C2(new_n804), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1005), .A2(new_n1009), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT47), .Z(new_n1023));
  OAI221_X1 g0823(.A(new_n1001), .B1(new_n1023), .B2(new_n865), .C1(new_n980), .C2(new_n845), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n999), .A2(new_n1024), .ZN(G387));
  OR2_X1    g0825(.A1(new_n721), .A2(new_n845), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n784), .B1(new_n233), .B2(new_n281), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n737), .B2(new_n781), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n248), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT50), .B1(new_n248), .B2(G50), .ZN(new_n1030));
  AOI21_X1  g0830(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n737), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1028), .A2(new_n1032), .B1(new_n268), .B2(new_n738), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n780), .B1(new_n1033), .B2(new_n794), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1018), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G317), .A2(new_n808), .B1(new_n874), .B2(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n868), .B2(new_n1011), .C1(new_n832), .C2(new_n816), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT48), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n821), .A2(G294), .B1(G283), .B2(new_n839), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n804), .A2(new_n512), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n265), .B(new_n1046), .C1(G326), .C2(new_n825), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n265), .B1(new_n798), .B2(new_n359), .C1(new_n202), .C2(new_n807), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n821), .B2(G77), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n440), .A2(new_n868), .B1(new_n816), .B2(new_n1008), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n811), .A2(new_n253), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n828), .A2(G97), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n825), .A2(G150), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1050), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1048), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1034), .B1(new_n1057), .B2(new_n792), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n995), .A2(new_n779), .B1(new_n1026), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n996), .A2(new_n739), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n995), .A2(new_n775), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(G393));
  OAI21_X1  g0862(.A(new_n996), .B1(new_n992), .B2(new_n993), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n997), .A2(new_n739), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n820), .A2(new_n867), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1065), .B(new_n805), .C1(G322), .C2(new_n825), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n265), .B1(new_n874), .B2(G294), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n512), .B2(new_n811), .C1(new_n868), .C2(new_n1018), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT52), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n816), .A2(new_n835), .B1(new_n807), .B2(new_n831), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1066), .B(new_n1071), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n811), .A2(new_n251), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n265), .B1(new_n798), .B2(new_n248), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(G50), .C2(new_n818), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n808), .A2(G159), .B1(G150), .B2(new_n815), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(KEYINPUT51), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n828), .A2(G87), .B1(G143), .B2(new_n825), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n359), .C2(new_n820), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n865), .B1(new_n1072), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n241), .A2(new_n784), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1083), .B(new_n793), .C1(new_n219), .C2(new_n570), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT115), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n848), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n971), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1082), .B(new_n1087), .C1(new_n1088), .C2(new_n791), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n992), .A2(new_n993), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n779), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1064), .A2(new_n1091), .ZN(G390));
  NAND2_X1  g0892(.A1(new_n769), .A2(new_n478), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(new_n963), .A3(new_n704), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n958), .A2(new_n857), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n768), .A2(G330), .A3(new_n859), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n901), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n768), .A2(G330), .A3(new_n901), .A4(new_n859), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1096), .A3(new_n1100), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1094), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n953), .B(new_n954), .C1(new_n959), .C2(new_n955), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n955), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n946), .A2(new_n921), .A3(new_n1107), .A4(new_n934), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1106), .A2(KEYINPUT116), .A3(new_n1108), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1100), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1100), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1105), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1100), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1106), .A2(KEYINPUT116), .A3(new_n1108), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT116), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n1114), .A3(new_n1104), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n739), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n863), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n839), .A2(G159), .B1(G128), .B2(new_n815), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n877), .B2(new_n868), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n430), .B1(new_n874), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1128), .B1(new_n882), .B2(new_n807), .C1(new_n1129), .C2(new_n824), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1125), .B(new_n1130), .C1(G50), .C2(new_n828), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n820), .A2(new_n876), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n430), .B1(new_n820), .B2(new_n643), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT117), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n804), .A2(new_n359), .B1(new_n487), .B2(new_n824), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n868), .A2(new_n268), .B1(new_n816), .B2(new_n867), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n807), .A2(new_n512), .B1(new_n798), .B2(new_n570), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1073), .A4(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1131), .A2(new_n1133), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n780), .B1(new_n304), .B2(new_n1123), .C1(new_n1140), .C2(new_n865), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n953), .A2(new_n954), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n789), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n779), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1122), .A2(new_n1145), .ZN(G378));
  INV_X1    g0946(.A(KEYINPUT123), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1094), .B(KEYINPUT122), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1121), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n957), .A2(new_n961), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n902), .A2(KEYINPUT111), .B1(new_n921), .B2(new_n920), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT40), .B1(new_n1152), .B2(new_n924), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n937), .A2(G330), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n325), .A2(new_n327), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n703), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n904), .A2(new_n308), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n703), .B(new_n1155), .C1(new_n308), .C2(new_n904), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1153), .A2(new_n1154), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1161), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1160), .B(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n727), .B1(new_n935), .B2(new_n936), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n927), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1151), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1162), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n927), .A2(new_n1166), .A3(new_n1165), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n962), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1147), .B(new_n1148), .C1(new_n1150), .C2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1121), .A2(new_n1149), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT123), .B1(new_n1174), .B2(KEYINPUT57), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n740), .B1(new_n1174), .B2(KEYINPUT57), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n265), .A2(G41), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G50), .B(new_n1178), .C1(new_n415), .C2(new_n280), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n808), .A2(G107), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT118), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n812), .A2(new_n868), .B1(new_n816), .B2(new_n512), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1178), .B1(new_n253), .B2(new_n798), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1006), .B(new_n1184), .C1(new_n821), .C2(G77), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n828), .A2(G58), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n825), .A2(G283), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1179), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT119), .Z(new_n1191));
  AOI22_X1  g0991(.A1(new_n874), .A2(G137), .B1(G125), .B2(new_n815), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n839), .A2(G150), .B1(G132), .B2(new_n818), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n821), .A2(new_n1127), .B1(G128), .B2(new_n808), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT120), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(KEYINPUT120), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1192), .B(new_n1193), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n828), .A2(G159), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n825), .C2(G124), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1191), .B(new_n1202), .C1(new_n1189), .C2(new_n1188), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n865), .B1(new_n1203), .B2(KEYINPUT121), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(KEYINPUT121), .B2(new_n1203), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1205), .B(new_n780), .C1(G50), .C2(new_n1123), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n789), .B2(new_n1162), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1208), .B2(new_n779), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1177), .A2(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1098), .A2(new_n789), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n780), .B1(G68), .B2(new_n1123), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1052), .B1(new_n815), .B2(G294), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n512), .B2(new_n868), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n821), .A2(G97), .B1(new_n825), .B2(G303), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n430), .B1(new_n807), .B2(new_n867), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G107), .B2(new_n874), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1004), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n825), .A2(G128), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1186), .B(new_n1220), .C1(new_n1008), .C2(new_n820), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n815), .A2(G132), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT124), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n265), .B1(new_n798), .B2(new_n876), .C1(new_n877), .C2(new_n807), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n868), .A2(new_n1126), .B1(new_n202), .B2(new_n811), .ZN(new_n1225));
  OR3_X1    g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1215), .A2(new_n1219), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1213), .B1(new_n1227), .B2(new_n792), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1211), .A2(new_n779), .B1(new_n1212), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n986), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1105), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1094), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1211), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1229), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT125), .ZN(G381));
  NAND2_X1  g1035(.A1(G378), .A2(KEYINPUT126), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT126), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1122), .A2(new_n1145), .A3(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n1209), .A3(new_n1177), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1241));
  OR4_X1    g1041(.A1(G387), .A2(new_n1240), .A3(new_n1241), .A4(G381), .ZN(G407));
  OAI211_X1 g1042(.A(G407), .B(G213), .C1(G343), .C2(new_n1240), .ZN(G409));
  XOR2_X1   g1043(.A(G393), .B(G396), .Z(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n999), .A2(new_n1024), .A3(G390), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G390), .B1(new_n999), .B2(new_n1024), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1245), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1248), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1177), .A2(G378), .A3(new_n1209), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1174), .A2(new_n1230), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1209), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1236), .A2(new_n1256), .A3(new_n1238), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n716), .A2(G343), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1094), .A4(new_n1103), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT127), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1233), .A2(KEYINPUT60), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1105), .A2(new_n739), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(G384), .A3(new_n1229), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G384), .B1(new_n1271), .B2(new_n1229), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G2897), .B(new_n1259), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1274), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1259), .A2(G2897), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1272), .A3(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1261), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1259), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1282), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1253), .A2(new_n1280), .A3(new_n1284), .A4(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1285), .A2(new_n1288), .A3(new_n1282), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1285), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1288), .B1(new_n1285), .B2(new_n1282), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1289), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1287), .B1(new_n1294), .B2(new_n1253), .ZN(G405));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1239), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1254), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1282), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1283), .A3(new_n1254), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(new_n1252), .ZN(G402));
endmodule


