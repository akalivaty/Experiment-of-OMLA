//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT66), .B(G238), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(new_n202), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G77), .A2(G244), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G50), .B2(G226), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G97), .A2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(G87), .A2(G250), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT65), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n230), .A2(G1), .A3(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n206), .A2(new_n207), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n214), .B(new_n227), .C1(new_n235), .C2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G226), .B(G232), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT68), .ZN(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n207), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n229), .A2(new_n231), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n260), .B1(new_n255), .B2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G50), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT74), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT72), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n201), .A2(KEYINPUT72), .A3(KEYINPUT8), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT73), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n234), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT73), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n267), .A2(new_n268), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n263), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n279), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n271), .A2(new_n274), .ZN(new_n282));
  INV_X1    g0082(.A(new_n268), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT8), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n264), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(KEYINPUT74), .B(new_n281), .C1(new_n282), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n208), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n280), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(KEYINPUT75), .A3(new_n260), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT75), .B1(new_n290), .B2(new_n260), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n258), .B(new_n262), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n290), .A2(new_n260), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT75), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n291), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(KEYINPUT9), .A3(new_n258), .A4(new_n262), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G77), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n229), .A2(new_n231), .B1(G33), .B2(G41), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G222), .A2(G1698), .ZN(new_n309));
  XOR2_X1   g0109(.A(KEYINPUT71), .B(G223), .Z(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n307), .B(new_n308), .C1(new_n311), .C2(new_n305), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n255), .A2(G274), .ZN(new_n313));
  INV_X1    g0113(.A(G41), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT69), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G41), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G45), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(G1), .B(G13), .C1(new_n269), .C2(new_n314), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT70), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n322), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G226), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n312), .B(new_n321), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n296), .A2(new_n301), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT10), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT76), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n294), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n336), .B1(new_n294), .B2(new_n338), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n330), .A2(G179), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n282), .A2(new_n306), .B1(new_n207), .B2(new_n277), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n234), .A2(G68), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n260), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT11), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n261), .A2(G68), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n257), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT12), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n256), .B2(G68), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT80), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n325), .A2(G238), .A3(new_n327), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  MUX2_X1   g0156(.A(G226), .B(G232), .S(G1698), .Z(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT3), .B(G33), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n357), .A2(new_n358), .B1(G33), .B2(G97), .ZN(new_n359));
  INV_X1    g0159(.A(new_n308), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n321), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n354), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n359), .A2(new_n360), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .A3(new_n321), .A4(new_n355), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n364), .A3(G200), .ZN(new_n365));
  OAI211_X1 g0165(.A(KEYINPUT79), .B(KEYINPUT13), .C1(new_n356), .C2(new_n361), .ZN(new_n366));
  NAND2_X1  g0166(.A1(KEYINPUT79), .A2(KEYINPUT13), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n363), .A2(new_n321), .A3(new_n355), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(G190), .A3(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n346), .A2(new_n353), .A3(new_n365), .A4(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n305), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(G232), .A2(G1698), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n215), .B2(G1698), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n308), .B(new_n373), .C1(new_n375), .C2(new_n305), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n325), .A2(G244), .A3(new_n327), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n321), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT77), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT77), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .A4(new_n321), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n371), .B1(new_n382), .B2(new_n332), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n256), .A2(G77), .ZN(new_n384));
  INV_X1    g0184(.A(new_n260), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n264), .A2(new_n285), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n387));
  OR2_X1    g0187(.A1(KEYINPUT15), .A2(G87), .ZN(new_n388));
  NAND2_X1  g0188(.A1(KEYINPUT15), .A2(G87), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n270), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n385), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n384), .B(new_n391), .C1(G77), .C2(new_n261), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n382), .B2(G200), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n379), .A2(new_n381), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT78), .A3(G190), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n383), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n362), .A2(new_n364), .A3(G169), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT14), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n366), .A2(G179), .A3(new_n368), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n362), .A2(new_n364), .A3(new_n401), .A4(G169), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n346), .A2(new_n353), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n382), .A2(new_n337), .ZN(new_n406));
  INV_X1    g0206(.A(G179), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n392), .B1(new_n395), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND4_X1   g0209(.A1(new_n370), .A2(new_n397), .A3(new_n405), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n358), .A2(new_n412), .A3(G20), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT7), .B1(new_n305), .B2(new_n234), .ZN(new_n414));
  OAI21_X1  g0214(.A(G68), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G58), .A2(G68), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n203), .A2(new_n205), .A3(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(KEYINPUT16), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n412), .B1(new_n358), .B2(G20), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n305), .A2(KEYINPUT7), .A3(new_n234), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n202), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n417), .A2(G20), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n276), .A2(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n420), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n419), .A2(new_n427), .A3(new_n260), .ZN(new_n428));
  INV_X1    g0228(.A(new_n287), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n261), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n287), .A2(new_n257), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT81), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n428), .A2(KEYINPUT81), .A3(new_n430), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OR2_X1    g0236(.A1(G223), .A2(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n329), .A2(G1698), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n358), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G87), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n308), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n322), .A2(G232), .A3(new_n323), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n321), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n407), .B2(new_n444), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n411), .B1(new_n436), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n444), .A2(new_n407), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(G169), .B2(new_n444), .ZN(new_n449));
  AOI211_X1 g0249(.A(KEYINPUT18), .B(new_n449), .C1(new_n434), .C2(new_n435), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n320), .B1(new_n441), .B2(new_n308), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n451), .A2(new_n332), .A3(new_n443), .ZN(new_n452));
  AOI21_X1  g0252(.A(G200), .B1(new_n451), .B2(new_n443), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT82), .ZN(new_n454));
  OR3_X1    g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n451), .A2(new_n454), .A3(new_n332), .A4(new_n443), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT17), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n428), .A2(new_n457), .A3(new_n430), .A4(new_n431), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n447), .A2(new_n450), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n335), .A2(new_n342), .A3(new_n410), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G200), .ZN(new_n467));
  AND2_X1   g0267(.A1(G264), .A2(G1698), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT86), .B1(new_n358), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n302), .A2(new_n304), .A3(new_n468), .A4(KEYINPUT86), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n302), .A2(new_n304), .A3(G257), .ZN(new_n473));
  INV_X1    g0273(.A(G1698), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n473), .A2(new_n474), .B1(G303), .B2(new_n305), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n360), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT5), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n255), .B(G45), .C1(new_n478), .C2(G41), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n315), .A2(new_n317), .A3(new_n478), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G270), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT69), .B(G41), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n479), .B1(new_n484), .B2(new_n478), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G274), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT87), .B1(new_n476), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n302), .A2(new_n304), .A3(new_n468), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n358), .A2(G257), .A3(new_n474), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n305), .A2(G303), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n470), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n308), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n482), .A2(G270), .B1(new_n485), .B2(G274), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT87), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n467), .B1(new_n488), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n255), .A2(G33), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n385), .A2(new_n256), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G116), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n256), .A2(G116), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G116), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  INV_X1    g0308(.A(G97), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n234), .C1(G33), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n260), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT20), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n507), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n503), .A2(new_n505), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT88), .B1(new_n499), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n497), .B1(new_n495), .B2(new_n496), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  OAI21_X1  g0321(.A(G200), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT88), .ZN(new_n523));
  INV_X1    g0323(.A(new_n516), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n517), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n302), .A2(new_n304), .A3(new_n234), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n358), .A2(new_n529), .A3(new_n234), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n270), .A2(G116), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n234), .A2(G107), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n533), .B(KEYINPUT23), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT24), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n531), .A2(KEYINPUT24), .A3(new_n532), .A4(new_n534), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n260), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n385), .A2(G107), .A3(new_n256), .A4(new_n500), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT25), .B1(new_n256), .B2(G107), .ZN(new_n541));
  OR3_X1    g0341(.A1(new_n256), .A2(KEYINPUT25), .A3(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT89), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n540), .A2(KEYINPUT89), .A3(new_n541), .A4(new_n542), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n302), .A2(new_n304), .A3(G250), .A4(new_n474), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n302), .A2(new_n304), .A3(G257), .A4(G1698), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G294), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n308), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n482), .A2(G264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n486), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n337), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n555), .A2(G179), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n548), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G169), .B(new_n516), .C1(new_n518), .C2(new_n519), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n476), .A2(new_n487), .A3(new_n407), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n516), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n488), .A2(new_n498), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(KEYINPUT21), .A3(G169), .A4(new_n516), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n558), .A2(new_n561), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n509), .A2(new_n372), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n372), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n573));
  OAI21_X1  g0373(.A(G107), .B1(new_n413), .B2(new_n414), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n385), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n501), .A2(new_n509), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n256), .A2(G97), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n302), .A2(new_n304), .A3(G244), .A4(new_n474), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n358), .A2(KEYINPUT4), .A3(G244), .A4(new_n474), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n358), .A2(G250), .A3(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n508), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n308), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n482), .A2(G257), .B1(new_n485), .B2(G274), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G190), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n584), .A2(KEYINPUT83), .A3(new_n308), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT83), .B1(new_n584), .B2(new_n308), .ZN(new_n590));
  INV_X1    g0390(.A(new_n586), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n578), .B(new_n588), .C1(new_n592), .C2(new_n467), .ZN(new_n593));
  INV_X1    g0393(.A(new_n590), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n584), .A2(KEYINPUT83), .A3(new_n308), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n407), .A3(new_n586), .A4(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n576), .ZN(new_n597));
  INV_X1    g0397(.A(new_n577), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n573), .A2(new_n574), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n385), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n585), .A2(new_n586), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n337), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n596), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n555), .A2(new_n467), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n553), .A2(new_n554), .A3(new_n332), .A4(new_n486), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(KEYINPUT90), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT90), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n555), .A2(new_n607), .A3(new_n467), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n606), .A2(new_n547), .A3(new_n539), .A4(new_n608), .ZN(new_n609));
  OR2_X1    g0409(.A1(G238), .A2(G1698), .ZN(new_n610));
  INV_X1    g0410(.A(G244), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G1698), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n302), .A2(new_n610), .A3(new_n304), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G33), .A2(G116), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n308), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n255), .A2(G45), .A3(G274), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n322), .B(G250), .C1(G1), .C2(new_n319), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  AND2_X1   g0420(.A1(KEYINPUT84), .A2(G87), .ZN(new_n621));
  NOR2_X1   g0421(.A1(KEYINPUT84), .A2(G87), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n569), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n234), .B1(new_n269), .B2(new_n509), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(KEYINPUT19), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n358), .A2(new_n234), .A3(G68), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT19), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n272), .B2(new_n509), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n388), .A2(new_n389), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n629), .A2(new_n260), .B1(new_n257), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n502), .A2(G87), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n616), .A2(G190), .A3(new_n617), .A4(new_n618), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n620), .A2(new_n631), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n629), .A2(new_n260), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n388), .A2(KEYINPUT85), .A3(new_n389), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(new_n385), .A3(new_n256), .A4(new_n500), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n630), .A2(new_n257), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n619), .A2(new_n337), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n616), .A2(new_n407), .A3(new_n617), .A4(new_n618), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n593), .A2(new_n603), .A3(new_n609), .A4(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n526), .A2(new_n566), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n466), .A2(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n342), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n432), .A2(new_n446), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(new_n411), .ZN(new_n652));
  INV_X1    g0452(.A(new_n405), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT92), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n406), .A2(new_n408), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(new_n406), .B2(new_n408), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n653), .B1(new_n657), .B2(new_n370), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n652), .B1(new_n658), .B2(new_n463), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n650), .B1(new_n659), .B2(new_n335), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n563), .A2(new_n558), .A3(new_n561), .A4(new_n565), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n645), .B1(new_n661), .B2(new_n647), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n634), .A2(new_n645), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n603), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n603), .B2(new_n663), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT91), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT91), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n668), .B(new_n664), .C1(new_n603), .C2(new_n663), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n660), .B1(new_n465), .B2(new_n671), .ZN(G369));
  INV_X1    g0472(.A(G13), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G20), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OR3_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .A3(G1), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT27), .B1(new_n675), .B2(G1), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n558), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n548), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n609), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n558), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n561), .A2(new_n565), .A3(new_n563), .ZN(new_n685));
  INV_X1    g0485(.A(new_n680), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n681), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT93), .Z(new_n689));
  NOR2_X1   g0489(.A1(new_n526), .A2(new_n685), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n524), .A2(new_n686), .ZN(new_n691));
  MUX2_X1   g0491(.A(new_n690), .B(new_n685), .S(new_n691), .Z(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(G330), .A3(new_n684), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n693), .ZN(G399));
  NOR2_X1   g0494(.A1(new_n621), .A2(new_n622), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n506), .A3(new_n569), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT94), .ZN(new_n698));
  INV_X1    g0498(.A(new_n212), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n484), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(G1), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n236), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n686), .B1(new_n662), .B2(new_n670), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n666), .ZN(new_n709));
  OAI221_X1 g0509(.A(new_n645), .B1(new_n709), .B2(new_n665), .C1(new_n661), .C2(new_n647), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n686), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n520), .A2(new_n592), .A3(G179), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n555), .A3(new_n619), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n553), .A2(new_n554), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n619), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n562), .A2(new_n587), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT30), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n686), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT95), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n722), .A3(KEYINPUT31), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n648), .B2(new_n686), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n721), .B(new_n723), .C1(new_n725), .C2(new_n719), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G330), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n712), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n705), .B1(new_n730), .B2(G1), .ZN(G364));
  AOI21_X1  g0531(.A(new_n255), .B1(new_n674), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n700), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n699), .A2(new_n358), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n250), .B2(G45), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G45), .B2(new_n703), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n358), .A2(G355), .A3(new_n212), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n739), .B(new_n740), .C1(G116), .C2(new_n212), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n233), .B1(G20), .B2(new_n337), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT97), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n750), .A2(new_n234), .A3(G190), .ZN(new_n751));
  NOR4_X1   g0551(.A1(new_n234), .A2(new_n407), .A3(new_n467), .A4(G190), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT33), .B(G317), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n751), .A2(G329), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n234), .A2(G190), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G179), .A3(new_n467), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G311), .ZN(new_n758));
  INV_X1    g0558(.A(G303), .ZN(new_n759));
  NAND2_X1  g0559(.A1(G20), .A2(G190), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n760), .A2(new_n467), .A3(G179), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n754), .B(new_n758), .C1(new_n759), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n234), .A2(new_n407), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(G326), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n760), .A2(new_n407), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n763), .A2(new_n358), .A3(new_n767), .A4(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n755), .A2(new_n407), .A3(G200), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT98), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT98), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  OAI21_X1  g0578(.A(G20), .B1(new_n750), .B2(new_n332), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n772), .B1(new_n773), .B2(new_n777), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT99), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  INV_X1    g0584(.A(new_n752), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n358), .B1(new_n696), .B2(new_n762), .C1(new_n785), .C2(new_n202), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n780), .A2(new_n509), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n751), .A2(G159), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n786), .B(new_n787), .C1(KEYINPUT32), .C2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n207), .B2(new_n765), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n777), .A2(new_n372), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n756), .A2(KEYINPUT96), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n756), .A2(KEYINPUT96), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n791), .B1(G77), .B2(new_n795), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n796), .B1(KEYINPUT32), .B2(new_n788), .C1(new_n201), .C2(new_n769), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n783), .A2(new_n784), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n735), .B(new_n747), .C1(new_n799), .C2(new_n742), .ZN(new_n800));
  INV_X1    g0600(.A(new_n745), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n692), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT101), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n734), .B1(new_n692), .B2(G330), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G330), .B2(new_n692), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  AOI22_X1  g0608(.A1(new_n751), .A2(G311), .B1(G107), .B2(new_n761), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n506), .B2(new_n794), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n787), .B1(G283), .B2(new_n752), .ZN(new_n811));
  INV_X1    g0611(.A(new_n777), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G87), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n358), .B1(new_n766), .B2(G303), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n810), .B(new_n815), .C1(G294), .C2(new_n768), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n812), .A2(G68), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n752), .A2(G150), .B1(G143), .B2(new_n768), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n766), .A2(G137), .ZN(new_n819));
  INV_X1    g0619(.A(G159), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n818), .B(new_n819), .C1(new_n794), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n751), .A2(G132), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n305), .B1(G50), .B2(new_n761), .ZN(new_n824));
  AND4_X1   g0624(.A1(new_n817), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n779), .A2(G58), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n816), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n742), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n734), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n742), .A2(new_n743), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT102), .Z(new_n831));
  AOI21_X1  g0631(.A(new_n829), .B1(new_n306), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT103), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n393), .A2(new_n680), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n655), .B2(new_n656), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n397), .A2(new_n409), .A3(new_n834), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n833), .B1(new_n744), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT104), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n727), .A2(new_n728), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n838), .B(KEYINPUT105), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n706), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n838), .B(new_n686), .C1(new_n662), .C2(new_n670), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n841), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n735), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n840), .A2(new_n847), .ZN(G384));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  INV_X1    g0649(.A(new_n678), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n432), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n447), .A2(new_n450), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n458), .A2(new_n462), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n460), .B2(new_n461), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n436), .B2(new_n446), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n436), .A2(new_n850), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(new_n651), .A3(new_n851), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n857), .A2(new_n858), .B1(new_n860), .B2(KEYINPUT37), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n849), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n857), .A2(new_n858), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(KEYINPUT38), .C1(new_n464), .C2(new_n851), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n653), .A2(new_n680), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n404), .A2(new_n680), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n405), .A2(new_n370), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n409), .A2(new_n680), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n872), .B1(new_n844), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n651), .B(KEYINPUT18), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n678), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n859), .A2(new_n651), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n678), .B1(new_n434), .B2(new_n435), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n863), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n881), .B1(new_n877), .B2(new_n463), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT107), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n866), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n436), .A2(new_n446), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT18), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n436), .A2(new_n411), .A3(new_n446), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n853), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n851), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n891), .A2(new_n892), .B1(new_n864), .B2(new_n863), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(KEYINPUT107), .A3(KEYINPUT38), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT39), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n866), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n405), .A2(new_n680), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n879), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n660), .B1(new_n712), .B2(new_n465), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  AND4_X1   g0701(.A1(new_n603), .A2(new_n593), .A3(new_n609), .A4(new_n646), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n517), .A2(new_n521), .A3(new_n525), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n661), .A2(new_n902), .A3(new_n903), .A4(new_n686), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT31), .ZN(new_n905));
  INV_X1    g0705(.A(new_n719), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n465), .B1(new_n720), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(G330), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n871), .A2(new_n838), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n907), .B2(new_n720), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n867), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n858), .A2(new_n859), .A3(new_n651), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .B1(new_n858), .B2(new_n857), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n858), .B1(new_n853), .B2(new_n652), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n849), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n918), .A2(KEYINPUT107), .B1(new_n893), .B2(KEYINPUT38), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n866), .A2(new_n886), .ZN(new_n920));
  OAI211_X1 g0720(.A(KEYINPUT40), .B(new_n911), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(new_n921), .A3(G330), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT40), .B1(new_n867), .B2(new_n911), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n870), .A2(new_n868), .B1(new_n836), .B2(new_n837), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n719), .B1(new_n904), .B2(KEYINPUT31), .ZN(new_n925));
  INV_X1    g0725(.A(new_n720), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n887), .B2(new_n894), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n923), .B1(KEYINPUT40), .B2(new_n928), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n909), .A2(new_n922), .B1(new_n929), .B2(new_n908), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n901), .B(new_n930), .Z(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n255), .B2(new_n674), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n236), .A2(G77), .A3(new_n416), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(G50), .B2(new_n202), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(G1), .A3(new_n673), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n506), .B1(new_n572), .B2(KEYINPUT35), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(new_n235), .C1(KEYINPUT35), .C2(new_n572), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT106), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n935), .A3(new_n939), .ZN(G367));
  AOI22_X1  g0740(.A1(new_n766), .A2(G311), .B1(G303), .B2(new_n768), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT46), .B1(new_n761), .B2(G116), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G294), .B2(new_n752), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT111), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(KEYINPUT111), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n941), .B1(new_n947), .B2(KEYINPUT112), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n947), .A2(KEYINPUT112), .B1(G317), .B2(new_n751), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(new_n305), .C1(new_n509), .C2(new_n777), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n948), .B(new_n950), .C1(G283), .C2(new_n795), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n372), .B2(new_n780), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n777), .A2(new_n306), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n780), .A2(new_n202), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n953), .B(new_n954), .C1(G137), .C2(new_n751), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n794), .A2(new_n207), .B1(new_n278), .B2(new_n769), .ZN(new_n956));
  INV_X1    g0756(.A(G143), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n762), .A2(new_n201), .B1(new_n765), .B2(new_n957), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n956), .A2(new_n305), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n955), .B(new_n959), .C1(new_n820), .C2(new_n785), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n952), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n742), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n631), .A2(new_n632), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n680), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n646), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(KEYINPUT108), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n645), .C2(new_n965), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(new_n801), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n746), .B1(new_n212), .B2(new_n630), .C1(new_n245), .C2(new_n737), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n963), .A2(new_n734), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT113), .Z(new_n973));
  OAI211_X1 g0773(.A(new_n593), .B(new_n603), .C1(new_n578), .C2(new_n686), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n603), .A2(new_n686), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n689), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT110), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n977), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n689), .A2(new_n976), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT45), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n693), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n687), .B1(new_n692), .B2(G330), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n684), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n730), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n729), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n700), .B(KEYINPUT41), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n732), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n684), .A2(new_n687), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n974), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT42), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n603), .B1(new_n974), .B2(new_n558), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n686), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n994), .A2(new_n996), .B1(KEYINPUT43), .B2(new_n969), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n976), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n693), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n999), .B(new_n1001), .Z(new_n1002));
  AOI21_X1  g0802(.A(new_n973), .B1(new_n991), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(G387));
  NAND2_X1  g0804(.A1(new_n986), .A2(new_n733), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n752), .A2(G311), .B1(G317), .B2(new_n768), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n770), .B2(new_n765), .C1(new_n794), .C2(new_n759), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT48), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n773), .B2(new_n780), .C1(new_n778), .C2(new_n762), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n812), .A2(G116), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n751), .A2(G326), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1010), .A2(new_n305), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n779), .A2(new_n639), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n761), .A2(G77), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n766), .A2(G159), .ZN(new_n1016));
  AND4_X1   g0816(.A1(new_n358), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n812), .A2(G97), .B1(new_n751), .B2(G150), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n768), .A2(G50), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n429), .A2(new_n752), .B1(new_n757), .B2(G68), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n828), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(G68), .A2(G77), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n386), .A2(new_n207), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT50), .Z(new_n1025));
  NAND4_X1  g0825(.A1(new_n698), .A2(new_n319), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n737), .B1(new_n242), .B2(G45), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n698), .A2(new_n699), .A3(new_n305), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(G107), .B2(new_n212), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n735), .B(new_n1022), .C1(new_n746), .C2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n684), .B2(new_n801), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n700), .B1(new_n730), .B2(new_n986), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1005), .B(new_n1032), .C1(new_n987), .C2(new_n1033), .ZN(G393));
  NAND2_X1  g0834(.A1(new_n984), .A2(new_n987), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n983), .B(new_n693), .Z(new_n1036));
  OAI211_X1 g0836(.A(new_n700), .B(new_n1035), .C1(new_n1036), .C2(new_n987), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n733), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n735), .B1(new_n1000), .B2(new_n745), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n756), .A2(new_n778), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1040), .B(new_n791), .C1(G322), .C2(new_n751), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n761), .A2(G283), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n766), .A2(G317), .B1(G311), .B2(new_n768), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  OAI21_X1  g0844(.A(new_n305), .B1(new_n780), .B2(new_n506), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G303), .B2(new_n752), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n795), .A2(new_n386), .B1(G50), .B2(new_n752), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1049), .A2(KEYINPUT114), .B1(G68), .B2(new_n761), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n305), .B1(new_n779), .B2(G77), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n751), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n813), .B1(new_n957), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n766), .A2(G150), .B1(G159), .B2(new_n768), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1050), .A2(new_n1051), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1049), .A2(KEYINPUT114), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1047), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n742), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n746), .B1(new_n509), .B2(new_n212), .C1(new_n253), .C2(new_n737), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1039), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1037), .A2(new_n1038), .A3(new_n1062), .ZN(G390));
  OAI21_X1  g0863(.A(G330), .B1(new_n925), .B2(new_n926), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n872), .B1(new_n1064), .B2(new_n842), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n726), .A2(G330), .A3(new_n924), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n710), .A2(new_n686), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n873), .B1(new_n1067), .B2(new_n838), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(G330), .B(new_n924), .C1(new_n925), .C2(new_n926), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n726), .A2(G330), .A3(new_n838), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n872), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n844), .A2(new_n874), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1069), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n900), .B1(G330), .B2(new_n908), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT116), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1075), .A2(KEYINPUT116), .A3(new_n1076), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n898), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n919), .B2(new_n920), .C1(new_n1068), .C2(new_n872), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT115), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n1082), .C1(new_n1074), .C2(new_n872), .ZN(new_n1085));
  OAI21_X1  g0885(.A(KEYINPUT115), .B1(new_n875), .B2(new_n898), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n897), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n1070), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1066), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1083), .B(new_n1090), .C1(new_n897), .C2(new_n1087), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1081), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1079), .A2(new_n1089), .A3(new_n1091), .A4(new_n1080), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n700), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n743), .B1(new_n895), .B2(new_n896), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n831), .A2(new_n287), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n761), .A2(G150), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1098), .A2(KEYINPUT53), .B1(G132), .B2(new_n768), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(KEYINPUT53), .B2(new_n1098), .C1(new_n780), .C2(new_n820), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT54), .B(G143), .Z(new_n1101));
  AOI22_X1  g0901(.A1(new_n795), .A2(new_n1101), .B1(G137), .B2(new_n752), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT117), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n751), .A2(G125), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n812), .A2(G50), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1103), .A2(new_n358), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1100), .B(new_n1106), .C1(G128), .C2(new_n766), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n779), .A2(G77), .B1(G116), .B2(new_n768), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT118), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n766), .A2(G283), .B1(G87), .B2(new_n761), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n509), .C2(new_n794), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n817), .B1(new_n372), .B2(new_n785), .C1(new_n778), .C2(new_n1052), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1111), .A2(new_n358), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n742), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1096), .A2(new_n734), .A3(new_n1097), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT119), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1092), .A2(new_n733), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1095), .A2(new_n1119), .ZN(G378));
  INV_X1    g0920(.A(new_n899), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n342), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n294), .A2(new_n850), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1127), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n335), .B2(new_n342), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1123), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n335), .A2(new_n342), .A3(new_n1129), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n1122), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n929), .B2(G330), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1135), .A2(new_n914), .A3(new_n921), .A4(G330), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1121), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1135), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n922), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n899), .A3(new_n1137), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1079), .A2(new_n1080), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n909), .B(new_n660), .C1(new_n465), .C2(new_n712), .ZN(new_n1145));
  OAI211_X1 g0945(.A(KEYINPUT57), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n700), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT122), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT123), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1093), .A2(new_n1076), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1141), .A2(new_n899), .A3(new_n1137), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n899), .B1(new_n1141), .B2(new_n1137), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT122), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT123), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n1157), .A3(new_n1150), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1152), .A2(new_n1153), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1147), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1152), .A2(new_n733), .A3(new_n1158), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n765), .A2(new_n506), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n954), .B1(G283), .B2(new_n751), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n639), .A2(new_n757), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n812), .A2(G58), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1164), .B(new_n1168), .C1(G107), .C2(new_n768), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n484), .A2(new_n358), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n752), .A2(G97), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1169), .A2(new_n1015), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT58), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n757), .A2(G137), .B1(new_n768), .B2(G128), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n766), .A2(G125), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n752), .A2(G132), .B1(new_n1101), .B2(new_n761), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G150), .B2(new_n779), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT59), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(G33), .A2(G41), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT120), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n777), .A2(new_n820), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G124), .C2(new_n751), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1170), .A2(G50), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1179), .A2(new_n1183), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n828), .B1(new_n1173), .B2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT121), .Z(new_n1187));
  AOI21_X1  g0987(.A(new_n735), .B1(new_n830), .B2(new_n207), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n744), .C2(new_n1135), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1163), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1162), .A2(new_n1191), .ZN(G375));
  NAND2_X1  g0992(.A1(new_n752), .A2(new_n1101), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n780), .B2(new_n207), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n305), .B(new_n1194), .C1(G132), .C2(new_n766), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n757), .A2(G150), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n751), .A2(G128), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G137), .A2(new_n768), .B1(new_n761), .B2(G159), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1167), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1014), .B1(new_n773), .B2(new_n769), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT124), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n785), .A2(new_n506), .B1(new_n509), .B2(new_n762), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n751), .B2(G303), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n305), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n953), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n372), .B2(new_n794), .C1(new_n778), .C2(new_n765), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1200), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n742), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n734), .B(new_n1209), .C1(new_n871), .C2(new_n744), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n202), .B2(new_n831), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1075), .B2(new_n733), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1079), .A2(new_n1080), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1212), .B1(new_n1215), .B2(new_n990), .ZN(G381));
  OR3_X1    g1016(.A1(new_n1161), .A2(G378), .A3(new_n1190), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(G396), .A2(G393), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1218), .A2(new_n1003), .A3(new_n1219), .A4(new_n1220), .ZN(G407));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G343), .C2(new_n1217), .ZN(G409));
  OAI21_X1  g1022(.A(G378), .B1(new_n1161), .B2(new_n1190), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1143), .A2(new_n733), .ZN(new_n1224));
  AND4_X1   g1024(.A1(new_n1119), .A2(new_n1095), .A3(new_n1189), .A4(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1152), .A2(new_n1158), .A3(new_n989), .A4(new_n1153), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1225), .A2(new_n1226), .B1(G213), .B2(new_n679), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1213), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n700), .B(new_n1229), .C1(new_n1214), .C2(new_n1228), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(G384), .A3(new_n1212), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G384), .B1(new_n1230), .B2(new_n1212), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1223), .A2(new_n1227), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT62), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1223), .A2(new_n1227), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n679), .A2(G213), .A3(G2897), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1232), .A2(new_n1233), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1230), .A2(new_n1212), .ZN(new_n1241));
  INV_X1    g1041(.A(G384), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1238), .B1(new_n1243), .B2(new_n1231), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1237), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1223), .A2(new_n1248), .A3(new_n1227), .A4(new_n1234), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1236), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(G396), .A2(G393), .ZN(new_n1251));
  OR3_X1    g1051(.A1(new_n1003), .A2(new_n1220), .A3(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1003), .A2(KEYINPUT126), .B1(new_n1251), .B2(new_n1220), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G390), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(G390), .A3(new_n1253), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1250), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT125), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1237), .A2(new_n1261), .A3(new_n1245), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1237), .B2(new_n1245), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1247), .B(new_n1258), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1235), .B(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1260), .B1(new_n1264), .B2(new_n1266), .ZN(G405));
  NAND2_X1  g1067(.A1(new_n1217), .A2(new_n1223), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT127), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1234), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1234), .A2(new_n1269), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1217), .A2(new_n1223), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1258), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1259), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(G402));
endmodule


