

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(n710), .A2(n971), .ZN(n709) );
  XNOR2_X1 U555 ( .A(KEYINPUT75), .B(n616), .ZN(n963) );
  XNOR2_X1 U556 ( .A(n537), .B(KEYINPUT89), .ZN(n697) );
  XOR2_X2 U557 ( .A(G2104), .B(KEYINPUT64), .Z(n522) );
  AND2_X2 U558 ( .A1(n907), .A2(G102), .ZN(n528) );
  XNOR2_X1 U559 ( .A(n722), .B(KEYINPUT100), .ZN(n725) );
  OR2_X2 U560 ( .A1(n810), .A2(n812), .ZN(n749) );
  NOR2_X1 U561 ( .A1(G651), .A2(n660), .ZN(n664) );
  INV_X1 U562 ( .A(KEYINPUT108), .ZN(n782) );
  XNOR2_X1 U563 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X2 U564 ( .A(n527), .B(n526), .ZN(n907) );
  AND2_X1 U565 ( .A1(n533), .A2(n532), .ZN(n520) );
  XOR2_X1 U566 ( .A(KEYINPUT74), .B(n614), .Z(n521) );
  AND2_X1 U567 ( .A1(n707), .A2(n706), .ZN(n523) );
  OR2_X1 U568 ( .A1(n840), .A2(n839), .ZN(n524) );
  AND2_X1 U569 ( .A1(n841), .A2(n524), .ZN(n525) );
  AND2_X1 U570 ( .A1(n708), .A2(n523), .ZN(n710) );
  AND2_X1 U571 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U572 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n738) );
  XNOR2_X1 U573 ( .A(n739), .B(n738), .ZN(n740) );
  INV_X1 U574 ( .A(n697), .ZN(n699) );
  NAND2_X1 U575 ( .A1(n699), .A2(n698), .ZN(n810) );
  INV_X1 U576 ( .A(KEYINPUT68), .ZN(n529) );
  XNOR2_X1 U577 ( .A(n529), .B(KEYINPUT17), .ZN(n530) );
  INV_X1 U578 ( .A(KEYINPUT65), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n534), .A2(n520), .ZN(n535) );
  OR2_X2 U580 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U581 ( .A(n543), .B(KEYINPUT66), .ZN(n544) );
  BUF_X1 U582 ( .A(n697), .Z(G164) );
  NOR2_X2 U583 ( .A1(n522), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U584 ( .A(n528), .B(KEYINPUT88), .ZN(n536) );
  AND2_X1 U585 ( .A1(n522), .A2(G2105), .ZN(n904) );
  NAND2_X1 U586 ( .A1(G126), .A2(n904), .ZN(n534) );
  AND2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n903) );
  NAND2_X1 U588 ( .A1(G114), .A2(n903), .ZN(n533) );
  NOR2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  XNOR2_X2 U590 ( .A(n531), .B(n530), .ZN(n567) );
  NAND2_X1 U591 ( .A1(G138), .A2(n567), .ZN(n532) );
  NAND2_X1 U592 ( .A1(G137), .A2(n567), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n903), .A2(G113), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U595 ( .A(n540), .B(KEYINPUT69), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G125), .A2(n904), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G101), .A2(n907), .ZN(n545) );
  XOR2_X1 U599 ( .A(KEYINPUT23), .B(KEYINPUT67), .Z(n543) );
  NOR2_X2 U600 ( .A1(n547), .A2(n546), .ZN(G160) );
  INV_X1 U601 ( .A(G651), .ZN(n551) );
  NOR2_X1 U602 ( .A1(G543), .A2(n551), .ZN(n548) );
  XOR2_X1 U603 ( .A(KEYINPUT1), .B(n548), .Z(n663) );
  NAND2_X1 U604 ( .A1(G60), .A2(n663), .ZN(n550) );
  XOR2_X1 U605 ( .A(KEYINPUT0), .B(G543), .Z(n660) );
  NAND2_X1 U606 ( .A1(G47), .A2(n664), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n555) );
  NOR2_X2 U608 ( .A1(n660), .A2(n551), .ZN(n667) );
  NAND2_X1 U609 ( .A1(G72), .A2(n667), .ZN(n553) );
  NOR2_X2 U610 ( .A1(G651), .A2(G543), .ZN(n672) );
  NAND2_X1 U611 ( .A1(G85), .A2(n672), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  OR2_X1 U613 ( .A1(n555), .A2(n554), .ZN(G290) );
  XNOR2_X1 U614 ( .A(G2443), .B(G2435), .ZN(n565) );
  XOR2_X1 U615 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n557) );
  XNOR2_X1 U616 ( .A(G2454), .B(G2430), .ZN(n556) );
  XNOR2_X1 U617 ( .A(n557), .B(n556), .ZN(n561) );
  XOR2_X1 U618 ( .A(G2427), .B(G2438), .Z(n559) );
  XNOR2_X1 U619 ( .A(G1348), .B(G1341), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U621 ( .A(n561), .B(n560), .Z(n563) );
  XNOR2_X1 U622 ( .A(G2451), .B(G2446), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U624 ( .A(n565), .B(n564), .ZN(n566) );
  AND2_X1 U625 ( .A1(n566), .A2(G14), .ZN(G401) );
  AND2_X1 U626 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U627 ( .A1(G111), .A2(n903), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G135), .A2(n567), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U630 ( .A1(n904), .A2(G123), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT18), .B(n570), .Z(n571) );
  NOR2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n907), .A2(G99), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n939) );
  XNOR2_X1 U635 ( .A(G2096), .B(n939), .ZN(n575) );
  OR2_X1 U636 ( .A1(G2100), .A2(n575), .ZN(G156) );
  INV_X1 U637 ( .A(G57), .ZN(G237) );
  INV_X1 U638 ( .A(G82), .ZN(G220) );
  NAND2_X1 U639 ( .A1(G64), .A2(n663), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT70), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G52), .A2(n664), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT71), .B(n577), .Z(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G77), .A2(n667), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G90), .A2(n672), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(KEYINPUT9), .B(n582), .Z(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(G171) );
  INV_X1 U649 ( .A(G171), .ZN(G301) );
  NAND2_X1 U650 ( .A1(G75), .A2(n667), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G88), .A2(n672), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(KEYINPUT87), .B(n587), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G62), .A2(n663), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G50), .A2(n664), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U657 ( .A(KEYINPUT86), .B(n590), .Z(n591) );
  NAND2_X1 U658 ( .A1(n592), .A2(n591), .ZN(G303) );
  NAND2_X1 U659 ( .A1(n672), .A2(G89), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n593), .B(KEYINPUT4), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G76), .A2(n667), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U663 ( .A(n596), .B(KEYINPUT5), .ZN(n602) );
  NAND2_X1 U664 ( .A1(n663), .A2(G63), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT78), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G51), .A2(n664), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U668 ( .A(KEYINPUT6), .B(n600), .Z(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n603), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U671 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U672 ( .A1(G7), .A2(G661), .ZN(n604) );
  XOR2_X1 U673 ( .A(n604), .B(KEYINPUT10), .Z(n854) );
  NAND2_X1 U674 ( .A1(n854), .A2(G567), .ZN(n605) );
  XOR2_X1 U675 ( .A(KEYINPUT11), .B(n605), .Z(G234) );
  NAND2_X1 U676 ( .A1(n663), .A2(G56), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT14), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G43), .A2(n664), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n615) );
  NAND2_X1 U680 ( .A1(G68), .A2(n667), .ZN(n612) );
  XOR2_X1 U681 ( .A(KEYINPUT12), .B(KEYINPUT73), .Z(n610) );
  NAND2_X1 U682 ( .A1(G81), .A2(n672), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n610), .B(n609), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n613), .B(KEYINPUT13), .ZN(n614) );
  NOR2_X1 U686 ( .A1(n615), .A2(n521), .ZN(n616) );
  INV_X1 U687 ( .A(G860), .ZN(n638) );
  OR2_X1 U688 ( .A1(n963), .A2(n638), .ZN(G153) );
  NAND2_X1 U689 ( .A1(G868), .A2(G301), .ZN(n627) );
  NAND2_X1 U690 ( .A1(G92), .A2(n672), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n617), .B(KEYINPUT76), .ZN(n624) );
  NAND2_X1 U692 ( .A1(G79), .A2(n667), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G66), .A2(n663), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G54), .A2(n664), .ZN(n620) );
  XNOR2_X1 U696 ( .A(KEYINPUT77), .B(n620), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U699 ( .A(KEYINPUT15), .B(n625), .ZN(n971) );
  OR2_X1 U700 ( .A1(n971), .A2(G868), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(G284) );
  NAND2_X1 U702 ( .A1(G65), .A2(n663), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G53), .A2(n664), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U705 ( .A1(G78), .A2(n667), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G91), .A2(n672), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n726) );
  INV_X1 U709 ( .A(n726), .ZN(G299) );
  INV_X1 U710 ( .A(G868), .ZN(n634) );
  NOR2_X1 U711 ( .A1(G286), .A2(n634), .ZN(n636) );
  NOR2_X1 U712 ( .A1(G868), .A2(G299), .ZN(n635) );
  NOR2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U714 ( .A(KEYINPUT79), .B(n637), .Z(G297) );
  NAND2_X1 U715 ( .A1(n638), .A2(G559), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n639), .A2(n971), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U718 ( .A1(G868), .A2(n963), .ZN(n641) );
  XNOR2_X1 U719 ( .A(KEYINPUT80), .B(n641), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G868), .A2(n971), .ZN(n642) );
  NOR2_X1 U721 ( .A1(G559), .A2(n642), .ZN(n643) );
  NOR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(G282) );
  NAND2_X1 U723 ( .A1(n672), .A2(G93), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n645), .B(KEYINPUT82), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G67), .A2(n663), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U727 ( .A1(G80), .A2(n667), .ZN(n649) );
  NAND2_X1 U728 ( .A1(G55), .A2(n664), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n682) );
  NAND2_X1 U731 ( .A1(G559), .A2(n971), .ZN(n652) );
  XOR2_X1 U732 ( .A(n963), .B(n652), .Z(n680) );
  XNOR2_X1 U733 ( .A(KEYINPUT81), .B(n680), .ZN(n653) );
  NOR2_X1 U734 ( .A1(G860), .A2(n653), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n682), .B(n654), .ZN(G145) );
  NAND2_X1 U736 ( .A1(n664), .A2(G49), .ZN(n655) );
  XOR2_X1 U737 ( .A(KEYINPUT83), .B(n655), .Z(n657) );
  NAND2_X1 U738 ( .A1(G651), .A2(G74), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U740 ( .A(KEYINPUT84), .B(n658), .ZN(n659) );
  NOR2_X1 U741 ( .A1(n663), .A2(n659), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n660), .A2(G87), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n662), .A2(n661), .ZN(G288) );
  NAND2_X1 U744 ( .A1(G61), .A2(n663), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G48), .A2(n664), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n671) );
  NAND2_X1 U747 ( .A1(G73), .A2(n667), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(KEYINPUT85), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n669), .B(KEYINPUT2), .ZN(n670) );
  NOR2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n674) );
  NAND2_X1 U751 ( .A1(n672), .A2(G86), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n674), .A2(n673), .ZN(G305) );
  XOR2_X1 U753 ( .A(G303), .B(G288), .Z(n679) );
  XOR2_X1 U754 ( .A(G299), .B(n682), .Z(n677) );
  XOR2_X1 U755 ( .A(KEYINPUT19), .B(G305), .Z(n675) );
  XNOR2_X1 U756 ( .A(G290), .B(n675), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U758 ( .A(n679), .B(n678), .ZN(n919) );
  XNOR2_X1 U759 ( .A(n680), .B(n919), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n681), .A2(G868), .ZN(n684) );
  OR2_X1 U761 ( .A1(G868), .A2(n682), .ZN(n683) );
  NAND2_X1 U762 ( .A1(n684), .A2(n683), .ZN(G295) );
  NAND2_X1 U763 ( .A1(G2084), .A2(G2078), .ZN(n685) );
  XOR2_X1 U764 ( .A(KEYINPUT20), .B(n685), .Z(n686) );
  NAND2_X1 U765 ( .A1(G2090), .A2(n686), .ZN(n687) );
  XNOR2_X1 U766 ( .A(KEYINPUT21), .B(n687), .ZN(n688) );
  NAND2_X1 U767 ( .A1(n688), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U768 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U769 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NOR2_X1 U770 ( .A1(G219), .A2(G220), .ZN(n689) );
  XOR2_X1 U771 ( .A(KEYINPUT22), .B(n689), .Z(n690) );
  NOR2_X1 U772 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U773 ( .A1(G96), .A2(n691), .ZN(n858) );
  NAND2_X1 U774 ( .A1(n858), .A2(G2106), .ZN(n695) );
  NAND2_X1 U775 ( .A1(G69), .A2(G120), .ZN(n692) );
  NOR2_X1 U776 ( .A1(G237), .A2(n692), .ZN(n693) );
  NAND2_X1 U777 ( .A1(G108), .A2(n693), .ZN(n859) );
  NAND2_X1 U778 ( .A1(n859), .A2(G567), .ZN(n694) );
  NAND2_X1 U779 ( .A1(n695), .A2(n694), .ZN(n932) );
  NAND2_X1 U780 ( .A1(G483), .A2(G661), .ZN(n696) );
  NOR2_X1 U781 ( .A1(n932), .A2(n696), .ZN(n857) );
  NAND2_X1 U782 ( .A1(n857), .A2(G36), .ZN(G176) );
  INV_X1 U783 ( .A(G1384), .ZN(n698) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n812) );
  NOR2_X2 U785 ( .A1(n810), .A2(n812), .ZN(n731) );
  NAND2_X1 U786 ( .A1(n731), .A2(G1996), .ZN(n700) );
  XNOR2_X1 U787 ( .A(n700), .B(KEYINPUT26), .ZN(n702) );
  AND2_X1 U788 ( .A1(KEYINPUT26), .A2(G1341), .ZN(n701) );
  NAND2_X1 U789 ( .A1(n749), .A2(n701), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n702), .A2(n705), .ZN(n704) );
  INV_X1 U791 ( .A(KEYINPUT101), .ZN(n703) );
  NAND2_X1 U792 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U793 ( .A1(n705), .A2(KEYINPUT101), .ZN(n707) );
  INV_X1 U794 ( .A(n963), .ZN(n706) );
  XNOR2_X1 U795 ( .A(n709), .B(KEYINPUT103), .ZN(n717) );
  NAND2_X1 U796 ( .A1(n710), .A2(n971), .ZN(n715) );
  INV_X1 U797 ( .A(G2067), .ZN(n860) );
  NOR2_X1 U798 ( .A1(n749), .A2(n860), .ZN(n711) );
  XOR2_X1 U799 ( .A(n711), .B(KEYINPUT102), .Z(n713) );
  NAND2_X1 U800 ( .A1(n749), .A2(G1348), .ZN(n712) );
  NAND2_X1 U801 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U803 ( .A1(n717), .A2(n716), .ZN(n724) );
  INV_X1 U804 ( .A(KEYINPUT27), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n731), .A2(G2072), .ZN(n718) );
  XNOR2_X1 U806 ( .A(n719), .B(n718), .ZN(n721) );
  NAND2_X1 U807 ( .A1(G1956), .A2(n749), .ZN(n720) );
  NAND2_X1 U808 ( .A1(n726), .A2(n725), .ZN(n723) );
  NAND2_X1 U809 ( .A1(n724), .A2(n723), .ZN(n729) );
  NOR2_X1 U810 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U811 ( .A(n727), .B(KEYINPUT28), .Z(n728) );
  NAND2_X1 U812 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U813 ( .A(n730), .B(KEYINPUT29), .ZN(n736) );
  XOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .Z(n1015) );
  NOR2_X1 U815 ( .A1(n1015), .A2(n749), .ZN(n733) );
  NOR2_X1 U816 ( .A1(n731), .A2(G1961), .ZN(n732) );
  NOR2_X1 U817 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U818 ( .A(KEYINPUT99), .B(n734), .ZN(n741) );
  AND2_X1 U819 ( .A1(G171), .A2(n741), .ZN(n735) );
  NOR2_X1 U820 ( .A1(n736), .A2(n735), .ZN(n746) );
  NAND2_X1 U821 ( .A1(G8), .A2(n749), .ZN(n840) );
  NOR2_X1 U822 ( .A1(G1966), .A2(n840), .ZN(n762) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n749), .ZN(n759) );
  NOR2_X1 U824 ( .A1(n762), .A2(n759), .ZN(n737) );
  NAND2_X1 U825 ( .A1(G8), .A2(n737), .ZN(n739) );
  NOR2_X1 U826 ( .A1(G168), .A2(n740), .ZN(n743) );
  NOR2_X1 U827 ( .A1(G171), .A2(n741), .ZN(n742) );
  NOR2_X1 U828 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U829 ( .A(n744), .B(KEYINPUT31), .ZN(n745) );
  NOR2_X1 U830 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U831 ( .A(n747), .B(KEYINPUT105), .ZN(n758) );
  AND2_X1 U832 ( .A1(G286), .A2(G8), .ZN(n748) );
  NAND2_X1 U833 ( .A1(n758), .A2(n748), .ZN(n756) );
  INV_X1 U834 ( .A(G8), .ZN(n754) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n840), .ZN(n751) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n749), .ZN(n750) );
  NOR2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n752), .A2(G303), .ZN(n753) );
  OR2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n755) );
  AND2_X1 U840 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U841 ( .A(n757), .B(KEYINPUT32), .ZN(n786) );
  XNOR2_X1 U842 ( .A(n758), .B(KEYINPUT106), .ZN(n764) );
  NAND2_X1 U843 ( .A1(n759), .A2(G8), .ZN(n760) );
  XOR2_X1 U844 ( .A(KEYINPUT98), .B(n760), .Z(n761) );
  NOR2_X1 U845 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U846 ( .A1(n764), .A2(n763), .ZN(n784) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n774) );
  INV_X1 U848 ( .A(n840), .ZN(n767) );
  NAND2_X1 U849 ( .A1(n774), .A2(n767), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n765), .A2(KEYINPUT33), .ZN(n775) );
  INV_X1 U851 ( .A(n775), .ZN(n770) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n976) );
  AND2_X1 U854 ( .A1(n766), .A2(n976), .ZN(n768) );
  AND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  OR2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n772) );
  AND2_X1 U857 ( .A1(n784), .A2(n772), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n786), .A2(n771), .ZN(n779) );
  INV_X1 U859 ( .A(n772), .ZN(n777) );
  NOR2_X1 U860 ( .A1(G1971), .A2(G303), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n972) );
  AND2_X1 U862 ( .A1(n972), .A2(n775), .ZN(n776) );
  OR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U865 ( .A(n780), .B(KEYINPUT107), .ZN(n781) );
  XNOR2_X1 U866 ( .A(G1981), .B(G305), .ZN(n961) );
  NOR2_X2 U867 ( .A1(n781), .A2(n961), .ZN(n783) );
  XNOR2_X1 U868 ( .A(n783), .B(n782), .ZN(n842) );
  BUF_X1 U869 ( .A(n784), .Z(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n789) );
  NOR2_X1 U871 ( .A1(G2090), .A2(G303), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G8), .A2(n787), .ZN(n788) );
  NAND2_X1 U873 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n790), .A2(n840), .ZN(n837) );
  XOR2_X1 U875 ( .A(KEYINPUT39), .B(KEYINPUT109), .Z(n820) );
  NAND2_X1 U876 ( .A1(n907), .A2(G105), .ZN(n791) );
  XNOR2_X1 U877 ( .A(KEYINPUT38), .B(n791), .ZN(n800) );
  NAND2_X1 U878 ( .A1(n567), .A2(G141), .ZN(n792) );
  XNOR2_X1 U879 ( .A(n792), .B(KEYINPUT97), .ZN(n798) );
  NAND2_X1 U880 ( .A1(n903), .A2(G117), .ZN(n793) );
  XOR2_X1 U881 ( .A(KEYINPUT95), .B(n793), .Z(n795) );
  NAND2_X1 U882 ( .A1(n904), .A2(G129), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U884 ( .A(KEYINPUT96), .B(n796), .ZN(n797) );
  NOR2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n898) );
  NOR2_X1 U887 ( .A1(G1996), .A2(n898), .ZN(n945) );
  XOR2_X1 U888 ( .A(KEYINPUT94), .B(G1991), .Z(n1016) );
  NAND2_X1 U889 ( .A1(G107), .A2(n903), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G119), .A2(n904), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n805) );
  NAND2_X1 U892 ( .A1(G131), .A2(n567), .ZN(n803) );
  XNOR2_X1 U893 ( .A(KEYINPUT93), .B(n803), .ZN(n804) );
  NOR2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n907), .A2(G95), .ZN(n806) );
  AND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n915) );
  NOR2_X1 U897 ( .A1(n1016), .A2(n915), .ZN(n809) );
  AND2_X1 U898 ( .A1(n898), .A2(G1996), .ZN(n808) );
  NOR2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n943) );
  INV_X1 U900 ( .A(n943), .ZN(n814) );
  INV_X1 U901 ( .A(n810), .ZN(n811) );
  NOR2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U903 ( .A(n813), .B(KEYINPUT90), .ZN(n844) );
  NAND2_X1 U904 ( .A1(n814), .A2(n844), .ZN(n847) );
  INV_X1 U905 ( .A(n847), .ZN(n817) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n815) );
  AND2_X1 U907 ( .A1(n1016), .A2(n915), .ZN(n941) );
  NOR2_X1 U908 ( .A1(n815), .A2(n941), .ZN(n816) );
  NOR2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U910 ( .A1(n945), .A2(n818), .ZN(n819) );
  XNOR2_X1 U911 ( .A(n820), .B(n819), .ZN(n832) );
  XOR2_X1 U912 ( .A(n860), .B(KEYINPUT37), .Z(n834) );
  NAND2_X1 U913 ( .A1(n907), .A2(G104), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G140), .A2(n567), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U916 ( .A(n823), .B(KEYINPUT91), .ZN(n824) );
  XNOR2_X1 U917 ( .A(n824), .B(KEYINPUT34), .ZN(n830) );
  XNOR2_X1 U918 ( .A(KEYINPUT92), .B(KEYINPUT35), .ZN(n828) );
  NAND2_X1 U919 ( .A1(G116), .A2(n903), .ZN(n826) );
  NAND2_X1 U920 ( .A1(G128), .A2(n904), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U924 ( .A(KEYINPUT36), .B(n831), .Z(n897) );
  NOR2_X1 U925 ( .A1(n834), .A2(n897), .ZN(n953) );
  NAND2_X1 U926 ( .A1(n953), .A2(n844), .ZN(n846) );
  NAND2_X1 U927 ( .A1(n832), .A2(n846), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n833), .B(KEYINPUT110), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n834), .A2(n897), .ZN(n950) );
  NAND2_X1 U930 ( .A1(n835), .A2(n950), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n836), .A2(n844), .ZN(n843) );
  AND2_X1 U932 ( .A1(n837), .A2(n843), .ZN(n841) );
  NOR2_X1 U933 ( .A1(G1981), .A2(G305), .ZN(n838) );
  XOR2_X1 U934 ( .A(n838), .B(KEYINPUT24), .Z(n839) );
  NAND2_X1 U935 ( .A1(n842), .A2(n525), .ZN(n852) );
  INV_X1 U936 ( .A(n843), .ZN(n850) );
  XNOR2_X1 U937 ( .A(G1986), .B(G290), .ZN(n968) );
  NAND2_X1 U938 ( .A1(n968), .A2(n844), .ZN(n845) );
  AND2_X1 U939 ( .A1(n846), .A2(n845), .ZN(n848) );
  AND2_X1 U940 ( .A1(n848), .A2(n847), .ZN(n849) );
  OR2_X1 U941 ( .A1(n850), .A2(n849), .ZN(n851) );
  AND2_X1 U942 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U943 ( .A(n853), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n854), .ZN(G217) );
  INV_X1 U945 ( .A(n854), .ZN(G223) );
  AND2_X1 U946 ( .A1(G15), .A2(G2), .ZN(n855) );
  NAND2_X1 U947 ( .A1(G661), .A2(n855), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n856) );
  NAND2_X1 U949 ( .A1(n857), .A2(n856), .ZN(G188) );
  INV_X1 U951 ( .A(G120), .ZN(G236) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  INV_X1 U953 ( .A(G69), .ZN(G235) );
  NOR2_X1 U954 ( .A1(n859), .A2(n858), .ZN(G325) );
  INV_X1 U955 ( .A(G325), .ZN(G261) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2090), .Z(n862) );
  XOR2_X1 U957 ( .A(G2084), .B(n860), .Z(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U959 ( .A(n863), .B(G2100), .Z(n865) );
  XNOR2_X1 U960 ( .A(G2078), .B(G2072), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U962 ( .A(G2096), .B(KEYINPUT43), .Z(n867) );
  XNOR2_X1 U963 ( .A(G2678), .B(KEYINPUT113), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U965 ( .A(n869), .B(n868), .Z(G227) );
  XOR2_X1 U966 ( .A(G1976), .B(G1971), .Z(n871) );
  XNOR2_X1 U967 ( .A(G1966), .B(G1956), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U969 ( .A(n872), .B(KEYINPUT41), .Z(n874) );
  XNOR2_X1 U970 ( .A(G1961), .B(G1986), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U972 ( .A(G2474), .B(G1991), .Z(n876) );
  XNOR2_X1 U973 ( .A(G1996), .B(G1981), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(G229) );
  NAND2_X1 U976 ( .A1(G124), .A2(n904), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n879), .B(KEYINPUT44), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n880), .B(KEYINPUT114), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G112), .A2(n903), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U981 ( .A1(n907), .A2(G100), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G136), .A2(n567), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(G162) );
  XOR2_X1 U985 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n888) );
  XNOR2_X1 U986 ( .A(G162), .B(KEYINPUT115), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U988 ( .A(G160), .B(n889), .ZN(n902) );
  NAND2_X1 U989 ( .A1(n907), .A2(G103), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G139), .A2(n567), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G115), .A2(n903), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G127), .A2(n904), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n933) );
  XNOR2_X1 U997 ( .A(n897), .B(n933), .ZN(n900) );
  XOR2_X1 U998 ( .A(G164), .B(n898), .Z(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n917) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n903), .ZN(n906) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n904), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n912) );
  NAND2_X1 U1004 ( .A1(n907), .A2(G106), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(G142), .A2(n567), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1007 ( .A(n910), .B(KEYINPUT45), .Z(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n913), .B(n939), .ZN(n914) );
  XOR2_X1 U1010 ( .A(n915), .B(n914), .Z(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n918), .ZN(G395) );
  XOR2_X1 U1013 ( .A(KEYINPUT116), .B(n919), .Z(n921) );
  XOR2_X1 U1014 ( .A(G301), .B(G286), .Z(n920) );
  XNOR2_X1 U1015 ( .A(n921), .B(n920), .ZN(n923) );
  XOR2_X1 U1016 ( .A(n963), .B(n971), .Z(n922) );
  XNOR2_X1 U1017 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n924), .ZN(G397) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n932), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(KEYINPUT117), .B(n925), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n926), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(KEYINPUT118), .B(n929), .ZN(n931) );
  NOR2_X1 U1025 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(n932), .ZN(G319) );
  INV_X1 U1029 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1030 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1033 ( .A(KEYINPUT50), .B(n936), .Z(n956) );
  XOR2_X1 U1034 ( .A(G160), .B(G2084), .Z(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT119), .B(n937), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n949) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1041 ( .A(KEYINPUT120), .B(n946), .Z(n947) );
  XOR2_X1 U1042 ( .A(KEYINPUT51), .B(n947), .Z(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(KEYINPUT121), .B(n954), .ZN(n955) );
  NOR2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n957), .ZN(n958) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n1029) );
  NAND2_X1 U1050 ( .A1(n958), .A2(n1029), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n959), .A2(G29), .ZN(n1038) );
  INV_X1 U1052 ( .A(G16), .ZN(n1009) );
  XOR2_X1 U1053 ( .A(n1009), .B(KEYINPUT56), .Z(n984) );
  XOR2_X1 U1054 ( .A(G168), .B(G1966), .Z(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1056 ( .A(KEYINPUT57), .B(n962), .Z(n982) );
  XNOR2_X1 U1057 ( .A(G1341), .B(KEYINPUT124), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(n963), .ZN(n980) );
  XOR2_X1 U1059 ( .A(G301), .B(G1961), .Z(n970) );
  XOR2_X1 U1060 ( .A(G299), .B(G1956), .Z(n966) );
  NAND2_X1 U1061 ( .A1(G1971), .A2(G303), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(G1348), .B(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT123), .B(n978), .Z(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n1011) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G22), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G1976), .B(G23), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1076 ( .A(KEYINPUT126), .B(n987), .Z(n989) );
  XNOR2_X1 U1077 ( .A(G1986), .B(G24), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT58), .B(n990), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G21), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G1961), .B(G5), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n1005) );
  XNOR2_X1 U1084 ( .A(KEYINPUT59), .B(G4), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(KEYINPUT125), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G1348), .B(n996), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G1981), .B(G6), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G20), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(n1006), .B(KEYINPUT127), .Z(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1036) );
  XNOR2_X1 U1099 ( .A(G1996), .B(G32), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G33), .B(G2072), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1022) );
  XOR2_X1 U1102 ( .A(G26), .B(G2067), .Z(n1014) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(G28), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(n1015), .B(G27), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(n1016), .B(G25), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(n1023), .B(KEYINPUT53), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(G2084), .B(G34), .Z(n1024) );
  XNOR2_X1 U1111 ( .A(KEYINPUT54), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(G35), .B(G2090), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1030) );
  XOR2_X1 U1115 ( .A(n1030), .B(n1029), .Z(n1032) );
  INV_X1 U1116 ( .A(G29), .ZN(n1031) );
  NAND2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1118 ( .A1(G11), .A2(n1033), .ZN(n1034) );
  XNOR2_X1 U1119 ( .A(KEYINPUT122), .B(n1034), .ZN(n1035) );
  NOR2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1121 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1039), .ZN(G150) );
  INV_X1 U1123 ( .A(G150), .ZN(G311) );
  INV_X1 U1124 ( .A(G303), .ZN(G166) );
endmodule

