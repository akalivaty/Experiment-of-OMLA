//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT69), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G116), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT68), .B(G119), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G116), .ZN(new_n201));
  INV_X1    g015(.A(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G113), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n197), .B1(new_n201), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n198), .A2(KEYINPUT68), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n210), .A3(G116), .ZN(new_n211));
  INV_X1    g025(.A(new_n199), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n206), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(KEYINPUT69), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT71), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT70), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n201), .A2(new_n218), .A3(new_n206), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n212), .A3(new_n206), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT70), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n216), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n217), .B1(new_n216), .B2(new_n222), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT0), .B(G128), .Z(new_n225));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G143), .B(G146), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT0), .B(G128), .C1(new_n233), .C2(KEYINPUT64), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT11), .ZN(new_n236));
  INV_X1    g050(.A(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G134), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n240), .A3(G137), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n237), .A2(G137), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n236), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n238), .A2(new_n240), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT11), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT65), .B(G134), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n236), .B1(new_n250), .B2(G137), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n242), .B1(new_n250), .B2(G137), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n249), .B(new_n251), .C1(new_n252), .C2(new_n236), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n235), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n228), .A3(new_n230), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n233), .A2(new_n259), .A3(new_n256), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n229), .A2(KEYINPUT1), .A3(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n231), .A2(new_n255), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n258), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n250), .A2(G137), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n246), .A2(G134), .ZN(new_n265));
  OAI21_X1  g079(.A(G131), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n253), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n223), .A2(new_n224), .B1(new_n254), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT69), .B1(new_n213), .B2(new_n214), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n197), .B(new_n206), .C1(new_n211), .C2(new_n212), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n218), .B1(new_n201), .B2(new_n206), .ZN(new_n271));
  AND4_X1   g085(.A1(new_n218), .A2(new_n211), .A3(new_n212), .A4(new_n206), .ZN(new_n272));
  OAI22_X1  g086(.A1(new_n269), .A2(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT71), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n216), .A2(new_n217), .A3(new_n222), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n248), .A2(new_n253), .ZN(new_n276));
  INV_X1    g090(.A(new_n235), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n253), .A2(new_n263), .A3(new_n266), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n274), .A2(new_n275), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n268), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT28), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n196), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n268), .B2(new_n280), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(KEYINPUT74), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT75), .B(new_n195), .C1(new_n285), .C2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n267), .A2(new_n254), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT67), .B1(new_n289), .B2(KEYINPUT30), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n291), .B(new_n292), .C1(new_n267), .C2(new_n254), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n278), .A2(KEYINPUT30), .A3(new_n279), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n289), .A2(KEYINPUT72), .A3(KEYINPUT30), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n290), .A2(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n274), .A2(new_n275), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n280), .A2(new_n194), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n280), .A2(KEYINPUT73), .A3(new_n194), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n298), .A2(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n290), .A2(new_n293), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n296), .A2(new_n297), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n299), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT31), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n288), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n280), .A2(new_n283), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT74), .B1(new_n286), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n282), .A2(new_n196), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT75), .B1(new_n317), .B2(new_n195), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n187), .B(new_n188), .C1(new_n313), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n282), .A2(new_n284), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n287), .B1(new_n323), .B2(KEYINPUT74), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n324), .B2(new_n194), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n307), .A2(new_n305), .A3(new_n310), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n305), .B1(new_n307), .B2(new_n310), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n328), .A3(new_n288), .ZN(new_n329));
  NOR2_X1   g143(.A1(G472), .A2(G902), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n320), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n282), .A2(KEYINPUT29), .A3(new_n284), .A4(new_n194), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n334));
  AOI21_X1  g148(.A(G902), .B1(new_n333), .B2(KEYINPUT76), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n336));
  INV_X1    g150(.A(new_n280), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n298), .B2(new_n299), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n338), .B2(new_n194), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n285), .A2(new_n287), .A3(new_n195), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n334), .B(new_n335), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n329), .A2(new_n332), .B1(new_n341), .B2(G472), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n321), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G214), .B1(G237), .B2(G902), .ZN(new_n344));
  XNOR2_X1  g158(.A(G110), .B(G122), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OR2_X1    g160(.A1(KEYINPUT85), .A2(G107), .ZN(new_n347));
  NAND2_X1  g161(.A1(KEYINPUT85), .A2(G107), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(G104), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G107), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT3), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT86), .B(G101), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT3), .B1(new_n350), .B2(G107), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n352), .A2(new_n356), .ZN(new_n359));
  INV_X1    g173(.A(G101), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n357), .A2(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(KEYINPUT4), .B(G101), .C1(new_n352), .C2(new_n356), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n274), .A2(new_n275), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n351), .ZN(new_n364));
  AND2_X1   g178(.A1(KEYINPUT85), .A2(G107), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT85), .A2(G107), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n367), .B2(G104), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n353), .B(new_n355), .C1(new_n368), .C2(KEYINPUT3), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n367), .A2(G104), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n350), .A2(G107), .ZN(new_n371));
  OAI21_X1  g185(.A(G101), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n211), .A2(KEYINPUT5), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(new_n202), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(new_n213), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n222), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n346), .B1(new_n363), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n361), .A2(new_n362), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n223), .B2(new_n224), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n345), .A3(new_n378), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n383), .A3(KEYINPUT6), .ZN(new_n384));
  AND2_X1   g198(.A1(KEYINPUT78), .A2(G125), .ZN(new_n385));
  NOR2_X1   g199(.A1(KEYINPUT78), .A2(G125), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n263), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n387), .B2(new_n235), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n190), .A2(G224), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n392), .B(new_n346), .C1(new_n363), .C2(new_n379), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G210), .B1(G237), .B2(G902), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n390), .A2(KEYINPUT7), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n389), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n373), .A2(new_n222), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n375), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n213), .A2(new_n376), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n374), .A2(KEYINPUT89), .A3(new_n202), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n377), .A2(new_n222), .ZN(new_n404));
  OAI22_X1  g218(.A1(new_n398), .A2(new_n403), .B1(new_n404), .B2(new_n373), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n345), .B(KEYINPUT8), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n397), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n407), .B2(new_n383), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n394), .A2(new_n395), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n395), .B1(new_n394), .B2(new_n408), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n344), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n189), .A2(new_n190), .A3(G214), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(new_n229), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT18), .A2(G131), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G125), .B(G140), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n417), .A2(new_n227), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n419));
  INV_X1    g233(.A(G125), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT78), .A2(G125), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n421), .A2(KEYINPUT79), .A3(G140), .A4(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G140), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n385), .A2(new_n386), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT79), .B1(new_n424), .B2(G125), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n423), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(new_n227), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n416), .B1(new_n418), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G113), .B(G122), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(G104), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT92), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n414), .A2(KEYINPUT17), .A3(G131), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n414), .A2(G131), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n414), .A2(G131), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n434), .B1(new_n437), .B2(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n428), .A2(KEYINPUT16), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n387), .A2(KEYINPUT16), .A3(G140), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(G146), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT16), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n421), .A2(G140), .A3(new_n422), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n426), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n445), .B2(new_n423), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n227), .B1(new_n446), .B2(new_n440), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n430), .B(new_n433), .C1(new_n438), .C2(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n446), .A2(new_n227), .A3(new_n440), .ZN(new_n450));
  OAI211_X1 g264(.A(KEYINPUT19), .B(new_n423), .C1(new_n425), .C2(new_n427), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n417), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n451), .A2(new_n227), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT90), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n227), .A3(new_n453), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n442), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n437), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n430), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n432), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n459), .B2(new_n430), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n449), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n465));
  NOR2_X1   g279(.A1(G475), .A2(G902), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(KEYINPUT93), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n470), .B(new_n449), .C1(new_n462), .C2(new_n463), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n468), .B1(new_n472), .B2(KEYINPUT20), .ZN(new_n473));
  INV_X1    g287(.A(new_n432), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n430), .B1(new_n438), .B2(new_n448), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n476), .B2(new_n475), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n449), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n188), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n480), .A2(G475), .ZN(new_n481));
  INV_X1    g295(.A(new_n367), .ZN(new_n482));
  XOR2_X1   g296(.A(G116), .B(G122), .Z(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n229), .A2(G128), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n255), .A2(G143), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n250), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT13), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n486), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n485), .A2(new_n489), .ZN(new_n492));
  OAI21_X1  g306(.A(G134), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n485), .A2(new_n486), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n245), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G116), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT14), .A3(G122), .ZN(new_n499));
  OAI211_X1 g313(.A(G107), .B(new_n499), .C1(new_n483), .C2(KEYINPUT14), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n497), .B(new_n500), .C1(new_n482), .C2(new_n483), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n488), .A2(new_n493), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n501), .A2(new_n494), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT9), .B(G234), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT82), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(G217), .A3(new_n190), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n504), .B(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(G902), .ZN(new_n510));
  INV_X1    g324(.A(G478), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(KEYINPUT15), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n509), .B2(G902), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n190), .A2(G952), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(G234), .B2(G237), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n188), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT21), .B(G898), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  NOR4_X1   g335(.A1(new_n412), .A2(new_n473), .A3(new_n481), .A4(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g339(.A(KEYINPUT77), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n200), .B2(G128), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n208), .A2(new_n210), .A3(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT23), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n209), .A2(G119), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n198), .A2(KEYINPUT68), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT77), .B(new_n255), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n198), .A2(G128), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT23), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n200), .B2(G128), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT24), .B(G110), .Z(new_n538));
  AOI22_X1  g352(.A1(new_n536), .A2(G110), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n448), .A2(new_n539), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n536), .A2(G110), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n440), .B1(new_n428), .B2(KEYINPUT16), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n418), .B1(new_n542), .B2(G146), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n540), .A2(new_n544), .A3(KEYINPUT80), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT80), .B1(new_n540), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n525), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n525), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n544), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT80), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G217), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(G234), .B2(new_n188), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G902), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n547), .A2(new_n188), .A3(new_n551), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n547), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n551), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n559), .A2(KEYINPUT81), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n562), .A3(new_n558), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n554), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n556), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n369), .A2(new_n263), .A3(new_n372), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT87), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n369), .A2(new_n263), .A3(KEYINPUT87), .A4(new_n372), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n355), .B1(new_n368), .B2(KEYINPUT3), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n369), .A2(KEYINPUT4), .B1(new_n574), .B2(G101), .ZN(new_n575));
  INV_X1    g389(.A(new_n362), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n277), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n276), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n373), .A2(KEYINPUT10), .A3(new_n263), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n573), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT88), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n568), .A2(new_n571), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n381), .B2(new_n277), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n584), .A2(KEYINPUT88), .A3(new_n578), .A4(new_n573), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n570), .B(new_n572), .C1(new_n263), .C2(new_n373), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n276), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(KEYINPUT12), .A3(new_n276), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n190), .A2(G227), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT83), .ZN(new_n594));
  XNOR2_X1  g408(.A(G110), .B(G140), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n586), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n584), .A2(new_n573), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n276), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n596), .B1(new_n586), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n567), .B(new_n188), .C1(new_n597), .C2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n586), .A2(new_n596), .A3(new_n599), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n582), .A2(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n596), .B(KEYINPUT84), .Z(new_n604));
  OAI211_X1 g418(.A(new_n602), .B(G469), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n567), .A2(new_n188), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n601), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G221), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n506), .B2(new_n188), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n343), .A2(new_n522), .A3(new_n566), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n354), .ZN(G3));
  INV_X1    g428(.A(new_n319), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n187), .B1(new_n329), .B2(new_n188), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n617), .A2(new_n566), .A3(new_n612), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n504), .B(new_n507), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n619), .A2(KEYINPUT33), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(KEYINPUT33), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(G478), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n511), .A2(new_n188), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n510), .B2(new_n511), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n472), .A2(KEYINPUT20), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n467), .ZN(new_n627));
  INV_X1    g441(.A(new_n481), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n394), .A2(new_n408), .ZN(new_n630));
  INV_X1    g444(.A(new_n395), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n409), .ZN(new_n634));
  INV_X1    g448(.A(new_n344), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n411), .B2(KEYINPUT96), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n634), .A2(new_n520), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT97), .B1(new_n629), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n625), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n473), .B2(new_n481), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n634), .A2(new_n520), .A3(new_n636), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n618), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND4_X1  g460(.A1(new_n469), .A2(new_n465), .A3(new_n466), .A4(new_n471), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n481), .B1(new_n626), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n512), .A2(new_n514), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n641), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n618), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  AND2_X1   g468(.A1(new_n563), .A2(new_n554), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n559), .A2(KEYINPUT81), .A3(new_n560), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n549), .B(new_n657), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n655), .A2(new_n656), .B1(new_n555), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n617), .A2(new_n522), .A3(new_n612), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  AND3_X1   g477(.A1(new_n612), .A2(new_n634), .A3(new_n636), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n659), .B1(new_n321), .B2(new_n342), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n516), .B1(new_n517), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n650), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n671));
  INV_X1    g485(.A(new_n281), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n311), .B1(new_n672), .B2(new_n194), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n187), .B1(new_n673), .B2(new_n188), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n329), .B2(new_n332), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n321), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n671), .B1(new_n321), .B2(new_n675), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n659), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n667), .B(KEYINPUT39), .Z(new_n680));
  NAND2_X1  g494(.A1(new_n612), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n410), .A2(new_n411), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n473), .A2(new_n481), .ZN(new_n686));
  INV_X1    g500(.A(new_n649), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n685), .A2(new_n635), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n679), .A2(new_n682), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n229), .ZN(G45));
  INV_X1    g506(.A(new_n667), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n639), .B(new_n693), .C1(new_n473), .C2(new_n481), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n664), .A2(new_n665), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  NOR2_X1   g511(.A1(new_n567), .A2(KEYINPUT100), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n586), .A2(new_n599), .ZN(new_n699));
  INV_X1    g513(.A(new_n596), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n582), .B2(new_n585), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n699), .A2(new_n700), .B1(new_n701), .B2(new_n592), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n698), .B1(new_n702), .B2(G902), .ZN(new_n703));
  INV_X1    g517(.A(new_n698), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n188), .B(new_n704), .C1(new_n597), .C2(new_n600), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n705), .A3(new_n611), .ZN(new_n706));
  AOI211_X1 g520(.A(new_n565), .B(new_n706), .C1(new_n321), .C2(new_n342), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n638), .B2(new_n643), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT41), .B(G113), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT101), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n708), .B(new_n710), .ZN(G15));
  AOI21_X1  g525(.A(new_n565), .B1(new_n321), .B2(new_n342), .ZN(new_n712));
  INV_X1    g526(.A(new_n706), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n651), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NAND4_X1  g529(.A1(new_n627), .A2(new_n628), .A3(new_n687), .A4(new_n520), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n634), .A2(new_n636), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n717), .A3(new_n706), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n665), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n665), .A3(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  AOI21_X1  g538(.A(new_n194), .B1(new_n282), .B2(new_n284), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n311), .B2(KEYINPUT31), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n326), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT103), .B1(new_n327), .B2(new_n725), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n331), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n616), .A2(new_n730), .A3(new_n706), .A4(new_n565), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n634), .A2(new_n649), .A3(new_n636), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n732), .A2(new_n686), .A3(new_n519), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NOR2_X1   g549(.A1(new_n717), .A2(new_n706), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n188), .B1(new_n313), .B2(new_n318), .ZN(new_n737));
  INV_X1    g551(.A(new_n725), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n312), .A2(new_n727), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n306), .A3(new_n729), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n737), .A2(G472), .B1(new_n740), .B2(new_n330), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT104), .B1(new_n741), .B2(new_n660), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n616), .A2(new_n730), .A3(new_n659), .A4(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n695), .B(new_n736), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  NAND2_X1  g560(.A1(new_n343), .A2(new_n566), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT107), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n712), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n605), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n586), .A2(new_n592), .ZN(new_n753));
  INV_X1    g567(.A(new_n604), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(KEYINPUT105), .A3(G469), .A4(new_n602), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n752), .A2(new_n601), .A3(new_n607), .A4(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n410), .A2(new_n635), .A3(new_n411), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n611), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n694), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n748), .A2(new_n750), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n757), .A2(new_n611), .A3(new_n758), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n343), .A2(new_n763), .A3(new_n566), .A4(new_n695), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n764), .A2(KEYINPUT106), .A3(new_n760), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT106), .B1(new_n764), .B2(new_n760), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NAND3_X1  g582(.A1(new_n712), .A2(new_n668), .A3(new_n763), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NAND2_X1  g584(.A1(new_n686), .A2(new_n639), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT43), .Z(new_n772));
  NOR2_X1   g586(.A1(new_n617), .A2(new_n659), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT110), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT110), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n758), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n777), .A2(KEYINPUT111), .A3(new_n778), .A4(new_n758), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n755), .A2(new_n602), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT108), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n567), .B1(new_n783), .B2(new_n784), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n788), .A2(new_n789), .A3(new_n606), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n789), .B1(new_n788), .B2(new_n606), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n601), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n611), .A3(new_n680), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT109), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n774), .A2(new_n775), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n781), .A2(new_n782), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  INV_X1    g611(.A(new_n758), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n343), .A2(new_n566), .A3(new_n694), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n792), .A2(new_n611), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n800), .B1(new_n792), .B2(new_n611), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n806));
  NOR2_X1   g620(.A1(G952), .A2(G953), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT120), .Z(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n757), .A2(new_n611), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n810), .A2(new_n732), .A3(new_n686), .A4(new_n667), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n811), .B(new_n659), .C1(new_n676), .C2(new_n677), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n664), .B(new_n665), .C1(new_n668), .C2(new_n695), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n745), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n737), .A2(G472), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n740), .A2(new_n330), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n660), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n743), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n741), .A2(KEYINPUT104), .A3(new_n660), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n694), .B(new_n759), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n344), .B(new_n520), .C1(new_n410), .C2(new_n411), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n627), .A2(new_n628), .A3(new_n649), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n823), .B2(new_n640), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n617), .A3(new_n566), .A4(new_n612), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n613), .A3(new_n661), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n649), .A2(new_n667), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n648), .A2(new_n827), .A3(new_n758), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n343), .A2(new_n828), .A3(new_n612), .A4(new_n660), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n769), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n821), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n812), .A2(new_n745), .A3(new_n813), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n815), .A2(new_n831), .A3(new_n767), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n718), .A2(new_n665), .A3(KEYINPUT102), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT102), .B1(new_n718), .B2(new_n665), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n638), .A2(new_n643), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n712), .A2(new_n713), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n734), .B(new_n714), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT114), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n707), .A2(new_n651), .B1(new_n731), .B2(new_n733), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n723), .A2(new_n842), .A3(new_n708), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n809), .B1(new_n834), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT115), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n848), .B(new_n809), .C1(new_n834), .C2(new_n845), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n834), .A2(new_n845), .A3(new_n809), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT54), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n834), .A2(new_n845), .A3(new_n809), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(KEYINPUT115), .B2(new_n846), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n854), .B1(new_n856), .B2(new_n849), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n837), .A2(new_n840), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n767), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n826), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n819), .A2(new_n820), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n695), .A3(new_n763), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n769), .A3(new_n864), .A4(new_n829), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n809), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n831), .A2(KEYINPUT117), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n815), .A3(new_n833), .A4(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n854), .B(new_n846), .C1(new_n861), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT116), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n853), .B1(new_n857), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n792), .A2(new_n611), .ZN(new_n874));
  INV_X1    g688(.A(new_n800), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n703), .A2(new_n705), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n610), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n801), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n616), .A2(new_n730), .A3(new_n565), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n772), .A2(new_n516), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n798), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n772), .A2(new_n516), .A3(new_n731), .ZN(new_n884));
  INV_X1    g698(.A(new_n685), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n344), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT50), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n881), .A2(new_n706), .A3(new_n798), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n566), .A2(new_n758), .A3(new_n516), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n678), .A2(new_n706), .A3(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n639), .A2(new_n473), .A3(new_n481), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n890), .A2(new_n863), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n873), .B1(new_n883), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(KEYINPUT51), .A3(new_n889), .A4(new_n894), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n884), .A2(new_n634), .A3(new_n636), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n892), .A2(new_n629), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n515), .B(KEYINPUT119), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n748), .A2(new_n750), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n890), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n904), .A2(KEYINPUT48), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(KEYINPUT48), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n896), .A2(new_n898), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n808), .B1(new_n872), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n566), .A2(new_n344), .A3(new_n611), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT113), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n771), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT49), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n885), .B1(new_n913), .B2(new_n877), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n912), .B(new_n914), .C1(new_n913), .C2(new_n877), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n678), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n806), .B1(new_n909), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n916), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n896), .A2(new_n898), .A3(new_n907), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(KEYINPUT116), .A3(new_n870), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n921), .B2(new_n853), .ZN(new_n922));
  OAI211_X1 g736(.A(KEYINPUT121), .B(new_n918), .C1(new_n922), .C2(new_n808), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n917), .A2(new_n923), .ZN(G75));
  NOR2_X1   g738(.A1(new_n190), .A2(G952), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT122), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n846), .B1(new_n861), .B2(new_n869), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(G902), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT56), .B1(new_n929), .B2(G210), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n384), .A2(new_n393), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n391), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  OR2_X1    g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n933), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n927), .B1(new_n934), .B2(new_n935), .ZN(G51));
  NAND2_X1  g750(.A1(new_n928), .A2(KEYINPUT54), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n870), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n928), .A2(KEYINPUT123), .A3(KEYINPUT54), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n606), .B(KEYINPUT57), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n600), .B2(new_n597), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n929), .A2(new_n788), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n925), .B1(new_n943), .B2(new_n944), .ZN(G54));
  NAND3_X1  g759(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n469), .A2(new_n471), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n925), .ZN(G60));
  NAND2_X1  g764(.A1(new_n620), .A2(new_n621), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n623), .B(KEYINPUT59), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n939), .A2(new_n940), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n926), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n872), .A2(new_n953), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n952), .ZN(G63));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n928), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(new_n552), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n658), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n926), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n926), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(G66));
  INV_X1    g783(.A(new_n518), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n190), .B1(new_n970), .B2(G224), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n841), .A2(new_n844), .A3(new_n862), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT125), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n971), .B1(new_n974), .B2(new_n190), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n931), .B1(G898), .B2(new_n190), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  NAND2_X1  g792(.A1(new_n451), .A2(new_n453), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n298), .B(new_n979), .Z(new_n980));
  NAND2_X1  g794(.A1(new_n745), .A2(new_n813), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n691), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n823), .A2(new_n640), .ZN(new_n985));
  OR4_X1    g799(.A1(new_n747), .A2(new_n985), .A3(new_n681), .A4(new_n798), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n804), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n982), .A2(new_n983), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT127), .B1(new_n982), .B2(new_n983), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n796), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n980), .B1(new_n993), .B2(new_n190), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n980), .B1(new_n666), .B2(new_n190), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n732), .A2(new_n686), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n794), .A2(new_n996), .A3(new_n903), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n745), .A2(new_n813), .A3(new_n769), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n804), .A2(new_n767), .A3(new_n998), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n796), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n995), .B1(new_n1000), .B2(new_n190), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1002));
  OR3_X1    g816(.A1(new_n994), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n994), .B2(new_n1001), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(G72));
  OR2_X1    g819(.A1(new_n338), .A2(new_n194), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n992), .A2(new_n796), .A3(new_n973), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  AOI21_X1  g823(.A(new_n338), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n796), .A2(new_n973), .A3(new_n999), .A4(new_n997), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n194), .B1(new_n1011), .B2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1006), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1009), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n1006), .B2(new_n311), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n925), .B1(new_n851), .B2(new_n1015), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n1013), .A2(new_n1016), .ZN(G57));
endmodule


