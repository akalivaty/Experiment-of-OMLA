//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011;
  NAND2_X1  g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  OR2_X1    g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G57gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G64gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT95), .ZN(new_n208));
  INV_X1    g007(.A(G64gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G57gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT96), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n205), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n207), .A2(new_n210), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n202), .B(new_n203), .C1(new_n213), .C2(new_n204), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(KEYINPUT21), .ZN(new_n216));
  NAND2_X1  g015(.A1(G231gat), .A2(G233gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(G127gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(G1gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT16), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G1gat), .B2(new_n220), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(G8gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n225), .B1(KEYINPUT21), .B2(new_n215), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n219), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G183gat), .B(G211gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT97), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n229), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n227), .B(new_n233), .Z(new_n234));
  XOR2_X1   g033(.A(KEYINPUT89), .B(KEYINPUT15), .Z(new_n235));
  INV_X1    g034(.A(G50gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT90), .A3(G43gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(G43gat), .ZN(new_n238));
  INV_X1    g037(.A(G43gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G50gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n235), .B(new_n237), .C1(KEYINPUT90), .C2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G29gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n244));
  AND2_X1   g043(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n244), .B1(new_n247), .B2(G36gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT15), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n248), .A2(KEYINPUT15), .A3(new_n238), .A4(new_n240), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT17), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G85gat), .A2(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT7), .ZN(new_n257));
  NAND2_X1  g056(.A1(G99gat), .A2(G106gat), .ZN(new_n258));
  INV_X1    g057(.A(G85gat), .ZN(new_n259));
  INV_X1    g058(.A(G92gat), .ZN(new_n260));
  AOI22_X1  g059(.A1(KEYINPUT8), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G99gat), .B(G106gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT98), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n255), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n266), .B(new_n267), .C1(new_n253), .C2(new_n265), .ZN(new_n268));
  XNOR2_X1  g067(.A(G190gat), .B(G218gat), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G134gat), .B(G162gat), .Z(new_n271));
  AOI21_X1  g070(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT100), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n273), .A2(KEYINPUT100), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT99), .B1(new_n268), .B2(new_n269), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n268), .A2(KEYINPUT99), .A3(new_n269), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n275), .A2(new_n277), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n270), .A2(new_n280), .A3(new_n274), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n276), .B1(new_n282), .B2(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G230gat), .ZN(new_n285));
  INV_X1    g084(.A(G233gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n212), .A2(new_n214), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n264), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n264), .A2(KEYINPUT98), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n264), .A2(KEYINPUT98), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n292), .A2(KEYINPUT10), .A3(new_n215), .A4(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n287), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n289), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(new_n287), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G120gat), .B(G148gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G176gat), .B(G204gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  OR2_X1    g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n295), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n287), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n234), .A2(new_n284), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n225), .A2(new_n251), .A3(new_n252), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n308), .B(KEYINPUT91), .Z(new_n309));
  INV_X1    g108(.A(new_n225), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n253), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G229gat), .A2(G233gat), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n313), .B(KEYINPUT13), .Z(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT92), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n255), .A2(new_n310), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n309), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT18), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT92), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(new_n321), .A3(new_n314), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n309), .A2(KEYINPUT18), .A3(new_n313), .A4(new_n317), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n316), .A2(new_n320), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G113gat), .B(G141gat), .Z(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT88), .B(G197gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT11), .B(G169gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  XOR2_X1   g128(.A(new_n329), .B(KEYINPUT12), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n322), .A3(new_n323), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n320), .A2(KEYINPUT93), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT93), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n335), .A3(new_n319), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n330), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n332), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G228gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(new_n286), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G141gat), .B(G148gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(G155gat), .B2(G162gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n344), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G141gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G148gat), .ZN(new_n350));
  INV_X1    g149(.A(G148gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G141gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G155gat), .B(G162gat), .ZN(new_n354));
  INV_X1    g153(.A(G162gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT2), .B1(new_n231), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359));
  INV_X1    g158(.A(G197gat), .ZN(new_n360));
  INV_X1    g159(.A(G204gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT22), .ZN(new_n364));
  NAND2_X1  g163(.A1(G211gat), .A2(G218gat), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n362), .A2(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n367));
  XNOR2_X1  g166(.A(G211gat), .B(G218gat), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n364), .ZN(new_n370));
  NOR2_X1   g169(.A1(G197gat), .A2(G204gat), .ZN(new_n371));
  AND2_X1   g170(.A1(G197gat), .A2(G204gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G211gat), .B(G218gat), .Z(new_n374));
  AOI21_X1  g173(.A(KEYINPUT74), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n373), .B2(new_n374), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n366), .A2(KEYINPUT75), .A3(new_n368), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n359), .B1(new_n381), .B2(KEYINPUT80), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n363), .ZN(new_n384));
  AND4_X1   g183(.A1(KEYINPUT75), .A2(new_n384), .A3(new_n368), .A4(new_n370), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT75), .B1(new_n366), .B2(new_n368), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT74), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n383), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n358), .B1(new_n382), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n348), .A2(new_n357), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n359), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n383), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n387), .A2(new_n390), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n341), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n380), .B1(new_n368), .B2(new_n366), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n383), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n395), .B1(new_n402), .B2(new_n359), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n341), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(G22gat), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT3), .B1(new_n391), .B2(new_n392), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n381), .A2(KEYINPUT80), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n395), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n399), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n340), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G22gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n405), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  NAND3_X1  g216(.A1(new_n406), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n406), .A2(new_n414), .A3(KEYINPUT81), .A4(new_n417), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n414), .ZN(new_n424));
  INV_X1    g223(.A(new_n417), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI211_X1 g225(.A(KEYINPUT82), .B(new_n417), .C1(new_n406), .C2(new_n414), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n420), .A2(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G120gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT69), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT69), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G120gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n432), .A3(G113gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT70), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n429), .B2(G113gat), .ZN(new_n435));
  INV_X1    g234(.A(G113gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G134gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G127gat), .ZN(new_n440));
  INV_X1    g239(.A(G127gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G134gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT1), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n442), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n429), .A2(G113gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n436), .A2(G120gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n438), .A2(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G169gat), .ZN(new_n450));
  INV_X1    g249(.A(G176gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT23), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT23), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(G169gat), .B2(G176gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(G169gat), .A2(G176gat), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT25), .B(new_n452), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT24), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT24), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(G183gat), .A3(G190gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(G183gat), .A2(G190gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT67), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n456), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G183gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(KEYINPUT24), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n466), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n457), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT65), .B1(new_n467), .B2(new_n462), .ZN(new_n468));
  INV_X1    g267(.A(new_n455), .ZN(new_n469));
  NAND2_X1  g268(.A1(G169gat), .A2(G176gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT23), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n453), .A2(G169gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n451), .A2(KEYINPUT66), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT66), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G176gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n462), .B1(new_n458), .B2(new_n460), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT65), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n468), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n483));
  AOI21_X1  g282(.A(new_n464), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT26), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n485), .A3(new_n470), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n455), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT68), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n465), .A2(KEYINPUT27), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT27), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G183gat), .ZN(new_n492));
  INV_X1    g291(.A(G190gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT28), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT27), .B(G183gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT28), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n493), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT68), .B1(new_n486), .B2(new_n487), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n489), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n449), .B1(new_n484), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n472), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n503));
  AOI211_X1 g302(.A(KEYINPUT65), .B(new_n462), .C1(new_n458), .C2(new_n460), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n483), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n464), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n430), .A2(new_n432), .A3(G113gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n435), .A2(new_n437), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n444), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n448), .A2(new_n445), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n499), .A2(new_n500), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n488), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n507), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n502), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G227gat), .A2(G233gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT34), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n517), .B2(KEYINPUT72), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n518), .B(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n502), .A2(new_n515), .A3(G227gat), .A4(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G43gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G99gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(KEYINPUT71), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(KEYINPUT71), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(KEYINPUT33), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n523), .A2(KEYINPUT32), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(KEYINPUT32), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT33), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n523), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n534), .A3(new_n527), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n522), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n531), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n518), .B(new_n520), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n398), .ZN(new_n542));
  NAND2_X1  g341(.A1(G226gat), .A2(G233gat), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n505), .A2(new_n506), .B1(new_n513), .B2(new_n488), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(KEYINPUT29), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT76), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n543), .B1(new_n507), .B2(new_n514), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n383), .B1(new_n484), .B2(new_n501), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n542), .B(new_n546), .C1(new_n549), .C2(KEYINPUT76), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n545), .B1(new_n543), .B2(new_n544), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n398), .ZN(new_n552));
  XNOR2_X1  g351(.A(G8gat), .B(G36gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(G64gat), .B(G92gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n550), .A2(new_n552), .ZN(new_n559));
  INV_X1    g358(.A(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n557), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n550), .A2(new_n552), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G1gat), .B(G29gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT0), .ZN(new_n566));
  XNOR2_X1  g365(.A(G57gat), .B(G85gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT5), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n449), .B(new_n395), .ZN(new_n571));
  NAND2_X1  g370(.A1(G225gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n570), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT3), .A2(new_n358), .B1(new_n510), .B2(new_n511), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n573), .B1(new_n576), .B2(new_n396), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT4), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n449), .A2(new_n395), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT77), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT4), .B1(new_n512), .B2(new_n358), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n449), .A2(new_n395), .A3(KEYINPUT77), .A4(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n577), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n580), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n583), .A3(new_n582), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT78), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n577), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n575), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(KEYINPUT79), .A3(new_n579), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT79), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n449), .A2(new_n395), .A3(new_n593), .A4(new_n578), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n577), .A2(new_n570), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(KEYINPUT6), .B(new_n569), .C1(new_n591), .C2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n569), .B1(new_n591), .B2(new_n598), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT6), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n588), .A2(new_n589), .A3(new_n577), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n589), .B1(new_n588), .B2(new_n577), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n574), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n568), .A3(new_n597), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n564), .B1(new_n599), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT35), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n428), .A2(new_n541), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n400), .A2(G22gat), .A3(new_n405), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n425), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT82), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n424), .A2(new_n423), .A3(new_n425), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n418), .A2(new_n419), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n613), .A2(new_n614), .B1(new_n615), .B2(new_n421), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n606), .A2(new_n599), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n555), .B1(new_n550), .B2(new_n552), .ZN(new_n618));
  INV_X1    g417(.A(new_n559), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(new_n562), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n558), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n537), .A2(KEYINPUT73), .A3(new_n522), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n522), .B1(new_n537), .B2(KEYINPUT73), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n616), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n609), .B1(new_n625), .B2(new_n608), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n576), .A2(new_n396), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n592), .A2(new_n627), .A3(new_n594), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n573), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT83), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT83), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n631), .A3(new_n573), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n571), .A2(new_n573), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n630), .A2(KEYINPUT39), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n628), .A2(new_n631), .A3(new_n573), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(new_n628), .B2(new_n573), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n638), .A3(new_n568), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT84), .B(KEYINPUT40), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT85), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n634), .A2(new_n638), .A3(KEYINPUT40), .A4(new_n568), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n644), .A2(new_n600), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n639), .A2(KEYINPUT85), .A3(new_n640), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n643), .A2(new_n645), .A3(new_n564), .A4(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n555), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n559), .B2(new_n560), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n550), .B2(new_n552), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT38), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n652), .A2(new_n599), .A3(new_n606), .A4(new_n556), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n398), .B(new_n546), .C1(new_n549), .C2(KEYINPUT76), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n648), .B1(new_n551), .B2(new_n542), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT38), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n618), .B2(new_n649), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT86), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT86), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n656), .B(new_n659), .C1(new_n618), .C2(new_n649), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n428), .B(new_n647), .C1(new_n653), .C2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT36), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n536), .B2(new_n539), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT36), .B1(new_n622), .B2(new_n623), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n616), .A2(new_n621), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n626), .A2(KEYINPUT87), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT87), .B1(new_n626), .B2(new_n667), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n338), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT94), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT87), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n665), .A2(new_n664), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n428), .B2(new_n607), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n653), .A2(new_n661), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n643), .A2(new_n646), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n645), .A2(new_n564), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n616), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n624), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n428), .A2(new_n607), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n613), .A2(new_n614), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n615), .A2(new_n421), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n540), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n621), .A2(KEYINPUT35), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n682), .A2(KEYINPUT35), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n673), .B1(new_n680), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n626), .A2(KEYINPUT87), .A3(new_n667), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(KEYINPUT94), .A3(new_n338), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n307), .B1(new_n672), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n617), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n564), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT101), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  OAI211_X1 g499(.A(KEYINPUT101), .B(new_n700), .C1(new_n696), .C2(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(G8gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(G1325gat));
  INV_X1    g502(.A(new_n674), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n692), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  INV_X1    g505(.A(G15gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n707), .A3(new_n541), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n706), .A2(KEYINPUT102), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1326gat));
  NAND2_X1  g512(.A1(new_n692), .A2(new_n616), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  NOR2_X1   g515(.A1(new_n234), .A2(new_n305), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n281), .A2(new_n283), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n672), .B2(new_n691), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n243), .A3(new_n693), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n668), .B2(new_n669), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT44), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n626), .A2(new_n667), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n718), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT103), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n284), .B1(new_n626), .B2(new_n667), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n731), .A3(new_n727), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n725), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n338), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n617), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n722), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n738), .A3(new_n739), .ZN(G1328gat));
  NAND3_X1  g539(.A1(new_n734), .A2(new_n564), .A3(new_n736), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G36gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743));
  INV_X1    g542(.A(new_n564), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(G36gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n720), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n719), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT94), .B1(new_n690), .B2(new_n338), .ZN(new_n748));
  INV_X1    g547(.A(new_n338), .ZN(new_n749));
  AOI211_X1 g548(.A(new_n671), .B(new_n749), .C1(new_n688), .C2(new_n689), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n747), .B(new_n745), .C1(new_n748), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT46), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n742), .A2(new_n746), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n742), .A2(new_n755), .A3(new_n746), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1329gat));
  OAI21_X1  g556(.A(G43gat), .B1(new_n737), .B2(new_n674), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n720), .A2(new_n239), .A3(new_n541), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT47), .B1(new_n759), .B2(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n758), .B(new_n759), .C1(KEYINPUT105), .C2(KEYINPUT47), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1330gat));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n731), .B1(new_n730), .B2(new_n727), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n682), .A2(KEYINPUT35), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n767), .A2(new_n609), .B1(new_n662), .B2(new_n666), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n768), .A2(KEYINPUT103), .A3(KEYINPUT44), .A4(new_n284), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n727), .B1(new_n690), .B2(new_n718), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n616), .B(new_n736), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n428), .A2(G50gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(G50gat), .B1(new_n720), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n765), .B1(new_n774), .B2(KEYINPUT106), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n735), .B1(new_n725), .B2(new_n733), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n236), .B1(new_n777), .B2(new_n616), .ZN(new_n778));
  INV_X1    g577(.A(new_n773), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n719), .B(new_n779), .C1(new_n672), .C2(new_n691), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n776), .B(KEYINPUT48), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n775), .A2(new_n781), .ZN(G1331gat));
  INV_X1    g581(.A(new_n234), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n783), .A2(new_n718), .A3(new_n338), .A4(new_n306), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n726), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n617), .B(KEYINPUT107), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(new_n206), .ZN(G1332gat));
  NOR2_X1   g587(.A1(new_n785), .A2(new_n744), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  AND2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(G1333gat));
  NOR3_X1   g592(.A1(new_n785), .A2(G71gat), .A3(new_n540), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n726), .A2(new_n784), .A3(new_n704), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(G71gat), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g596(.A1(new_n785), .A2(new_n428), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT108), .B(G78gat), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1335gat));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n749), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n306), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n725), .B2(new_n733), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G85gat), .B1(new_n805), .B2(new_n617), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n730), .A2(new_n749), .A3(new_n783), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n306), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n259), .A3(new_n693), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n812), .ZN(G1336gat));
  NOR2_X1   g612(.A1(new_n744), .A2(G92gat), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n260), .B1(new_n804), .B2(new_n564), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n815), .B2(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1337gat));
  XNOR2_X1  g620(.A(KEYINPUT109), .B(G99gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n811), .A2(new_n541), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n805), .A2(new_n674), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n822), .ZN(G1338gat));
  NAND3_X1  g624(.A1(new_n734), .A2(new_n616), .A3(new_n802), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n804), .A2(KEYINPUT111), .A3(new_n616), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(G106gat), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n428), .A2(G106gat), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n811), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n826), .A2(G106gat), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT53), .B1(new_n836), .B2(new_n832), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1339gat));
  NOR2_X1   g637(.A1(new_n749), .A2(G113gat), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT114), .Z(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n334), .A2(new_n330), .A3(new_n336), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n316), .A2(new_n322), .A3(new_n323), .ZN(new_n843));
  INV_X1    g642(.A(new_n329), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n309), .A2(new_n317), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n845), .A2(new_n313), .B1(new_n312), .B2(new_n314), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n842), .A2(new_n843), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n718), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n291), .A2(new_n287), .A3(new_n294), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n302), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n300), .B1(new_n295), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(KEYINPUT55), .A3(new_n852), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n304), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n304), .A4(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n848), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n338), .A2(new_n858), .A3(new_n859), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n305), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n718), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n783), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n307), .A2(new_n338), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n564), .B(new_n786), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n616), .A2(new_n624), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n867), .A2(KEYINPUT113), .A3(new_n868), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n841), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n865), .A2(new_n866), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(new_n685), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n617), .A2(new_n564), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G113gat), .B1(new_n879), .B2(new_n749), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n874), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n880), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT115), .B1(new_n873), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1340gat));
  OAI21_X1  g683(.A(G120gat), .B1(new_n879), .B2(new_n306), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n871), .A2(new_n872), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n305), .A2(new_n430), .A3(new_n432), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT116), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(G1341gat));
  INV_X1    g688(.A(new_n869), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n441), .A3(new_n234), .ZN(new_n891));
  OAI21_X1  g690(.A(G127gat), .B1(new_n879), .B2(new_n783), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1342gat));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n439), .A3(new_n718), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n879), .B2(new_n284), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1343gat));
  NOR2_X1   g697(.A1(new_n307), .A2(new_n338), .ZN(new_n899));
  INV_X1    g698(.A(new_n856), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n338), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n718), .B1(new_n901), .B2(new_n863), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT117), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n338), .A2(new_n900), .B1(new_n847), .B2(new_n305), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n718), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n848), .A2(new_n860), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n899), .B1(new_n908), .B2(new_n783), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n428), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n674), .A2(new_n878), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n428), .B1(new_n865), .B2(new_n866), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G141gat), .B1(new_n915), .B2(new_n749), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n867), .A2(new_n616), .A3(new_n674), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n349), .A3(new_n338), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT58), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT58), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n916), .A2(new_n921), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1344gat));
  NAND3_X1  g722(.A1(new_n917), .A2(new_n351), .A3(new_n305), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925));
  AND4_X1   g724(.A1(new_n283), .A2(new_n847), .A3(new_n281), .A4(new_n900), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n783), .B1(new_n902), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n428), .B1(new_n927), .B2(new_n866), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT119), .B1(new_n928), .B2(KEYINPUT57), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n876), .A2(KEYINPUT57), .A3(new_n616), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n905), .A2(new_n718), .B1(new_n848), .B2(new_n856), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n899), .B1(new_n932), .B2(new_n783), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n931), .B(new_n913), .C1(new_n933), .C2(new_n428), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n306), .B1(new_n911), .B2(KEYINPUT118), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n935), .B(new_n936), .C1(KEYINPUT118), .C2(new_n911), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n925), .B1(new_n937), .B2(G148gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n910), .A2(new_n305), .A3(new_n914), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(new_n925), .A3(G148gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n924), .B1(new_n938), .B2(new_n940), .ZN(G1345gat));
  OAI21_X1  g740(.A(G155gat), .B1(new_n915), .B2(new_n783), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n917), .A2(new_n231), .A3(new_n234), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1346gat));
  NOR3_X1   g743(.A1(new_n915), .A2(new_n355), .A3(new_n284), .ZN(new_n945));
  AOI21_X1  g744(.A(G162gat), .B1(new_n917), .B2(new_n718), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(G1347gat));
  NAND2_X1  g746(.A1(new_n786), .A2(new_n564), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n877), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n950), .A2(new_n450), .A3(new_n749), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n876), .A2(KEYINPUT120), .A3(new_n617), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT120), .B1(new_n876), .B2(new_n617), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n868), .A2(new_n564), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT121), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n954), .A2(new_n338), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n951), .B1(new_n957), .B2(new_n450), .ZN(G1348gat));
  AOI211_X1 g757(.A(new_n306), .B(new_n950), .C1(new_n474), .C2(new_n476), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n305), .B(new_n956), .C1(new_n952), .C2(new_n953), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n962), .B2(G176gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(KEYINPUT122), .A3(new_n451), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(G1349gat));
  NAND4_X1  g764(.A1(new_n876), .A2(new_n685), .A3(new_n234), .A4(new_n949), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n465), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n234), .A2(new_n496), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n956), .B(new_n970), .C1(new_n952), .C2(new_n953), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n969), .A2(KEYINPUT124), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT60), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT60), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n969), .A2(KEYINPUT124), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n877), .A2(new_n718), .A3(new_n949), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n977), .A2(new_n978), .A3(G190gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n977), .B2(G190gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n954), .A2(new_n956), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n718), .A2(new_n493), .ZN(new_n982));
  OAI22_X1  g781(.A1(new_n979), .A2(new_n980), .B1(new_n981), .B2(new_n982), .ZN(G1351gat));
  NOR2_X1   g782(.A1(new_n948), .A2(new_n704), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n935), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n985), .A2(new_n360), .A3(new_n749), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n704), .A2(new_n428), .A3(new_n744), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n954), .A2(new_n338), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n986), .B1(new_n360), .B2(new_n988), .ZN(G1352gat));
  XNOR2_X1  g788(.A(KEYINPUT125), .B(G204gat), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n306), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n987), .B(new_n991), .C1(new_n952), .C2(new_n953), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(KEYINPUT126), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n990), .B1(new_n985), .B2(new_n306), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n992), .A2(new_n997), .A3(KEYINPUT62), .ZN(new_n998));
  NAND4_X1  g797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n998), .ZN(G1353gat));
  NAND3_X1  g798(.A1(new_n935), .A2(new_n234), .A3(new_n984), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n1000), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1001));
  AOI21_X1  g800(.A(KEYINPUT63), .B1(new_n1000), .B2(G211gat), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n954), .A2(new_n987), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n783), .A2(G211gat), .ZN(new_n1004));
  OAI22_X1  g803(.A1(new_n1001), .A2(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(G1354gat));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n935), .A2(new_n1006), .A3(new_n984), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1006), .B1(new_n935), .B2(new_n984), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n1007), .A2(new_n1008), .A3(new_n284), .ZN(new_n1009));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n718), .A2(new_n1010), .ZN(new_n1011));
  OAI22_X1  g810(.A1(new_n1009), .A2(new_n1010), .B1(new_n1003), .B2(new_n1011), .ZN(G1355gat));
endmodule


