//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G15gat), .ZN(new_n204));
  INV_X1    g003(.A(G15gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT91), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(new_n206), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n202), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(new_n202), .A3(new_n211), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n217));
  OAI21_X1  g016(.A(G29gat), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT88), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT88), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n220), .B(G29gat), .C1(new_n216), .C2(new_n217), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT14), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n219), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(G43gat), .A2(G50gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(G43gat), .A2(G50gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT15), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n219), .A2(new_n221), .A3(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT89), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n229), .A2(new_n230), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(G43gat), .A2(G50gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(G43gat), .A2(G50gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n239), .A2(new_n235), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n224), .A2(new_n226), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n224), .B2(new_n226), .ZN(new_n245));
  OAI22_X1  g044(.A1(new_n238), .A2(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n233), .B1(new_n234), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT17), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT87), .B(G36gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n220), .B1(new_n249), .B2(G29gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n221), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n226), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT90), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n224), .A2(new_n226), .A3(new_n243), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n237), .A3(new_n240), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT89), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n241), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n252), .A2(new_n231), .A3(new_n256), .A4(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT17), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n233), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n215), .B1(new_n248), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G229gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n260), .A2(new_n233), .B1(new_n213), .B2(new_n214), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n264), .B(KEYINPUT13), .Z(new_n268));
  NOR2_X1   g067(.A1(new_n247), .A2(new_n215), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(new_n266), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT93), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n247), .A2(new_n215), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n209), .A2(new_n202), .A3(new_n211), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(new_n212), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n233), .A3(new_n260), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n268), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n267), .A2(KEYINPUT18), .B1(new_n271), .B2(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n254), .A2(new_n255), .B1(new_n258), .B2(new_n241), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n219), .A2(new_n221), .A3(new_n231), .ZN(new_n281));
  AOI221_X4 g080(.A(KEYINPUT17), .B1(new_n228), .B2(new_n232), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n261), .B1(new_n260), .B2(new_n233), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n274), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(new_n264), .A3(new_n272), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT18), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G141gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G197gat), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT11), .B(G169gat), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(KEYINPUT12), .Z(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n279), .B(new_n287), .C1(KEYINPUT92), .C2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n284), .A2(KEYINPUT18), .A3(new_n264), .A4(new_n272), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n277), .B1(new_n276), .B2(new_n268), .ZN(new_n296));
  INV_X1    g095(.A(new_n268), .ZN(new_n297));
  AOI211_X1 g096(.A(KEYINPUT93), .B(new_n297), .C1(new_n272), .C2(new_n275), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n295), .B(KEYINPUT92), .C1(new_n296), .C2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n263), .A2(new_n266), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT18), .B1(new_n301), .B2(new_n264), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n299), .B(new_n292), .C1(new_n300), .C2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G232gat), .A2(G233gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT41), .ZN(new_n306));
  XNOR2_X1  g105(.A(G134gat), .B(G162gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT98), .ZN(new_n310));
  XNOR2_X1  g109(.A(G99gat), .B(G106gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G99gat), .A2(G106gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT8), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G85gat), .B2(G92gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n315));
  OAI211_X1 g114(.A(G85gat), .B(G92gat), .C1(new_n315), .C2(KEYINPUT96), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT97), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT96), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT7), .ZN(new_n319));
  AND2_X1   g118(.A1(G85gat), .A2(G92gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT97), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n315), .A2(KEYINPUT96), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n314), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n317), .A2(new_n322), .A3(KEYINPUT96), .A4(new_n315), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n311), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n321), .B1(new_n319), .B2(new_n320), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n314), .ZN(new_n331));
  AND4_X1   g130(.A1(new_n311), .A2(new_n330), .A3(new_n326), .A4(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n310), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n326), .A3(new_n331), .ZN(new_n334));
  INV_X1    g133(.A(new_n311), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n325), .A2(new_n311), .A3(new_n326), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT98), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n333), .B(new_n338), .C1(new_n282), .C2(new_n283), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n327), .A2(new_n332), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n340), .A2(new_n247), .B1(KEYINPUT41), .B2(new_n305), .ZN(new_n341));
  XNOR2_X1  g140(.A(G190gat), .B(G218gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n342), .B(KEYINPUT99), .Z(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n339), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n344), .B1(new_n339), .B2(new_n341), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n309), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n339), .A2(new_n341), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n343), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n339), .A2(new_n341), .A3(new_n344), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n308), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G120gat), .B(G148gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G176gat), .B(G204gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G64gat), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g157(.A1(G71gat), .A2(G78gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(G71gat), .A2(G78gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT94), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n363), .A3(new_n360), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n358), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n361), .B(KEYINPUT94), .C1(new_n356), .C2(new_n357), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(new_n327), .B2(new_n332), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n336), .A2(new_n337), .A3(new_n367), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n340), .A2(KEYINPUT10), .A3(new_n367), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G230gat), .A2(G233gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n369), .B2(new_n370), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n355), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n375), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n372), .B2(new_n373), .ZN(new_n381));
  INV_X1    g180(.A(new_n355), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n381), .A2(new_n377), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n385));
  INV_X1    g184(.A(G155gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n367), .A2(KEYINPUT21), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n274), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n274), .A2(new_n390), .A3(new_n389), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n393), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n395), .A2(new_n391), .A3(new_n387), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G183gat), .B(G211gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT21), .ZN(new_n400));
  NAND2_X1  g199(.A1(G231gat), .A2(G233gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n368), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(G231gat), .B(G233gat), .C1(new_n367), .C2(KEYINPUT21), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G127gat), .ZN(new_n405));
  INV_X1    g204(.A(G127gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n406), .A3(new_n403), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n399), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n399), .A3(new_n407), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n397), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n405), .A2(new_n399), .A3(new_n407), .ZN(new_n412));
  OAI22_X1  g211(.A1(new_n412), .A2(new_n408), .B1(new_n396), .B2(new_n394), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n352), .A2(new_n384), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  XNOR2_X1  g215(.A(G155gat), .B(G162gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G141gat), .B(G148gat), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(KEYINPUT2), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(G141gat), .B(G148gat), .Z(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT75), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT75), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n417), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT2), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT76), .B(G162gat), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(G155gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n420), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(G211gat), .B(G218gat), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT71), .B(G197gat), .ZN(new_n433));
  INV_X1    g232(.A(G204gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT72), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT22), .ZN(new_n437));
  INV_X1    g236(.A(G211gat), .ZN(new_n438));
  INV_X1    g237(.A(G218gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n436), .B1(new_n435), .B2(new_n440), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n432), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n443), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n431), .A3(new_n441), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT29), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n430), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n449), .B(new_n420), .C1(new_n425), .C2(new_n428), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n444), .A2(new_n446), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G228gat), .ZN(new_n453));
  INV_X1    g252(.A(G233gat), .ZN(new_n454));
  OAI22_X1  g253(.A1(new_n450), .A2(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g255(.A1(new_n450), .A2(new_n453), .A3(new_n454), .A4(new_n452), .ZN(new_n457));
  OAI21_X1  g256(.A(G22gat), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n448), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n429), .ZN(new_n461));
  INV_X1    g260(.A(new_n452), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(G228gat), .A3(G233gat), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n203), .A3(new_n455), .ZN(new_n464));
  XOR2_X1   g263(.A(G78gat), .B(G106gat), .Z(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT31), .B(G50gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n458), .A2(new_n459), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n470), .A2(new_n467), .B1(new_n458), .B2(new_n464), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT80), .ZN(new_n473));
  INV_X1    g272(.A(G113gat), .ZN(new_n474));
  INV_X1    g273(.A(G120gat), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT1), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G127gat), .B(G134gat), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT67), .B(G113gat), .Z(new_n478));
  OAI211_X1 g277(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n475), .ZN(new_n479));
  INV_X1    g278(.A(new_n476), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(G113gat), .B2(G120gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n481), .B2(new_n477), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n429), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n429), .A2(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT77), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n451), .A2(new_n482), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT77), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n429), .A2(new_n488), .A3(KEYINPUT3), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT78), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT78), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n486), .A2(new_n487), .A3(new_n492), .A4(new_n489), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n484), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g294(.A1(G225gat), .A2(G233gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G1gat), .B(G29gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT0), .ZN(new_n499));
  XNOR2_X1  g298(.A(G57gat), .B(G85gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n499), .B(new_n500), .Z(new_n501));
  INV_X1    g300(.A(new_n496), .ZN(new_n502));
  AOI211_X1 g301(.A(new_n502), .B(new_n484), .C1(new_n491), .C2(new_n493), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n429), .B(new_n482), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n502), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n497), .B(new_n501), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n493), .ZN(new_n510));
  INV_X1    g309(.A(new_n484), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n496), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(KEYINPUT5), .A3(new_n505), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n501), .B1(new_n513), .B2(new_n497), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n473), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n501), .ZN(new_n516));
  INV_X1    g315(.A(new_n497), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n506), .B1(new_n494), .B2(new_n496), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT80), .A3(new_n508), .A4(new_n507), .ZN(new_n520));
  AOI211_X1 g319(.A(new_n501), .B(new_n508), .C1(new_n513), .C2(new_n497), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G8gat), .B(G36gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G64gat), .B(G92gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n524), .B(new_n525), .Z(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G183gat), .ZN(new_n528));
  INV_X1    g327(.A(G190gat), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT24), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT24), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(G183gat), .A3(G190gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G183gat), .B2(G190gat), .ZN(new_n534));
  INV_X1    g333(.A(G169gat), .ZN(new_n535));
  INV_X1    g334(.A(G176gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT23), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT23), .B1(new_n535), .B2(new_n536), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT25), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT64), .B(G190gat), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n528), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n533), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(KEYINPUT25), .A3(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT26), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n537), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n540), .ZN(new_n553));
  OAI22_X1  g352(.A1(new_n537), .A2(new_n551), .B1(new_n528), .B2(new_n529), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G183gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT66), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n546), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n546), .B2(new_n556), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n550), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT73), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G226gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n454), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT29), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n550), .A2(KEYINPUT73), .A3(new_n561), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT65), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n545), .A2(new_n570), .A3(new_n549), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n545), .B2(new_n549), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n566), .B(new_n561), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n444), .A2(new_n446), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n561), .B1(new_n571), .B2(new_n572), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n567), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n550), .A2(KEYINPUT73), .A3(new_n561), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT73), .B1(new_n550), .B2(new_n561), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n566), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n580), .B(new_n576), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n575), .B1(new_n574), .B2(new_n577), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n527), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n567), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n581), .A2(new_n582), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n573), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n577), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT74), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n593), .A2(new_n585), .A3(new_n578), .A4(new_n526), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n588), .A2(KEYINPUT30), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n586), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT30), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n596), .A2(new_n597), .A3(new_n593), .A4(new_n526), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n472), .B1(new_n523), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n482), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n579), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G227gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n454), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n482), .B(new_n561), .C1(new_n571), .C2(new_n572), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT32), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT68), .B(G71gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G99gat), .ZN(new_n611));
  XOR2_X1   g410(.A(G15gat), .B(G43gat), .Z(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n606), .B(KEYINPUT32), .C1(new_n608), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n605), .ZN(new_n618));
  INV_X1    g417(.A(new_n604), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n618), .B2(new_n619), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n617), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n614), .A3(new_n616), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT36), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n617), .A2(new_n624), .A3(KEYINPUT70), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n617), .B2(KEYINPUT70), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT36), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n416), .B1(new_n600), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n628), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n626), .B1(new_n635), .B2(KEYINPUT36), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n595), .A2(new_n598), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n519), .A2(new_n508), .A3(new_n507), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n521), .B1(new_n638), .B2(new_n473), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n639), .B2(new_n520), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n636), .B(KEYINPUT82), .C1(new_n640), .C2(new_n472), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n642));
  OR3_X1    g441(.A1(new_n494), .A2(new_n496), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT39), .B1(new_n504), .B2(new_n502), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n644), .A2(KEYINPUT84), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(KEYINPUT84), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n645), .B(new_n646), .C1(new_n494), .C2(new_n496), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n643), .A2(new_n501), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(KEYINPUT85), .B2(KEYINPUT40), .ZN(new_n649));
  NOR2_X1   g448(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n643), .A2(new_n501), .A3(new_n650), .A4(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n513), .A2(KEYINPUT86), .A3(new_n497), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT86), .B1(new_n513), .B2(new_n497), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n516), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n513), .A2(new_n497), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT86), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n501), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n522), .B1(new_n661), .B2(new_n509), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT37), .ZN(new_n663));
  INV_X1    g462(.A(new_n583), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n664), .A2(new_n566), .B1(new_n567), .B2(new_n579), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n665), .B2(new_n577), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n574), .A2(new_n576), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT38), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n596), .A2(new_n593), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n668), .B(new_n527), .C1(new_n669), .C2(KEYINPUT37), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n527), .A2(KEYINPUT37), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n669), .A2(KEYINPUT37), .B1(new_n588), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT38), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n670), .B(new_n594), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n657), .B(new_n472), .C1(new_n662), .C2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n633), .A2(new_n641), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n623), .A2(new_n625), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n599), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n470), .A2(new_n467), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n458), .A2(new_n464), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n468), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n678), .A2(new_n682), .A3(KEYINPUT35), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n662), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n629), .A2(new_n630), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n523), .A2(new_n685), .A3(new_n472), .A4(new_n599), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT35), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n304), .B(new_n415), .C1(new_n676), .C2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n523), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g491(.A(KEYINPUT16), .B(G8gat), .Z(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT101), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(KEYINPUT101), .B2(KEYINPUT42), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n689), .A2(new_n637), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n689), .A2(new_n637), .A3(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n202), .B1(new_n689), .B2(new_n637), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT102), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n696), .B(new_n702), .C1(new_n698), .C2(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(G1325gat));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n205), .A3(new_n677), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n689), .A2(new_n632), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n205), .ZN(G1326gat));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n682), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(KEYINPUT103), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(KEYINPUT103), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT43), .B(G22gat), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n709), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(new_n600), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n675), .A3(new_n636), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n688), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n347), .A2(new_n351), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n352), .B1(new_n676), .B2(new_n688), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(new_n718), .ZN(new_n722));
  INV_X1    g521(.A(new_n384), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n304), .A2(new_n414), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n690), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n222), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n726), .B2(new_n725), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n721), .A2(new_n724), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n222), .A3(new_n690), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT45), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n722), .A2(new_n637), .A3(new_n724), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n249), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n249), .B(new_n599), .C1(new_n735), .C2(KEYINPUT46), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n724), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(KEYINPUT46), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n734), .A2(new_n739), .A3(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1329gat));
  NAND2_X1  g543(.A1(new_n676), .A2(new_n688), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n718), .B1(new_n745), .B2(new_n719), .ZN(new_n746));
  AOI211_X1 g545(.A(KEYINPUT44), .B(new_n352), .C1(new_n716), .C2(new_n688), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n632), .B(new_n724), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n722), .A2(KEYINPUT107), .A3(new_n632), .A4(new_n724), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(G43gat), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(G43gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n729), .A2(new_n753), .A3(new_n677), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n748), .A2(G43gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n754), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(G1330gat));
  OAI211_X1 g560(.A(new_n682), .B(new_n724), .C1(new_n746), .C2(new_n747), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n722), .A2(KEYINPUT109), .A3(new_n682), .A4(new_n724), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(G50gat), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n472), .A2(G50gat), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n745), .A2(new_n719), .A3(new_n724), .A4(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(KEYINPUT48), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n762), .A2(G50gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n768), .B(KEYINPUT108), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n770), .A2(new_n775), .ZN(G1331gat));
  NAND2_X1  g575(.A1(new_n294), .A2(new_n303), .ZN(new_n777));
  INV_X1    g576(.A(new_n414), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n777), .A2(new_n778), .A3(new_n719), .A4(new_n384), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n717), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n690), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G57gat), .ZN(G1332gat));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n717), .A2(new_n779), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n599), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  AND2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(G1333gat));
  INV_X1    g591(.A(G71gat), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n677), .B(KEYINPUT111), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n780), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n784), .A2(new_n632), .A3(new_n786), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(G71gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g597(.A1(new_n787), .A2(new_n472), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g599(.A1(new_n777), .A2(new_n414), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n715), .A2(new_n675), .A3(new_n636), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n662), .A2(new_n683), .B1(new_n686), .B2(KEYINPUT35), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n719), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n717), .A2(KEYINPUT51), .A3(new_n719), .A4(new_n801), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(G85gat), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n808), .A2(new_n809), .A3(new_n690), .A4(new_n723), .ZN(new_n810));
  INV_X1    g609(.A(new_n722), .ZN(new_n811));
  INV_X1    g610(.A(new_n801), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n384), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n811), .A2(new_n523), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n810), .B1(new_n815), .B2(new_n809), .ZN(G1336gat));
  OAI211_X1 g615(.A(new_n637), .B(new_n813), .C1(new_n746), .C2(new_n747), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT113), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n722), .A2(new_n819), .A3(new_n637), .A4(new_n813), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(G92gat), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n599), .A2(G92gat), .A3(new_n384), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(new_n808), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n817), .A2(G92gat), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n826), .A3(new_n807), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n804), .A2(KEYINPUT112), .A3(new_n805), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n822), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n824), .A2(new_n831), .ZN(G1337gat));
  INV_X1    g631(.A(G99gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n677), .A2(new_n833), .A3(new_n723), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT114), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n808), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n811), .A2(new_n636), .A3(new_n814), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n833), .ZN(G1338gat));
  NAND3_X1  g637(.A1(new_n722), .A2(new_n682), .A3(new_n813), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G106gat), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n472), .A2(G106gat), .A3(new_n384), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n827), .A2(new_n828), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT53), .B1(new_n808), .B2(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(G1339gat));
  NAND2_X1  g646(.A1(new_n271), .A2(new_n278), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n287), .A2(new_n848), .A3(new_n295), .A4(new_n293), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n272), .A2(new_n275), .A3(new_n297), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n850), .B(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n264), .B1(new_n284), .B2(new_n272), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n291), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n383), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n372), .A2(new_n380), .A3(new_n373), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n376), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n355), .B1(new_n381), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(KEYINPUT55), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n372), .A2(new_n380), .A3(new_n373), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n381), .A3(new_n859), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n374), .A2(new_n859), .A3(new_n375), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n382), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n862), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n855), .A2(new_n856), .A3(new_n861), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n414), .B1(new_n868), .B2(new_n719), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n861), .A2(new_n856), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n777), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n849), .A2(new_n854), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n352), .B1(new_n872), .B2(new_n384), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n415), .B2(new_n777), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n352), .A2(new_n384), .A3(new_n414), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n304), .A3(KEYINPUT115), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n869), .A2(new_n875), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(new_n682), .A3(new_n635), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n690), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n637), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n478), .A3(new_n777), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n880), .A2(new_n682), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(new_n690), .A3(new_n599), .A4(new_n677), .ZN(new_n886));
  OAI21_X1  g685(.A(G113gat), .B1(new_n886), .B2(new_n304), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(G1340gat));
  NOR3_X1   g687(.A1(new_n886), .A2(new_n475), .A3(new_n384), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n723), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n475), .ZN(G1341gat));
  NAND3_X1  g690(.A1(new_n883), .A2(new_n406), .A3(new_n414), .ZN(new_n892));
  OAI21_X1  g691(.A(G127gat), .B1(new_n886), .B2(new_n778), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1342gat));
  NAND2_X1  g693(.A1(new_n599), .A2(new_n719), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT117), .Z(new_n896));
  OR3_X1    g695(.A1(new_n882), .A2(G134gat), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n886), .B2(new_n352), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G1343gat));
  NOR2_X1   g700(.A1(new_n632), .A2(new_n523), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n869), .A2(new_n875), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n879), .A2(new_n877), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n472), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT121), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n637), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n304), .A2(G141gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT58), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(G141gat), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n880), .A2(new_n912), .A3(new_n472), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT118), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(new_n912), .C1(new_n880), .C2(new_n472), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n599), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(new_n304), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n910), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n913), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n861), .A2(new_n856), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT55), .B1(new_n858), .B2(new_n860), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n922), .A2(new_n923), .A3(new_n872), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n778), .B1(new_n924), .B2(new_n352), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n294), .B2(new_n303), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n873), .B1(new_n870), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n904), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n682), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n915), .B1(new_n929), .B2(new_n912), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT118), .B(KEYINPUT57), .C1(new_n928), .C2(new_n682), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n921), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n918), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(KEYINPUT119), .A3(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n917), .B2(new_n918), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n936), .A3(new_n777), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(G141gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n937), .B2(G141gat), .ZN(new_n940));
  NOR4_X1   g739(.A1(new_n906), .A2(G141gat), .A3(new_n637), .A4(new_n304), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT58), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n920), .B1(new_n942), .B2(new_n943), .ZN(G1344gat));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n945));
  AOI211_X1 g744(.A(new_n945), .B(G148gat), .C1(new_n908), .C2(new_n723), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n934), .A2(new_n936), .A3(new_n945), .A4(new_n723), .ZN(new_n947));
  INV_X1    g746(.A(G148gat), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n869), .A2(new_n875), .B1(new_n304), .B2(new_n878), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n912), .B1(new_n949), .B2(new_n472), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n921), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n723), .A3(new_n933), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n952), .B2(KEYINPUT59), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n946), .B1(new_n947), .B2(new_n953), .ZN(G1345gat));
  NAND2_X1  g753(.A1(new_n934), .A2(new_n936), .ZN(new_n955));
  OAI21_X1  g754(.A(G155gat), .B1(new_n955), .B2(new_n778), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n908), .A2(new_n386), .A3(new_n414), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1346gat));
  OAI21_X1  g757(.A(new_n427), .B1(new_n955), .B2(new_n352), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n896), .A2(new_n427), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n907), .B2(new_n960), .ZN(G1347gat));
  NAND2_X1  g760(.A1(new_n523), .A2(new_n637), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(new_n794), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n885), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n965), .A2(new_n535), .A3(new_n304), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n881), .A2(new_n963), .ZN(new_n967));
  AOI21_X1  g766(.A(G169gat), .B1(new_n967), .B2(new_n777), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n966), .A2(new_n968), .ZN(G1348gat));
  INV_X1    g768(.A(new_n965), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(G176gat), .A3(new_n723), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(KEYINPUT122), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(KEYINPUT122), .ZN(new_n973));
  AOI21_X1  g772(.A(G176gat), .B1(new_n967), .B2(new_n723), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(G1349gat));
  OAI21_X1  g774(.A(G183gat), .B1(new_n965), .B2(new_n778), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n967), .A2(new_n556), .A3(new_n414), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(KEYINPUT123), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g778(.A1(new_n967), .A2(new_n546), .A3(new_n719), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n970), .A2(new_n719), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(G190gat), .ZN(new_n983));
  AOI211_X1 g782(.A(KEYINPUT61), .B(new_n529), .C1(new_n970), .C2(new_n719), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(G1351gat));
  NOR2_X1   g784(.A1(new_n632), .A2(new_n962), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n987), .B1(new_n921), .B2(new_n950), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n988), .A2(new_n777), .ZN(new_n989));
  OR2_X1    g788(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n990), .A2(G197gat), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n987), .A2(new_n929), .ZN(new_n993));
  INV_X1    g792(.A(G197gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n993), .A2(new_n994), .A3(new_n777), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n992), .A2(new_n995), .ZN(G1352gat));
  NAND3_X1  g795(.A1(new_n993), .A2(new_n434), .A3(new_n723), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n997), .B(KEYINPUT62), .Z(new_n998));
  AND2_X1   g797(.A1(new_n988), .A2(new_n723), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n999), .B2(new_n434), .ZN(G1353gat));
  NAND3_X1  g799(.A1(new_n993), .A2(new_n438), .A3(new_n414), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n988), .A2(new_n414), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT63), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1003), .A2(KEYINPUT125), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n438), .B1(KEYINPUT125), .B2(new_n1003), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1004), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n439), .A3(new_n719), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n988), .A2(new_n719), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1009), .B1(new_n1010), .B2(new_n439), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1011), .B(KEYINPUT126), .ZN(G1355gat));
endmodule


