//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(G1gat), .ZN(new_n209));
  AOI21_X1  g008(.A(G8gat), .B1(new_n209), .B2(KEYINPUT86), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(new_n211), .B2(G1gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n209), .B(new_n212), .C1(KEYINPUT86), .C2(G8gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(KEYINPUT84), .B(G50gat), .Z(new_n218));
  INV_X1    g017(.A(G43gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT83), .B(G43gat), .ZN(new_n221));
  INV_X1    g020(.A(G50gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT15), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT15), .ZN(new_n226));
  NAND2_X1  g025(.A1(G29gat), .A2(G36gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  NOR3_X1   g027(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(KEYINPUT85), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n229), .A2(KEYINPUT85), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n226), .B(new_n227), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OR3_X1    g031(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n233), .A2(new_n228), .B1(G29gat), .B2(G36gat), .ZN(new_n234));
  OAI22_X1  g033(.A1(new_n224), .A2(new_n232), .B1(new_n234), .B2(new_n226), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n235), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n216), .A2(KEYINPUT87), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT87), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n240), .A3(new_n215), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n207), .B(new_n236), .C1(new_n238), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT89), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n206), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n235), .B(KEYINPUT17), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(new_n239), .A3(new_n241), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n249), .A2(KEYINPUT18), .A3(new_n207), .A4(new_n236), .ZN(new_n250));
  INV_X1    g049(.A(new_n235), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT88), .B1(new_n251), .B2(new_n216), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n236), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n207), .B(KEYINPUT13), .Z(new_n254));
  NAND3_X1  g053(.A1(new_n217), .A2(KEYINPUT88), .A3(new_n235), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n245), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n247), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n247), .A2(new_n257), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G120gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  XNOR2_X1  g061(.A(G127gat), .B(G134gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n263), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(KEYINPUT1), .B2(new_n261), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  INV_X1    g067(.A(G169gat), .ZN(new_n269));
  INV_X1    g068(.A(G176gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT26), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(new_n269), .A3(new_n270), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n268), .B(new_n272), .C1(new_n276), .C2(KEYINPUT26), .ZN(new_n277));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n284), .B(KEYINPUT28), .Z(new_n285));
  NAND3_X1  g084(.A1(new_n277), .A2(KEYINPUT68), .A3(new_n278), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n268), .A2(KEYINPUT23), .ZN(new_n289));
  MUX2_X1   g088(.A(KEYINPUT23), .B(new_n289), .S(new_n271), .Z(new_n290));
  OAI21_X1  g089(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n278), .ZN(new_n292));
  NAND3_X1  g091(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n288), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n288), .B1(new_n289), .B2(new_n271), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n274), .A2(KEYINPUT23), .A3(new_n275), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n292), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT66), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(new_n305), .A3(new_n292), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n298), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n295), .B1(new_n307), .B2(KEYINPUT67), .ZN(new_n308));
  INV_X1    g107(.A(new_n298), .ZN(new_n309));
  AOI221_X4 g108(.A(KEYINPUT66), .B1(new_n291), .B2(new_n278), .C1(new_n300), .C2(new_n301), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(new_n302), .B2(new_n292), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n309), .B(KEYINPUT67), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n267), .B(new_n287), .C1(new_n308), .C2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(new_n312), .A3(new_n295), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n320), .A2(KEYINPUT69), .A3(new_n267), .A4(new_n287), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n287), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n264), .A2(new_n266), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n316), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT33), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT32), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n325), .B2(new_n327), .ZN(new_n330));
  XNOR2_X1  g129(.A(G15gat), .B(G43gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G71gat), .B(G99gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n328), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n325), .A2(new_n327), .ZN(new_n335));
  INV_X1    g134(.A(new_n333), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT33), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(KEYINPUT32), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n316), .A2(new_n324), .A3(new_n326), .A4(new_n321), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT34), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n339), .A2(KEYINPUT34), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT70), .B1(new_n334), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n328), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n335), .A2(KEYINPUT32), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n336), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT34), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n339), .B(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .A4(new_n338), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n353));
  XOR2_X1   g152(.A(G141gat), .B(G148gat), .Z(new_n354));
  INV_X1    g153(.A(G155gat), .ZN(new_n355));
  INV_X1    g154(.A(G162gat), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT2), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G155gat), .B(G162gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n359), .A3(new_n357), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(new_n323), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n353), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n361), .A2(new_n362), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n267), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT4), .B1(new_n363), .B2(new_n323), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n363), .A2(KEYINPUT3), .B1(new_n264), .B2(new_n266), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n361), .A2(new_n375), .A3(new_n362), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT76), .B(KEYINPUT4), .C1(new_n363), .C2(new_n323), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n365), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n367), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT5), .B1(new_n370), .B2(new_n371), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n366), .B1(new_n374), .B2(new_n376), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G1gat), .B(G29gat), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT78), .ZN(new_n386));
  XOR2_X1   g185(.A(G57gat), .B(G85gat), .Z(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT79), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n386), .B(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n389), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n352), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n384), .A2(new_n393), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n382), .B(new_n378), .C1(new_n372), .C2(KEYINPUT76), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n398), .A2(new_n367), .B1(new_n382), .B2(new_n381), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT6), .B1(new_n399), .B2(new_n392), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT80), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n384), .A2(KEYINPUT6), .A3(new_n393), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n407), .B(KEYINPUT75), .Z(new_n408));
  NAND3_X1  g207(.A1(new_n320), .A2(new_n408), .A3(new_n287), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(G211gat), .A2(G218gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G211gat), .A2(G218gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(KEYINPUT72), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT72), .ZN(new_n415));
  INV_X1    g214(.A(new_n413), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(new_n411), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n416), .A2(KEYINPUT22), .ZN(new_n420));
  INV_X1    g219(.A(G197gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT71), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT71), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G197gat), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n422), .A2(new_n424), .A3(G204gat), .ZN(new_n425));
  AOI21_X1  g224(.A(G204gat), .B1(new_n422), .B2(new_n424), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n420), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT73), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n416), .A2(new_n411), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT73), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n422), .A2(new_n424), .ZN(new_n432));
  INV_X1    g231(.A(G204gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n422), .A2(new_n424), .A3(G204gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n418), .B1(new_n436), .B2(new_n420), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n429), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT74), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(new_n429), .C1(new_n431), .C2(new_n437), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n408), .A2(KEYINPUT29), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n320), .B2(new_n287), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n410), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n438), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n322), .A2(new_n443), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(new_n409), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n406), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n438), .B1(new_n410), .B2(new_n445), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n439), .A2(new_n441), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n452), .A3(new_n409), .ZN(new_n453));
  INV_X1    g252(.A(new_n406), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(KEYINPUT30), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n457), .B(new_n406), .C1(new_n446), .C2(new_n449), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n402), .A2(new_n403), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n349), .B1(new_n346), .B2(new_n338), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT81), .Z(new_n463));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n376), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n439), .A2(new_n441), .A3(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n464), .B(new_n429), .C1(new_n431), .C2(new_n437), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n375), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n363), .ZN(new_n469));
  INV_X1    g268(.A(G228gat), .ZN(new_n470));
  INV_X1    g269(.A(G233gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G22gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n430), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n436), .A2(new_n420), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n436), .B2(new_n420), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n368), .B1(new_n479), .B2(new_n375), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n438), .A2(new_n465), .ZN(new_n481));
  OAI22_X1  g280(.A1(new_n480), .A2(new_n481), .B1(new_n470), .B2(new_n471), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n473), .A2(new_n474), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n474), .B1(new_n473), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n463), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n473), .A2(new_n482), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G22gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n463), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n474), .A3(new_n482), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G50gat), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n485), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n485), .B2(new_n490), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n351), .A2(new_n459), .A3(new_n461), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n460), .A2(new_n492), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n400), .A2(new_n397), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n456), .A2(new_n458), .B1(new_n498), .B2(new_n403), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT35), .B1(new_n499), .B2(new_n500), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n497), .A2(new_n501), .A3(new_n351), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n351), .A2(new_n461), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT36), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n399), .A2(new_n392), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n450), .B(new_n403), .C1(new_n394), .C2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n446), .B2(new_n449), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n442), .B1(new_n410), .B2(new_n445), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n448), .A2(new_n447), .A3(new_n409), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT37), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n454), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT38), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n451), .A2(new_n453), .A3(KEYINPUT37), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n510), .A2(KEYINPUT38), .A3(new_n517), .A4(new_n454), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n508), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n456), .A2(new_n458), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT40), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n365), .B1(new_n372), .B2(new_n377), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n392), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT39), .B1(new_n364), .B2(new_n366), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n521), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n522), .A2(new_n526), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(KEYINPUT40), .A3(new_n392), .A4(new_n524), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n397), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n494), .B1(new_n519), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n402), .A2(new_n403), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n534), .B(new_n520), .C1(new_n492), .C2(new_n493), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n351), .A2(new_n537), .A3(new_n461), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n506), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n260), .B1(new_n504), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT98), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT97), .ZN(new_n542));
  INV_X1    g341(.A(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n542), .B(KEYINPUT7), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT7), .ZN(new_n546));
  OAI211_X1 g345(.A(G85gat), .B(G92gat), .C1(new_n546), .C2(KEYINPUT97), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n543), .B2(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G99gat), .B(G106gat), .Z(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n548), .B2(new_n550), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n541), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n552), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n548), .A3(new_n550), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT98), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n235), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n560), .A2(KEYINPUT99), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT99), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(new_n559), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n562), .A2(new_n563), .B1(new_n238), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT101), .ZN(new_n567));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n566), .A2(new_n568), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT96), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n571), .B(new_n572), .C1(KEYINPUT100), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n566), .A2(new_n568), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT101), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n572), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(KEYINPUT100), .A3(new_n581), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n576), .ZN(new_n584));
  OR2_X1    g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT9), .B1(new_n589), .B2(KEYINPUT90), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT90), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n587), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT9), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n586), .B1(new_n585), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT91), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n589), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n593), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G127gat), .B(G155gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT21), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n216), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n604), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT94), .ZN(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT93), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT95), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n607), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n578), .A2(new_n584), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT102), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n578), .A2(new_n584), .A3(new_n619), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n557), .A2(new_n558), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n557), .A2(KEYINPUT103), .A3(new_n558), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n600), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n597), .A2(new_n599), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n628), .A2(new_n623), .A3(new_n624), .A4(new_n593), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT10), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n564), .A2(new_n631), .A3(new_n600), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n622), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n622), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n627), .A2(new_n634), .A3(new_n629), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n636), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n621), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n540), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n534), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(G1gat), .Z(G1324gat));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645));
  INV_X1    g444(.A(new_n520), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n540), .A2(new_n646), .A3(new_n641), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(G8gat), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  NAND4_X1  g448(.A1(new_n540), .A2(new_n646), .A3(new_n641), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n645), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n648), .B2(new_n650), .ZN(new_n656));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT104), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n658), .ZN(G1325gat));
  AOI211_X1 g458(.A(KEYINPUT36), .B(new_n460), .C1(new_n343), .C2(new_n350), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n537), .B1(new_n351), .B2(new_n461), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n642), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n505), .A2(G15gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(new_n642), .B2(new_n664), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n642), .A2(new_n494), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT43), .B(G22gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  NAND2_X1  g467(.A1(new_n578), .A2(new_n584), .ZN(new_n669));
  INV_X1    g468(.A(new_n616), .ZN(new_n670));
  INV_X1    g469(.A(new_n640), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT105), .Z(new_n673));
  AND2_X1   g472(.A1(new_n540), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(G29gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n534), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  NOR2_X1   g477(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n662), .A2(new_n536), .B1(new_n496), .B2(new_n503), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n578), .A2(new_n584), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n504), .A2(new_n539), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n669), .A3(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n260), .A2(new_n616), .A3(new_n640), .ZN(new_n686));
  AND4_X1   g485(.A1(new_n676), .A2(new_n682), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n678), .B1(new_n675), .B2(new_n687), .ZN(G1328gat));
  INV_X1    g487(.A(G36gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n689), .A3(new_n646), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT46), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT46), .ZN(new_n692));
  AND4_X1   g491(.A1(new_n646), .A2(new_n682), .A3(new_n685), .A4(new_n686), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n691), .B(new_n692), .C1(new_n689), .C2(new_n693), .ZN(G1329gat));
  NOR2_X1   g493(.A1(new_n505), .A2(new_n221), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n540), .A2(new_n673), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT107), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n662), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n682), .A2(new_n699), .A3(new_n685), .A4(new_n686), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n221), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n701), .A3(KEYINPUT47), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  INV_X1    g502(.A(new_n701), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n697), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(G1330gat));
  INV_X1    g505(.A(new_n494), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n674), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n218), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n494), .A2(new_n709), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n682), .A2(new_n685), .A3(new_n686), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT48), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(new_n715), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1331gat));
  INV_X1    g516(.A(new_n260), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n621), .A2(new_n718), .A3(new_n671), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n683), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n534), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(G57gat), .Z(G1332gat));
  NAND2_X1  g521(.A1(new_n720), .A2(KEYINPUT108), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n683), .A2(new_n724), .A3(new_n719), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n646), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT49), .B(G64gat), .Z(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(G1333gat));
  NOR3_X1   g529(.A1(new_n720), .A2(G71gat), .A3(new_n505), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n723), .A2(new_n699), .A3(new_n725), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(G71gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n726), .A2(new_n707), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g535(.A(new_n681), .B1(new_n504), .B2(new_n539), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n718), .A2(new_n616), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT51), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n683), .A2(KEYINPUT51), .A3(new_n669), .A4(new_n738), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n737), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n738), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n676), .A2(new_n543), .A3(new_n640), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n718), .A2(new_n616), .A3(new_n671), .ZN(new_n746));
  AND4_X1   g545(.A1(new_n676), .A2(new_n682), .A3(new_n685), .A4(new_n746), .ZN(new_n747));
  OAI22_X1  g546(.A1(new_n744), .A2(new_n745), .B1(new_n747), .B2(new_n543), .ZN(G1336gat));
  NAND4_X1  g547(.A1(new_n682), .A2(new_n646), .A3(new_n685), .A4(new_n746), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G92gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n737), .B2(new_n738), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n742), .B2(new_n743), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n520), .A2(new_n671), .A3(G92gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT110), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT52), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n758));
  OAI211_X1 g557(.A(new_n750), .B(new_n758), .C1(new_n744), .C2(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1337gat));
  XOR2_X1   g559(.A(KEYINPUT113), .B(G99gat), .Z(new_n761));
  NAND4_X1  g560(.A1(new_n351), .A2(new_n461), .A3(new_n640), .A4(new_n761), .ZN(new_n762));
  AND4_X1   g561(.A1(new_n699), .A2(new_n682), .A3(new_n685), .A4(new_n746), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n744), .A2(new_n762), .B1(new_n763), .B2(new_n761), .ZN(G1338gat));
  NAND4_X1  g563(.A1(new_n682), .A2(new_n707), .A3(new_n685), .A4(new_n746), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G106gat), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n494), .A2(G106gat), .A3(new_n671), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT114), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT115), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n753), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT53), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n772));
  OAI211_X1 g571(.A(new_n766), .B(new_n772), .C1(new_n744), .C2(new_n768), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1339gat));
  NAND4_X1  g573(.A1(new_n618), .A2(new_n260), .A3(new_n620), .A4(new_n671), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n627), .A2(new_n629), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n631), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n564), .A2(new_n631), .A3(new_n600), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n634), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n780), .A2(KEYINPUT54), .A3(new_n633), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n782), .B(new_n622), .C1(new_n630), .C2(new_n632), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n639), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n776), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n636), .A2(new_n639), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n783), .A2(new_n639), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n780), .A2(KEYINPUT54), .A3(new_n633), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n785), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n245), .A2(new_n250), .A3(new_n206), .A4(new_n256), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n207), .B1(new_n249), .B2(new_n236), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n254), .B1(new_n253), .B2(new_n255), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n205), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n260), .A2(new_n790), .B1(new_n671), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n790), .B1(new_n578), .B2(new_n584), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n791), .A2(new_n794), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n681), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n775), .B1(new_n799), .B2(new_n616), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n497), .A2(new_n351), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n534), .A2(new_n646), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT117), .ZN(new_n804));
  OAI21_X1  g603(.A(G113gat), .B1(new_n804), .B2(new_n260), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n800), .A2(new_n801), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n260), .A2(G113gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT118), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT119), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n805), .A2(new_n812), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1340gat));
  OAI21_X1  g613(.A(G120gat), .B1(new_n804), .B2(new_n671), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n671), .A2(G120gat), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT120), .Z(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n803), .B2(new_n817), .ZN(G1341gat));
  OAI21_X1  g617(.A(G127gat), .B1(new_n804), .B2(new_n670), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n803), .A2(G127gat), .A3(new_n670), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(KEYINPUT121), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1342gat));
  NOR3_X1   g624(.A1(new_n803), .A2(G134gat), .A3(new_n681), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT56), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n804), .B2(new_n681), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1343gat));
  AND2_X1   g628(.A1(new_n662), .A2(new_n802), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n494), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT122), .B1(new_n798), .B2(new_n640), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n789), .A2(new_n786), .ZN(new_n835));
  INV_X1    g634(.A(new_n259), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n247), .A2(new_n257), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n787), .B2(new_n788), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT123), .B(KEYINPUT55), .C1(new_n787), .C2(new_n788), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n834), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n798), .A2(KEYINPUT122), .A3(new_n640), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n669), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n797), .A2(new_n798), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n670), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n833), .B1(new_n849), .B2(new_n775), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n800), .B2(new_n707), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n718), .B(new_n830), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853));
  INV_X1    g652(.A(new_n775), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n796), .A2(new_n681), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n616), .B1(new_n855), .B2(new_n847), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n853), .B(new_n676), .C1(new_n854), .C2(new_n856), .ZN(new_n857));
  NOR4_X1   g656(.A1(new_n660), .A2(new_n661), .A3(new_n646), .A4(new_n494), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n853), .B1(new_n800), .B2(new_n676), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n260), .A2(G141gat), .ZN(new_n862));
  AOI22_X1  g661(.A1(G141gat), .A2(new_n852), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n852), .B2(G141gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n863), .A2(new_n865), .A3(KEYINPUT58), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n852), .A2(G141gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(new_n862), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n867), .B(new_n868), .C1(KEYINPUT125), .C2(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n866), .A2(new_n870), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n671), .A2(KEYINPUT59), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n830), .B(new_n872), .C1(new_n850), .C2(new_n851), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n830), .A2(new_n640), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n875), .B1(new_n671), .B2(new_n795), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n786), .B(new_n789), .C1(new_n258), .C2(new_n259), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n785), .A2(KEYINPUT123), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n839), .A2(new_n840), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n845), .B(new_n876), .C1(new_n877), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n681), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883));
  INV_X1    g682(.A(new_n790), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n669), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n798), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n797), .A2(new_n883), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n854), .B1(new_n888), .B2(new_n670), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n831), .B1(new_n889), .B2(new_n494), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n800), .A2(new_n832), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n874), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n873), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n860), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n895), .A2(new_n640), .A3(new_n857), .A4(new_n858), .ZN(new_n896));
  AOI21_X1  g695(.A(G148gat), .B1(new_n896), .B2(KEYINPUT59), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT127), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(KEYINPUT59), .ZN(new_n899));
  INV_X1    g698(.A(G148gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n891), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n795), .B1(new_n797), .B2(new_n883), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT126), .B1(new_n681), .B2(new_n790), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n616), .B1(new_n905), .B2(new_n882), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n707), .B1(new_n906), .B2(new_n854), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n902), .B1(new_n907), .B2(new_n831), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT59), .B(G148gat), .C1(new_n908), .C2(new_n874), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n901), .A2(new_n909), .A3(new_n910), .A4(new_n873), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n898), .A2(new_n911), .ZN(G1345gat));
  OAI21_X1  g711(.A(new_n830), .B1(new_n850), .B2(new_n851), .ZN(new_n913));
  OAI21_X1  g712(.A(G155gat), .B1(new_n913), .B2(new_n670), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n861), .A2(new_n355), .A3(new_n616), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1346gat));
  NOR3_X1   g715(.A1(new_n913), .A2(new_n356), .A3(new_n681), .ZN(new_n917));
  AOI21_X1  g716(.A(G162gat), .B1(new_n861), .B2(new_n669), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n676), .A2(new_n520), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n806), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n260), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(new_n269), .ZN(G1348gat));
  NOR2_X1   g722(.A1(new_n921), .A2(new_n671), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(new_n270), .ZN(G1349gat));
  INV_X1    g724(.A(G183gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n921), .B2(new_n670), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n806), .A2(new_n616), .A3(new_n920), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n282), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(G1350gat));
  OAI22_X1  g730(.A1(new_n921), .A2(new_n681), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n932), .B(new_n933), .ZN(G1351gat));
  INV_X1    g733(.A(new_n920), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n935), .A2(new_n660), .A3(new_n661), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(new_n800), .A3(new_n707), .ZN(new_n937));
  AOI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n718), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n908), .A2(new_n699), .A3(new_n935), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n260), .A2(new_n421), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(G1352gat));
  NAND3_X1  g740(.A1(new_n937), .A2(new_n433), .A3(new_n640), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT62), .Z(new_n943));
  AND2_X1   g742(.A1(new_n939), .A2(new_n640), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n433), .ZN(G1353gat));
  INV_X1    g744(.A(G211gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n937), .A2(new_n946), .A3(new_n616), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n890), .A2(new_n891), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n616), .A3(new_n936), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  INV_X1    g751(.A(G218gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n953), .A3(new_n669), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n939), .A2(new_n669), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n953), .ZN(G1355gat));
endmodule


