//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202));
  XOR2_X1   g001(.A(G134gat), .B(G162gat), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT99), .ZN(new_n206));
  INV_X1    g005(.A(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G43gat), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G50gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT15), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT88), .ZN(new_n213));
  OR3_X1    g012(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(KEYINPUT88), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n212), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n220), .A2(new_n211), .A3(new_n217), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n209), .A2(G50gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT15), .B1(new_n222), .B2(KEYINPUT89), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT89), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n210), .A3(new_n224), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n223), .A2(KEYINPUT90), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT90), .B1(new_n223), .B2(new_n225), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT7), .ZN(new_n230));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231));
  INV_X1    g030(.A(G85gat), .ZN(new_n232));
  INV_X1    g031(.A(G92gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(KEYINPUT8), .A2(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT98), .ZN(new_n235));
  XNOR2_X1  g034(.A(G99gat), .B(G106gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n230), .B(new_n234), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n235), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n236), .A2(new_n235), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n241), .A2(new_n238), .A3(new_n230), .A4(new_n234), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n219), .A2(new_n228), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n206), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n242), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n220), .A2(new_n211), .A3(new_n217), .ZN(new_n248));
  INV_X1    g047(.A(new_n227), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n223), .A2(KEYINPUT90), .A3(new_n225), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n247), .B1(new_n251), .B2(new_n218), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(KEYINPUT99), .A3(new_n244), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n219), .A2(new_n228), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT17), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n219), .A2(new_n228), .A3(KEYINPUT17), .ZN(new_n258));
  INV_X1    g057(.A(new_n247), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(KEYINPUT100), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT100), .B1(new_n254), .B2(new_n260), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n205), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n254), .A2(new_n260), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT100), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(G190gat), .A3(new_n261), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(G218gat), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT97), .ZN(new_n270));
  AOI21_X1  g069(.A(G218gat), .B1(new_n264), .B2(new_n268), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT101), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n264), .A2(new_n268), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT101), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n277), .A2(KEYINPUT97), .A3(new_n278), .A4(new_n269), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n272), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n274), .B1(new_n272), .B2(new_n279), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n204), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n272), .A2(new_n279), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n273), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n272), .A2(new_n274), .A3(new_n279), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n203), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n288));
  INV_X1    g087(.A(G57gat), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n289), .A2(G64gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(G64gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G71gat), .ZN(new_n293));
  INV_X1    g092(.A(G78gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(G71gat), .A2(G78gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT94), .ZN(new_n297));
  OAI22_X1  g096(.A1(new_n295), .A2(new_n296), .B1(new_n288), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n292), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT95), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT21), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G127gat), .B(G155gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305));
  INV_X1    g104(.A(G1gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT16), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G1gat), .B2(new_n305), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(G8gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(new_n300), .B2(new_n301), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n304), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G231gat), .A2(G233gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT96), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G183gat), .B(G211gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n313), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n202), .B1(new_n287), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n282), .A2(new_n286), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT102), .A3(new_n320), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G230gat), .A2(G233gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n259), .A2(new_n299), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(new_n300), .B2(new_n247), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OR3_X1    g130(.A1(new_n300), .A2(new_n330), .A3(new_n259), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT103), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n327), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n334), .B2(new_n333), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n329), .A2(new_n326), .ZN(new_n337));
  XOR2_X1   g136(.A(G120gat), .B(G148gat), .Z(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT104), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT105), .ZN(new_n340));
  XNOR2_X1  g139(.A(G176gat), .B(G204gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n333), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(new_n327), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n342), .B1(new_n346), .B2(new_n337), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n325), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT31), .B(G50gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G141gat), .ZN(new_n353));
  INV_X1    g152(.A(G148gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358));
  INV_X1    g157(.A(G155gat), .ZN(new_n359));
  INV_X1    g158(.A(G162gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT2), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(KEYINPUT78), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n357), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(KEYINPUT2), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT78), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n358), .ZN(new_n368));
  NOR3_X1   g167(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n364), .A2(new_n355), .A3(new_n356), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G197gat), .B(G204gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT73), .B(G218gat), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n375), .A2(G211gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n376), .B2(KEYINPUT22), .ZN(new_n377));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n374), .B(new_n378), .C1(new_n376), .C2(KEYINPUT22), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n373), .B1(new_n382), .B2(KEYINPUT3), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n381), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n363), .A2(new_n365), .B1(new_n370), .B2(new_n371), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n385), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G22gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n395), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n383), .B(new_n393), .C1(new_n384), .C2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n396), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n396), .B2(new_n399), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n352), .B(new_n400), .C1(new_n401), .C2(KEYINPUT82), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n401), .A2(KEYINPUT82), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n352), .B(KEYINPUT80), .Z(new_n405));
  INV_X1    g204(.A(new_n400), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n401), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(G8gat), .B(G36gat), .Z(new_n410));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT28), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT27), .ZN(new_n415));
  INV_X1    g214(.A(G183gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT67), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(KEYINPUT67), .A3(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n423), .B2(new_n205), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT64), .B(G183gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n417), .B1(new_n425), .B2(new_n415), .ZN(new_n426));
  NOR2_X1   g225(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429));
  INV_X1    g228(.A(G169gat), .ZN(new_n430));
  INV_X1    g229(.A(G176gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT26), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT26), .B1(new_n430), .B2(new_n431), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n424), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n429), .A2(KEYINPUT24), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT24), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(G183gat), .A3(G190gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(G183gat), .B2(G190gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT23), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT23), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(G169gat), .B2(G176gat), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n445), .A2(new_n447), .A3(new_n435), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT25), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n416), .A2(KEYINPUT64), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT64), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(G183gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n452), .A3(new_n205), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n443), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT65), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n443), .A3(KEYINPUT65), .ZN(new_n457));
  AND4_X1   g256(.A1(KEYINPUT25), .A2(new_n445), .A3(new_n447), .A4(new_n435), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT66), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n449), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT66), .A4(new_n458), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n439), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n413), .B1(new_n463), .B2(KEYINPUT29), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n425), .A2(new_n205), .B1(new_n440), .B2(new_n442), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n458), .B1(new_n465), .B2(KEYINPUT65), .ZN(new_n466));
  INV_X1    g265(.A(new_n457), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n449), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n439), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n413), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n464), .A2(new_n474), .A3(new_n386), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n464), .A2(KEYINPUT75), .A3(new_n474), .A4(new_n386), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT74), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n464), .B2(new_n474), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n391), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT74), .B1(new_n482), .B2(new_n413), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n387), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n412), .B1(new_n485), .B2(KEYINPUT37), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n464), .A2(new_n480), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n413), .B1(new_n470), .B2(new_n471), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n482), .B2(new_n413), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n490), .B2(new_n480), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n491), .A2(new_n387), .B1(new_n477), .B2(new_n478), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND4_X1   g293(.A1(new_n487), .A2(new_n479), .A3(new_n493), .A4(new_n484), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n486), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT38), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT5), .ZN(new_n498));
  INV_X1    g297(.A(G113gat), .ZN(new_n499));
  INV_X1    g298(.A(G120gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G113gat), .A2(G120gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT1), .B1(new_n503), .B2(KEYINPUT69), .ZN(new_n504));
  XNOR2_X1  g303(.A(G127gat), .B(G134gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT69), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n504), .B1(new_n507), .B2(new_n503), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT1), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n501), .A2(new_n510), .A3(new_n502), .ZN(new_n511));
  INV_X1    g310(.A(G134gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G127gat), .ZN(new_n513));
  INV_X1    g312(.A(G127gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G134gat), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT68), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n509), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n373), .A2(new_n508), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n508), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n388), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT79), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n498), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n525));
  INV_X1    g324(.A(new_n519), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n390), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT4), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n519), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n523), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n524), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n527), .A2(new_n529), .A3(new_n532), .A4(new_n530), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(new_n498), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT84), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G1gat), .B(G29gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT0), .ZN(new_n538));
  XNOR2_X1  g337(.A(G57gat), .B(G85gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n538), .B(new_n539), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n524), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n534), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n531), .A2(KEYINPUT5), .A3(new_n532), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT84), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n544), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT6), .B1(new_n548), .B2(new_n540), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n544), .A2(new_n543), .A3(KEYINPUT6), .A4(new_n541), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n479), .A2(new_n484), .A3(new_n412), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n492), .A2(new_n487), .A3(new_n493), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n479), .A2(new_n493), .A3(new_n484), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT86), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n491), .A2(new_n386), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n493), .B1(new_n490), .B2(new_n387), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT38), .B(new_n412), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n553), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n409), .B1(new_n497), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n479), .A2(new_n484), .A3(KEYINPUT30), .A4(new_n412), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n492), .B2(new_n412), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n552), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT76), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT76), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n564), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT85), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n521), .A2(new_n523), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT83), .Z(new_n573));
  OR2_X1    g372(.A1(new_n531), .A2(new_n532), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT39), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n574), .A2(KEYINPUT39), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n540), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT40), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT40), .A4(new_n540), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n547), .A3(new_n580), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n570), .A2(new_n571), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n412), .B1(new_n479), .B2(new_n484), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n479), .A2(new_n484), .A3(new_n412), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(KEYINPUT30), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n552), .A2(new_n568), .A3(new_n565), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n568), .B1(new_n552), .B2(new_n565), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n579), .A2(new_n547), .A3(new_n580), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT85), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n562), .B1(new_n582), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n472), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n463), .A2(KEYINPUT70), .A3(new_n526), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n594), .A2(new_n595), .A3(G227gat), .A4(G233gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT32), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G15gat), .B(G43gat), .Z(new_n600));
  XNOR2_X1  g399(.A(G71gat), .B(G99gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n596), .B(KEYINPUT32), .C1(new_n598), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n594), .A2(new_n595), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n608));
  NAND2_X1  g407(.A1(G227gat), .A2(G233gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT71), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT71), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n607), .A2(new_n612), .A3(new_n608), .A4(new_n609), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n609), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT34), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n606), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n608), .B1(new_n607), .B2(new_n609), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(KEYINPUT71), .B2(new_n610), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n619), .A2(new_n603), .A3(new_n605), .A4(new_n613), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT72), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OR3_X1    g421(.A1(new_n606), .A2(new_n616), .A3(new_n621), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n617), .A2(new_n620), .A3(KEYINPUT36), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n549), .B1(new_n540), .B2(new_n548), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n551), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n585), .B(new_n629), .C1(new_n586), .C2(new_n587), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n409), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n408), .A2(new_n620), .A3(new_n617), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT35), .B1(new_n633), .B2(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n622), .A2(new_n623), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT35), .B1(new_n550), .B2(new_n551), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n635), .A2(new_n570), .A3(new_n408), .A4(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n591), .A2(new_n632), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G169gat), .B(G197gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n255), .A2(new_n310), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT91), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n255), .A2(new_n310), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT13), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT18), .ZN(new_n652));
  INV_X1    g451(.A(new_n646), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n257), .A2(new_n311), .A3(new_n258), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n651), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n652), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n644), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT92), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n644), .B1(new_n657), .B2(KEYINPUT93), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT93), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n656), .B1(new_n664), .B2(new_n658), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n661), .A2(new_n662), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n638), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n349), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n629), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n306), .ZN(G1324gat));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n570), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(G8gat), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  MUX2_X1   g474(.A(new_n673), .B(new_n675), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g475(.A(new_n635), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n668), .A2(G15gat), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G15gat), .B1(new_n668), .B2(new_n627), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT106), .ZN(G1326gat));
  NAND3_X1  g480(.A1(new_n349), .A2(new_n409), .A3(new_n667), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT107), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT43), .B(G22gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  NAND2_X1  g484(.A1(new_n591), .A2(new_n632), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n634), .A2(new_n637), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n323), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n666), .ZN(new_n689));
  INV_X1    g488(.A(new_n348), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n320), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n629), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT108), .B1(new_n688), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n560), .B1(new_n494), .B2(new_n495), .ZN(new_n699));
  INV_X1    g498(.A(new_n553), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT38), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n557), .B2(new_n486), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n408), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n571), .B1(new_n570), .B2(new_n581), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n588), .A2(KEYINPUT85), .A3(new_n589), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n631), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n630), .A2(KEYINPUT109), .A3(new_n409), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n627), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n687), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n697), .A3(new_n287), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n714), .B(KEYINPUT44), .C1(new_n638), .C2(new_n323), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n693), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n629), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n696), .A2(new_n718), .ZN(G1328gat));
  OAI21_X1  g518(.A(G36gat), .B1(new_n717), .B2(new_n570), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n694), .A2(G36gat), .A3(new_n570), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(G1329gat));
  OAI21_X1  g522(.A(new_n209), .B1(new_n694), .B2(new_n677), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n625), .A2(G43gat), .A3(new_n626), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n717), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n715), .A2(new_n713), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n627), .A2(new_n631), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n705), .A2(new_n706), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(new_n562), .ZN(new_n732));
  INV_X1    g531(.A(new_n687), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n287), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n714), .B1(new_n734), .B2(KEYINPUT44), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n409), .B(new_n693), .C1(new_n729), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT110), .B1(new_n736), .B2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n409), .A2(new_n207), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n691), .B1(new_n740), .B2(KEYINPUT111), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n741), .B(new_n323), .C1(KEYINPUT111), .C2(new_n740), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n667), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(KEYINPUT48), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n738), .A2(new_n739), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n716), .A2(KEYINPUT112), .A3(new_n409), .A4(new_n693), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n736), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n743), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n728), .B(new_n745), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(G50gat), .A3(new_n746), .ZN(new_n753));
  INV_X1    g552(.A(new_n743), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n744), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n737), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT113), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n752), .A2(new_n758), .ZN(G1331gat));
  NAND4_X1  g558(.A1(new_n325), .A2(new_n666), .A3(new_n690), .A4(new_n712), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n629), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n289), .ZN(G1332gat));
  AOI21_X1  g561(.A(new_n570), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT114), .Z(new_n764));
  NOR2_X1   g563(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1333gat));
  OAI21_X1  g566(.A(G71gat), .B1(new_n760), .B2(new_n627), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n635), .A2(new_n293), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n760), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1334gat));
  NOR2_X1   g571(.A1(new_n760), .A2(new_n408), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n294), .ZN(G1335gat));
  INV_X1    g573(.A(new_n716), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n666), .A2(new_n321), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n690), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT116), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n775), .A2(new_n781), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n629), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n712), .A2(new_n287), .A3(new_n777), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT51), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n348), .A2(G85gat), .A3(new_n629), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT118), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(G1336gat));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(G92gat), .C1(new_n780), .C2(new_n570), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n787), .A2(new_n348), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n570), .A2(G92gat), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(KEYINPUT52), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n793), .A2(new_n795), .A3(new_n794), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n588), .A3(new_n783), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(G92gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n800), .B2(new_n791), .ZN(G1337gat));
  AOI21_X1  g600(.A(G99gat), .B1(new_n793), .B2(new_n635), .ZN(new_n802));
  INV_X1    g601(.A(new_n784), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n625), .A2(G99gat), .A3(new_n626), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(G1338gat));
  XNOR2_X1  g604(.A(KEYINPUT120), .B(G106gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n780), .B2(new_n408), .ZN(new_n807));
  NOR4_X1   g606(.A1(new_n787), .A2(G106gat), .A3(new_n408), .A4(new_n348), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n782), .A2(new_n409), .A3(new_n783), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(new_n806), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(G1339gat));
  NAND4_X1  g613(.A1(new_n322), .A2(new_n666), .A3(new_n324), .A4(new_n348), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n345), .B2(new_n327), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n336), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n346), .A2(new_n816), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n342), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n342), .A4(new_n819), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n823), .A3(new_n344), .ZN(new_n824));
  INV_X1    g623(.A(new_n655), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n825), .A2(KEYINPUT18), .B1(new_n648), .B2(new_n650), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n655), .A2(new_n664), .A3(new_n652), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n663), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n648), .A2(new_n650), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n643), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n323), .A2(new_n824), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n824), .A2(new_n666), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n348), .A2(new_n832), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n834), .A2(new_n835), .B1(new_n282), .B2(new_n286), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n321), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n629), .B1(new_n815), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n633), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n838), .A2(new_n570), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n689), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n409), .B1(new_n815), .B2(new_n837), .ZN(new_n842));
  INV_X1    g641(.A(new_n629), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n570), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n635), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n499), .A3(new_n666), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n841), .A2(new_n847), .ZN(G1340gat));
  AOI21_X1  g647(.A(G120gat), .B1(new_n840), .B2(new_n690), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n846), .A2(new_n500), .A3(new_n348), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(G1341gat));
  NAND3_X1  g650(.A1(new_n840), .A2(new_n514), .A3(new_n320), .ZN(new_n852));
  OAI21_X1  g651(.A(G127gat), .B1(new_n846), .B2(new_n321), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1342gat));
  NAND3_X1  g653(.A1(new_n840), .A2(new_n512), .A3(new_n287), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n846), .B2(new_n323), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(G1343gat));
  NOR2_X1   g658(.A1(new_n348), .A2(new_n832), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT123), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n834), .A2(new_n861), .B1(new_n286), .B2(new_n282), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n321), .B1(new_n833), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n815), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(KEYINPUT57), .A3(new_n409), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n408), .B1(new_n815), .B2(new_n837), .ZN(new_n866));
  XOR2_X1   g665(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n845), .A2(new_n627), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT121), .Z(new_n870));
  NAND4_X1  g669(.A1(new_n868), .A2(G141gat), .A3(new_n689), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n627), .A2(new_n409), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n588), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n838), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n353), .B1(new_n874), .B2(new_n666), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n876), .B(new_n877), .ZN(G1344gat));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n833), .B2(new_n862), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n834), .A2(new_n861), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n323), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n824), .A2(new_n832), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n287), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT124), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n880), .A2(new_n885), .A3(new_n321), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n815), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n409), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n866), .A2(new_n867), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n690), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT59), .B(G148gat), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT59), .B1(new_n874), .B2(new_n348), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n891), .A2(KEYINPUT59), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n893), .A2(new_n354), .B1(new_n868), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1345gat));
  INV_X1    g695(.A(new_n874), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n359), .A3(new_n320), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n868), .A2(new_n320), .A3(new_n870), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n900), .B2(new_n359), .ZN(G1346gat));
  NAND3_X1  g700(.A1(new_n897), .A2(new_n360), .A3(new_n287), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n868), .A2(new_n287), .A3(new_n870), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n902), .B1(new_n904), .B2(new_n360), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n570), .A2(new_n843), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n677), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n842), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n430), .A3(new_n666), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n815), .B2(new_n837), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n839), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n689), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n430), .B2(new_n914), .ZN(G1348gat));
  OAI21_X1  g714(.A(G176gat), .B1(new_n909), .B2(new_n348), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n690), .A2(new_n431), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n912), .B2(new_n917), .ZN(G1349gat));
  NAND3_X1  g717(.A1(new_n913), .A2(new_n423), .A3(new_n320), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n909), .A2(new_n321), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n425), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n921), .B(new_n922), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n913), .A2(new_n205), .A3(new_n287), .ZN(new_n924));
  OAI21_X1  g723(.A(G190gat), .B1(new_n909), .B2(new_n323), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n627), .A2(new_n906), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n689), .B(new_n930), .C1(new_n888), .C2(new_n889), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G197gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n872), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n911), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n666), .A2(G197gat), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n929), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT126), .B(new_n936), .C1(new_n931), .C2(G197gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(G1352gat));
  INV_X1    g739(.A(G204gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n941), .A3(new_n690), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT62), .Z(new_n943));
  OAI21_X1  g742(.A(new_n930), .B1(new_n888), .B2(new_n889), .ZN(new_n944));
  OAI21_X1  g743(.A(G204gat), .B1(new_n944), .B2(new_n348), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1353gat));
  INV_X1    g745(.A(G211gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n934), .A2(new_n947), .A3(new_n320), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n320), .B(new_n930), .C1(new_n888), .C2(new_n889), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  AOI21_X1  g751(.A(G218gat), .B1(new_n934), .B2(new_n287), .ZN(new_n953));
  OAI211_X1 g752(.A(KEYINPUT127), .B(new_n930), .C1(new_n888), .C2(new_n889), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(new_n375), .A3(new_n287), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n944), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n953), .B1(new_n955), .B2(new_n957), .ZN(G1355gat));
endmodule


