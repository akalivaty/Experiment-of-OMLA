//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G116), .A2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n213), .B(new_n214), .C1(new_n202), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT65), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n216), .A2(new_n217), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G87), .A2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n205), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  INV_X1    g0026(.A(G1), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT64), .Z(new_n234));
  AOI211_X1 g0034(.A(new_n212), .B(new_n226), .C1(new_n232), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G222), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n252), .B1(new_n253), .B2(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n229), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n259), .B(new_n263), .C1(G77), .C2(new_n252), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n227), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n262), .A2(new_n265), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n264), .B(new_n268), .C1(new_n215), .C2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT68), .ZN(new_n272));
  INV_X1    g0072(.A(G200), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n274), .A2(KEYINPUT73), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(KEYINPUT73), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(G190), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n227), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n227), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n209), .A2(new_n260), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n229), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n282), .B(new_n284), .C1(G1), .C2(new_n231), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n285), .A2(new_n202), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n203), .A2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  XOR2_X1   g0090(.A(KEYINPUT8), .B(G58), .Z(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n231), .A2(G33), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n287), .B1(new_n288), .B2(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n284), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n282), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n202), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n286), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT9), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n275), .A2(new_n276), .A3(new_n277), .A4(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT10), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n272), .A2(G169), .ZN(new_n303));
  INV_X1    g0103(.A(new_n299), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n272), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G238), .ZN(new_n310));
  INV_X1    g0110(.A(G232), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n252), .B1(new_n310), .B2(new_n254), .C1(new_n257), .C2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(new_n263), .C1(G107), .C2(new_n252), .ZN(new_n313));
  INV_X1    g0113(.A(G244), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n268), .C1(new_n314), .C2(new_n270), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(G179), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT71), .ZN(new_n317));
  INV_X1    g0117(.A(new_n285), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n291), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n319));
  OR2_X1    g0119(.A1(KEYINPUT15), .A2(G87), .ZN(new_n320));
  NAND2_X1  g0120(.A1(KEYINPUT15), .A2(G87), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT70), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT70), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n319), .B1(new_n326), .B2(new_n293), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n318), .A2(G77), .B1(new_n295), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G77), .B2(new_n282), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n315), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n332), .A2(KEYINPUT72), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(KEYINPUT72), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n317), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT67), .B(G1698), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n338), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n337), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n263), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n269), .A2(G238), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n268), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT13), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n345), .A2(new_n349), .A3(new_n268), .A4(new_n346), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G169), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n350), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT74), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n347), .A2(new_n355), .A3(KEYINPUT13), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G179), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G77), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n293), .A2(new_n361), .B1(new_n231), .B2(G68), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT75), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n290), .A2(new_n202), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n295), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT11), .ZN(new_n366));
  INV_X1    g0166(.A(G68), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT12), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n297), .B2(new_n367), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n282), .A2(KEYINPUT12), .A3(G68), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n366), .B1(new_n367), .B2(new_n285), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n360), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n341), .ZN(new_n373));
  AND2_X1   g0173(.A1(KEYINPUT76), .A2(G33), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT76), .A2(G33), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT7), .B1(new_n377), .B2(G20), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT76), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n260), .ZN(new_n380));
  NAND2_X1  g0180(.A1(KEYINPUT76), .A2(G33), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(KEYINPUT3), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n341), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(new_n231), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(G68), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(G58), .B(G68), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(KEYINPUT16), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n384), .A2(G20), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT3), .B1(new_n380), .B2(new_n381), .ZN(new_n391));
  INV_X1    g0191(.A(new_n342), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n384), .B1(new_n252), .B2(G20), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n367), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n388), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n389), .B(new_n295), .C1(KEYINPUT16), .C2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n267), .B1(new_n269), .B2(G232), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n257), .A2(new_n253), .B1(new_n215), .B2(new_n254), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(new_n377), .B1(G33), .B2(G87), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n262), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G190), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n292), .A2(new_n282), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n318), .B2(new_n292), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(G200), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n398), .A2(new_n404), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n398), .A2(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n402), .A2(new_n330), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n399), .B(new_n305), .C1(new_n262), .C2(new_n401), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n410), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n414), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .A3(new_n410), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n329), .B1(G200), .B2(new_n315), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n315), .A2(new_n403), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n372), .A2(new_n409), .A3(new_n423), .A4(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n371), .B1(new_n357), .B2(G190), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n351), .A2(G200), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR4_X1   g0232(.A1(new_n309), .A2(new_n336), .A3(new_n428), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n282), .A2(G97), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n227), .A2(G33), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n282), .A2(new_n284), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n434), .B1(new_n437), .B2(G97), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n206), .B1(new_n393), .B2(new_n394), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT78), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(KEYINPUT6), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT6), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(KEYINPUT78), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n442), .A2(new_n444), .B1(new_n205), .B2(G107), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(KEYINPUT78), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n441), .A2(KEYINPUT6), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G97), .A2(G107), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n207), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(G20), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n289), .A2(G77), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n295), .B1(new_n440), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT79), .B(new_n295), .C1(new_n440), .C2(new_n452), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n439), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n458));
  NAND2_X1  g0258(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n314), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(new_n341), .A3(new_n382), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT4), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n341), .A2(new_n342), .A3(G250), .A4(G1698), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(KEYINPUT4), .B(G244), .C1(new_n255), .C2(new_n256), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT80), .B1(new_n468), .B2(new_n343), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n460), .A2(new_n470), .A3(KEYINPUT4), .A4(new_n252), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n463), .A2(new_n467), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n263), .ZN(new_n473));
  INV_X1    g0273(.A(G45), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G41), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n266), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n262), .A2(new_n479), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n480), .B1(new_n482), .B2(G257), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n457), .B1(new_n403), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n473), .A2(KEYINPUT81), .A3(new_n483), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(G200), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n487), .A2(new_n491), .A3(G200), .A4(new_n488), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n485), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT22), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n231), .A2(G87), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n343), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n206), .A2(G20), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT23), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n498), .B(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(G116), .B1(new_n374), .B2(new_n375), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n497), .B(new_n500), .C1(G20), .C2(new_n501), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n383), .A2(new_n495), .A3(new_n496), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n494), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n501), .ZN(new_n505));
  INV_X1    g0305(.A(new_n496), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n252), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n505), .A2(new_n231), .B1(new_n507), .B2(new_n495), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n377), .A2(KEYINPUT22), .A3(new_n506), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT24), .A4(new_n500), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n295), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n437), .A2(G107), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n282), .A2(G107), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT25), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n338), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n516));
  INV_X1    g0316(.A(G294), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n516), .A2(new_n383), .B1(new_n517), .B2(new_n376), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(new_n263), .B1(G264), .B2(new_n482), .ZN(new_n519));
  INV_X1    g0319(.A(new_n480), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n515), .B1(G200), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n521), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G190), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n390), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n340), .B1(new_n374), .B2(new_n375), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n342), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT7), .B1(new_n343), .B2(new_n231), .ZN(new_n530));
  OAI21_X1  g0330(.A(G107), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(new_n451), .A3(new_n450), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT79), .B1(new_n532), .B2(new_n295), .ZN(new_n533));
  INV_X1    g0333(.A(new_n456), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n438), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n473), .A2(new_n305), .A3(new_n483), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n469), .A2(new_n471), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n466), .B1(new_n461), .B2(new_n462), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n262), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n483), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n330), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n493), .A2(new_n526), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n523), .A2(new_n305), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n521), .A2(new_n330), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n515), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G20), .ZN(new_n549));
  AOI21_X1  g0349(.A(G20), .B1(G33), .B2(G283), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n260), .A2(G97), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT85), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT85), .B1(new_n550), .B2(new_n551), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n295), .B(new_n549), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT20), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n552), .B(new_n553), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n295), .A4(new_n549), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n297), .A2(new_n548), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT84), .B1(new_n436), .B2(new_n548), .ZN(new_n563));
  OR3_X1    g0363(.A1(new_n436), .A2(KEYINPUT84), .A3(new_n548), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n338), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(G303), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n566), .A2(new_n383), .B1(new_n567), .B2(new_n252), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n263), .B1(G270), .B2(new_n482), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n520), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n565), .A2(new_n571), .A3(G179), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(KEYINPUT21), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n330), .B1(new_n569), .B2(new_n520), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n565), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n574), .B1(new_n565), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n547), .B(new_n572), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n570), .A2(G200), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n561), .A2(new_n562), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n564), .A2(new_n563), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n569), .A2(G190), .A3(new_n520), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n475), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n266), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n262), .A2(G250), .A3(new_n584), .ZN(new_n587));
  OAI21_X1  g0387(.A(G238), .B1(new_n255), .B2(new_n256), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n314), .A2(new_n254), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n505), .B1(new_n377), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n586), .B(new_n587), .C1(new_n592), .C2(new_n262), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G200), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n589), .B1(new_n338), .B2(G238), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n501), .B1(new_n595), .B2(new_n383), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n263), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n597), .A2(G190), .A3(new_n586), .A4(new_n587), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT19), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(new_n231), .A3(G33), .A4(G97), .ZN(new_n600));
  NOR2_X1   g0400(.A1(G97), .A2(G107), .ZN(new_n601));
  INV_X1    g0401(.A(G87), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n601), .A2(new_n602), .B1(new_n337), .B2(new_n231), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n600), .B1(new_n603), .B2(new_n599), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n382), .A2(new_n231), .A3(G68), .A4(new_n341), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n284), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(G87), .A2(new_n282), .A3(new_n284), .A4(new_n435), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n282), .B1(new_n325), .B2(new_n323), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n594), .A2(new_n598), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n593), .A2(G169), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n597), .A2(G179), .A3(new_n586), .A4(new_n587), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n436), .A2(new_n326), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n615), .A2(new_n606), .A3(new_n608), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n613), .B1(new_n611), .B2(new_n612), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n583), .B(new_n610), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n578), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n433), .A2(new_n544), .A3(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n490), .A2(new_n492), .ZN(new_n623));
  INV_X1    g0423(.A(new_n485), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n543), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n594), .A2(new_n598), .A3(new_n609), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n616), .B1(new_n611), .B2(new_n612), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n587), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n596), .B2(new_n263), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n330), .B1(new_n631), .B2(new_n586), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n310), .B1(new_n458), .B2(new_n459), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n341), .B(new_n382), .C1(new_n633), .C2(new_n589), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n262), .B1(new_n634), .B2(new_n501), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n635), .A2(new_n305), .A3(new_n585), .A4(new_n630), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n617), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n610), .A3(KEYINPUT87), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n629), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n625), .A2(new_n525), .A3(new_n578), .A4(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n610), .B1(new_n618), .B2(new_n619), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT26), .B1(new_n641), .B2(new_n542), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n535), .A2(KEYINPUT88), .A3(new_n536), .A4(new_n541), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT88), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n541), .A2(new_n536), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n457), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(new_n639), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n640), .A2(new_n637), .A3(new_n642), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n433), .A2(new_n650), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n431), .A2(new_n336), .B1(new_n371), .B2(new_n360), .ZN(new_n652));
  INV_X1    g0452(.A(new_n409), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n423), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n307), .B1(new_n302), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(new_n547), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n227), .A2(new_n231), .A3(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT89), .ZN(new_n660));
  INV_X1    g0460(.A(G213), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n658), .B2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(KEYINPUT89), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n515), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n657), .B1(new_n525), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n666), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n657), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(new_n673));
  INV_X1    g0473(.A(new_n583), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n565), .A2(new_n666), .ZN(new_n675));
  OR3_X1    g0475(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n676), .A2(KEYINPUT90), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n673), .A2(KEYINPUT90), .A3(new_n675), .ZN(new_n678));
  OAI211_X1 g0478(.A(G330), .B(new_n672), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n672), .A2(new_n673), .A3(new_n669), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n670), .A3(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n210), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n233), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n646), .A4(new_n643), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT92), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT92), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n647), .A2(new_n692), .A3(KEYINPUT26), .A4(new_n639), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n648), .B1(new_n641), .B2(new_n542), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT93), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g0496(.A(KEYINPUT93), .B(new_n648), .C1(new_n641), .C2(new_n542), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n691), .A2(new_n693), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n637), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT94), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(KEYINPUT94), .A3(new_n637), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n640), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n689), .B1(new_n703), .B2(new_n669), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n625), .A2(new_n525), .A3(new_n621), .A4(new_n669), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT91), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n484), .A2(new_n521), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(new_n569), .A3(new_n636), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n569), .A4(new_n636), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n484), .A2(new_n570), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n305), .A3(new_n521), .A4(new_n593), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n666), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(new_n666), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT91), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n544), .A2(new_n720), .A3(new_n621), .A4(new_n669), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n706), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G330), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n650), .A2(new_n669), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n704), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n688), .B1(new_n728), .B2(G1), .ZN(G364));
  OR2_X1    g0529(.A1(new_n677), .A2(new_n678), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(G330), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n228), .A2(new_n474), .A3(G20), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(KEYINPUT95), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(G1), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n683), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n731), .A2(new_n732), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n231), .A2(new_n305), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n403), .A2(new_n273), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT99), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n743), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n231), .A2(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n403), .A3(G200), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n747), .A2(new_n202), .B1(new_n206), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n740), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n750), .B1(G77), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n740), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n755), .A2(new_n273), .A3(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n403), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n231), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n754), .B1(new_n367), .B2(new_n757), .C1(new_n205), .C2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n740), .A2(G190), .A3(new_n273), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT98), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n761), .B(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G58), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n741), .A2(new_n748), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G87), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n748), .A2(new_n751), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n769), .B1(new_n773), .B2(KEYINPUT32), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT32), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n252), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n760), .A2(new_n766), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n756), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n770), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n780), .A2(KEYINPUT100), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(KEYINPUT100), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n252), .B(new_n779), .C1(new_n784), .C2(G329), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n785), .B1(new_n517), .B2(new_n759), .C1(new_n567), .C2(new_n767), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n761), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G326), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n747), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n749), .B1(new_n752), .B2(new_n792), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n786), .A2(new_n788), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n777), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n230), .B1(G20), .B2(new_n330), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n247), .A2(G45), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n234), .A2(new_n474), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n377), .A2(new_n682), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(G355), .B(KEYINPUT96), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(new_n210), .A3(new_n252), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n800), .B(new_n802), .C1(G116), .C2(new_n210), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT97), .Z(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n796), .A2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n795), .A2(new_n796), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n807), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n730), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n739), .B1(new_n738), .B2(new_n811), .ZN(G396));
  NOR2_X1   g0612(.A1(new_n336), .A2(new_n427), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n329), .A2(new_n666), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n335), .A2(KEYINPUT101), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n335), .B2(KEYINPUT101), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n813), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n726), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n817), .A2(new_n650), .A3(new_n669), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(new_n725), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n738), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n818), .A2(new_n805), .ZN(new_n824));
  INV_X1    g0624(.A(new_n747), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n825), .A2(G137), .B1(G143), .B2(new_n763), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n288), .B2(new_n757), .C1(new_n771), .C2(new_n752), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT34), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n202), .B2(new_n767), .C1(new_n829), .C2(new_n783), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n749), .A2(new_n367), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n759), .A2(new_n765), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n830), .A2(new_n383), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n343), .B1(new_n517), .B2(new_n761), .C1(new_n757), .C2(new_n791), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n825), .A2(G303), .B1(G107), .B2(new_n768), .ZN(new_n835));
  INV_X1    g0635(.A(new_n759), .ZN(new_n836));
  INV_X1    g0636(.A(new_n749), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(G97), .B1(new_n837), .B2(G87), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n835), .B(new_n838), .C1(new_n792), .C2(new_n783), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n834), .B(new_n839), .C1(G116), .C2(new_n753), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n796), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n796), .A2(new_n805), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n361), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n824), .A2(new_n841), .A3(new_n737), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n823), .A2(new_n844), .ZN(G384));
  NAND2_X1  g0645(.A1(new_n445), .A2(new_n449), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT35), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n231), .B(new_n230), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n848), .B(G116), .C1(new_n847), .C2(new_n846), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT36), .ZN(new_n850));
  OAI21_X1  g0650(.A(G77), .B1(new_n765), .B2(new_n367), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n851), .A2(new_n233), .B1(G50), .B2(new_n367), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(G1), .A3(new_n228), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n433), .A2(new_n725), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n372), .A2(new_n669), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT102), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n372), .B(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n429), .A2(new_n430), .B1(new_n371), .B2(new_n666), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n723), .A2(new_n859), .A3(KEYINPUT40), .A4(new_n818), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  INV_X1    g0661(.A(new_n664), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n410), .A2(new_n862), .ZN(new_n863));
  AND4_X1   g0663(.A1(new_n861), .A2(new_n417), .A3(new_n408), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n389), .A2(new_n295), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT16), .B1(new_n386), .B2(new_n388), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n406), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n421), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n862), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n408), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n864), .B1(KEYINPUT37), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n423), .B2(new_n409), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n423), .A2(new_n409), .ZN(new_n875));
  INV_X1    g0675(.A(new_n869), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n410), .B1(new_n421), .B2(new_n862), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n861), .A3(new_n408), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n861), .B1(new_n879), .B2(new_n408), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n864), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n863), .B1(new_n423), .B2(new_n409), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n873), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n877), .A2(new_n881), .A3(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n372), .A2(new_n856), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT102), .B1(new_n360), .B2(new_n371), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n858), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n855), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n890), .A2(new_n895), .A3(new_n722), .A4(new_n817), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n860), .A2(new_n884), .B1(KEYINPUT40), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n854), .B1(new_n897), .B2(new_n724), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(new_n723), .ZN(new_n899));
  INV_X1    g0699(.A(new_n433), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n433), .B1(new_n704), .B2(new_n727), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n655), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n901), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n857), .A2(new_n666), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n888), .A2(new_n889), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n873), .B1(new_n871), .B2(new_n872), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n909), .B2(new_n889), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT103), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT103), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n888), .A2(new_n889), .A3(new_n907), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(new_n883), .C2(new_n907), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n906), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n336), .A2(new_n669), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n859), .B1(new_n820), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n917), .A2(new_n884), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n423), .A2(new_n862), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n915), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n904), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n227), .B1(G13), .B2(new_n231), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n850), .B(new_n853), .C1(new_n922), .C2(new_n923), .ZN(G367));
  OAI21_X1  g0724(.A(new_n639), .B1(new_n609), .B2(new_n669), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT104), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n637), .A2(new_n609), .A3(new_n669), .ZN(new_n928));
  MUX2_X1   g0728(.A(new_n927), .B(new_n926), .S(new_n928), .Z(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n666), .B(new_n493), .C1(new_n542), .C2(new_n547), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n625), .ZN(new_n933));
  INV_X1    g0733(.A(new_n578), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n680), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n930), .B(new_n932), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n535), .A2(new_n666), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n625), .A2(new_n941), .B1(new_n543), .B2(new_n666), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n679), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n944));
  INV_X1    g0744(.A(new_n930), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n940), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n943), .B1(new_n940), .B2(new_n947), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT109), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n673), .A2(new_n669), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n670), .B1(new_n668), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n942), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT45), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT44), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT106), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n942), .A2(new_n958), .A3(new_n954), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n958), .B1(new_n942), .B2(new_n954), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n961), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(KEYINPUT44), .A3(new_n959), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n956), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n679), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n679), .B(KEYINPUT107), .Z(new_n968));
  AND2_X1   g0768(.A1(new_n968), .A2(new_n965), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n967), .B1(new_n969), .B2(KEYINPUT108), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n965), .A3(KEYINPUT108), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n672), .B(new_n953), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n732), .B(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n728), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n728), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n683), .B(KEYINPUT41), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n951), .B(new_n952), .C1(new_n977), .C2(new_n736), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n736), .B1(new_n975), .B2(new_n976), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n940), .A2(new_n947), .ZN(new_n980));
  INV_X1    g0780(.A(new_n943), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n948), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT109), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n799), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n808), .B1(new_n210), .B2(new_n326), .C1(new_n986), .C2(new_n242), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n377), .B1(G107), .B2(new_n836), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n749), .A2(new_n205), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G283), .B2(new_n753), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(new_n764), .C2(new_n567), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n768), .A2(G116), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT46), .ZN(new_n993));
  INV_X1    g0793(.A(G317), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n992), .A2(new_n993), .B1(new_n994), .B2(new_n770), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n747), .A2(new_n792), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n992), .A2(new_n993), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n995), .B(new_n996), .C1(KEYINPUT110), .C2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(KEYINPUT110), .B2(new_n997), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n991), .B(new_n999), .C1(G294), .C2(new_n756), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n756), .A2(G159), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n836), .A2(G68), .ZN(new_n1002));
  INV_X1    g0802(.A(G143), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n765), .B2(new_n767), .C1(new_n747), .C2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n749), .A2(new_n361), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n252), .B1(new_n752), .B2(new_n202), .ZN(new_n1006));
  INV_X1    g0806(.A(G137), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n761), .A2(new_n288), .B1(new_n770), .B2(new_n1007), .ZN(new_n1008));
  NOR4_X1   g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1000), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT47), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n796), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n737), .B(new_n987), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n929), .A2(new_n810), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n985), .A2(new_n1016), .ZN(G387));
  AOI22_X1  g0817(.A1(new_n763), .A2(G317), .B1(G303), .B2(new_n753), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT112), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n792), .B2(new_n757), .C1(new_n787), .C2(new_n747), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n791), .B2(new_n759), .C1(new_n517), .C2(new_n767), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT49), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n749), .A2(new_n548), .B1(new_n770), .B2(new_n789), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n383), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n326), .A2(new_n759), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G68), .B2(new_n753), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n288), .B2(new_n770), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n761), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n989), .B(new_n1029), .C1(G50), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n756), .A2(new_n291), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n767), .A2(new_n361), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n383), .B1(new_n825), .B2(G159), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1012), .B1(new_n1026), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n672), .A2(new_n810), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1037), .A2(new_n738), .A3(new_n1038), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n292), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n685), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(G68), .A2(G77), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT50), .B1(new_n292), .B2(G50), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1042), .A2(new_n474), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1045), .B(new_n799), .C1(new_n474), .C2(new_n239), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1041), .A2(new_n210), .A3(new_n252), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(G107), .C2(new_n210), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT111), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n808), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1039), .A2(new_n1050), .B1(new_n736), .B2(new_n973), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n728), .A2(new_n973), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n683), .B1(new_n728), .B2(new_n973), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(G393));
  XNOR2_X1  g0855(.A(new_n965), .B(new_n679), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n683), .B1(new_n970), .B2(new_n974), .C1(new_n1053), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n736), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n747), .A2(new_n994), .B1(new_n792), .B2(new_n761), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT52), .Z(new_n1060));
  NOR2_X1   g0860(.A1(new_n757), .A2(new_n567), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n749), .A2(new_n206), .B1(new_n770), .B2(new_n787), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n343), .B1(new_n759), .B2(new_n548), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n791), .B2(new_n767), .C1(new_n517), .C2(new_n752), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT114), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n377), .B1(new_n1003), .B2(new_n770), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n747), .A2(new_n288), .B1(new_n771), .B2(new_n761), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT51), .Z(new_n1069));
  AOI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(G87), .C2(new_n837), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n759), .A2(new_n361), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G50), .B2(new_n756), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(new_n367), .C2(new_n767), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n291), .B2(new_n753), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n796), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n942), .A2(new_n807), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n808), .B1(new_n205), .B2(new_n210), .C1(new_n986), .C2(new_n250), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n737), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT113), .Z(new_n1079));
  NAND3_X1  g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1057), .A2(new_n1058), .A3(new_n1080), .ZN(G390));
  OAI211_X1 g0881(.A(new_n911), .B(new_n914), .C1(new_n917), .C2(new_n905), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n703), .A2(new_n669), .A3(new_n817), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n859), .B1(new_n1083), .B2(new_n916), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n906), .A2(new_n890), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n895), .A2(new_n722), .A3(G330), .A4(new_n817), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1082), .B(new_n1087), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n902), .A2(new_n655), .A3(new_n854), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n722), .A2(G330), .A3(new_n817), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n859), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT115), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n1087), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n820), .A2(new_n916), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(KEYINPUT115), .A3(new_n859), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1083), .A2(new_n916), .A3(new_n1087), .A4(new_n1093), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT116), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n902), .A2(new_n655), .A3(new_n854), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1091), .A2(new_n1100), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n683), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n911), .A2(new_n914), .A3(new_n805), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  AOI22_X1  g0914(.A1(new_n756), .A2(G137), .B1(new_n753), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n784), .A2(G125), .B1(KEYINPUT117), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(G128), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n747), .C1(new_n771), .C2(new_n759), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n343), .B1(new_n1030), .B2(G132), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1119), .B1(new_n202), .B2(new_n749), .C1(new_n1115), .C2(KEYINPUT117), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n768), .A2(G150), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT53), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n252), .B(new_n1071), .C1(G97), .C2(new_n753), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1030), .A2(G116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n756), .A2(G107), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n769), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n783), .A2(new_n517), .B1(new_n747), .B2(new_n791), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1127), .A2(new_n831), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n796), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n842), .A2(new_n292), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1113), .A2(new_n737), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT118), .Z(new_n1133));
  NAND3_X1  g0933(.A1(new_n1089), .A2(new_n736), .A3(new_n1090), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1112), .A2(new_n1133), .A3(new_n1134), .ZN(G378));
  NOR2_X1   g0935(.A1(new_n304), .A2(new_n664), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n309), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n309), .A2(new_n1136), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n805), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n326), .A2(new_n752), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n784), .B2(G283), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n765), .B2(new_n749), .C1(new_n548), .C2(new_n747), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n757), .A2(new_n205), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n761), .A2(new_n206), .ZN(new_n1149));
  NOR4_X1   g0949(.A1(new_n1147), .A2(new_n1033), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1150), .A2(new_n261), .A3(new_n383), .A4(new_n1002), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT119), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT58), .Z(new_n1153));
  INV_X1    g0953(.A(G124), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n260), .B1(new_n770), .B2(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n757), .A2(new_n829), .B1(new_n1117), .B2(new_n761), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G150), .B2(new_n836), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n825), .A2(G125), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G137), .A2(new_n753), .B1(new_n768), .B2(new_n1114), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G41), .B(new_n1155), .C1(new_n1160), .C2(KEYINPUT59), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(KEYINPUT59), .B2(new_n1160), .C1(new_n771), .C2(new_n749), .ZN(new_n1162));
  AOI21_X1  g0962(.A(G41), .B1(new_n374), .B2(KEYINPUT3), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(G50), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n796), .B1(new_n1153), .B2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT120), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n842), .A2(new_n202), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1144), .A2(new_n1166), .A3(new_n737), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1143), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n897), .A2(new_n724), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1143), .B1(new_n897), .B2(new_n724), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1171), .A2(new_n920), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n920), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n736), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1168), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1108), .A2(new_n1091), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1174), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1171), .A2(new_n920), .A3(new_n1172), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n684), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1104), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1179), .B1(new_n1184), .B2(new_n1175), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1177), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n1110), .A3(new_n976), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n859), .A2(new_n805), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n784), .A2(G128), .B1(G137), .B2(new_n763), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n756), .A2(new_n1114), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G150), .A2(new_n753), .B1(new_n768), .B2(G159), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n383), .B1(G58), .B2(new_n837), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT122), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n747), .A2(new_n829), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1196), .B1(KEYINPUT121), .B2(new_n1197), .C1(new_n202), .C2(new_n759), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1194), .B(new_n1198), .C1(KEYINPUT121), .C2(new_n1197), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n784), .A2(G303), .B1(G116), .B2(new_n756), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n206), .B2(new_n752), .C1(new_n517), .C2(new_n747), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n343), .B1(new_n767), .B2(new_n205), .C1(new_n791), .C2(new_n761), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(new_n1201), .A2(new_n1005), .A3(new_n1027), .A4(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n796), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n842), .A2(new_n367), .ZN(new_n1205));
  AND4_X1   g1005(.A1(new_n737), .A2(new_n1190), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1100), .B2(new_n736), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1189), .A2(new_n1207), .ZN(G381));
  NOR2_X1   g1008(.A1(G375), .A2(G378), .ZN(new_n1209));
  INV_X1    g1009(.A(G390), .ZN(new_n1210));
  INV_X1    g1010(.A(G381), .ZN(new_n1211));
  OR2_X1    g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G387), .A2(G384), .A3(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(G407));
  AOI21_X1  g1014(.A(new_n661), .B1(new_n1209), .B2(new_n665), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(G407), .ZN(G409));
  AOI21_X1  g1016(.A(new_n1015), .B1(new_n978), .B2(new_n984), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(G390), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT125), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1212), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1212), .A2(new_n1220), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(G387), .A2(new_n1210), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1221), .B1(new_n1217), .B2(G390), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n1226), .B2(new_n1218), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1184), .A2(new_n1175), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1177), .B1(new_n1228), .B2(new_n976), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(G378), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT123), .B1(new_n1186), .B2(G378), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1177), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n683), .B1(new_n1184), .B2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G378), .B(new_n1233), .C1(new_n1235), .C2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT123), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1231), .B1(new_n1232), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n661), .A2(G343), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT60), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n683), .B(new_n1110), .C1(new_n1188), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT60), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1207), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G384), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1241), .A2(new_n1243), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1227), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1256));
  INV_X1    g1056(.A(G2897), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1251), .B1(new_n1257), .B2(new_n1243), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1249), .A2(G2897), .A3(new_n1242), .A4(new_n1250), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT124), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1243), .A4(new_n1252), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(KEYINPUT123), .A3(G378), .A4(new_n1233), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1242), .B1(new_n1269), .B2(new_n1231), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1270), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1252), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1255), .A2(new_n1262), .A3(new_n1265), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1260), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1270), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1270), .B2(new_n1252), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1230), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(new_n1278), .A2(KEYINPUT62), .A3(new_n1242), .A4(new_n1251), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1275), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1226), .A2(new_n1218), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1222), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1272), .B1(new_n1280), .B2(new_n1283), .ZN(G405));
  OR2_X1    g1084(.A1(new_n1186), .A2(G378), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1269), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1283), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT127), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1227), .A2(new_n1269), .A3(new_n1285), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1288), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1251), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1289), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1227), .B1(new_n1269), .B2(new_n1285), .ZN(new_n1295));
  OAI21_X1  g1095(.A(KEYINPUT127), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n1252), .A3(new_n1290), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1293), .A2(new_n1297), .ZN(G402));
endmodule


