//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT0), .A3(G128), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G137), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  AOI21_X1  g014(.A(G131), .B1(new_n193), .B2(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n201), .A3(new_n196), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n194), .A2(new_n201), .A3(new_n204), .A4(new_n196), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n199), .A2(new_n200), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n198), .A2(G131), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n191), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n195), .A2(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n197), .ZN(new_n211));
  AOI22_X1  g025(.A1(new_n203), .A2(new_n205), .B1(G131), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(new_n188), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  OR3_X1    g032(.A1(new_n209), .A2(new_n218), .A3(KEYINPUT30), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n203), .A2(new_n205), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n198), .A2(new_n200), .A3(G131), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n208), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n191), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n217), .B1(new_n212), .B2(KEYINPUT67), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n211), .A2(G131), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n220), .A2(KEYINPUT67), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n224), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT30), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT2), .B(G113), .Z(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n234), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT66), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n233), .A2(new_n239), .A3(KEYINPUT66), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n230), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n242), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(new_n240), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n224), .B(new_n246), .C1(new_n225), .C2(new_n227), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(G237), .A2(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(KEYINPUT27), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n260));
  OAI21_X1  g074(.A(new_n243), .B1(new_n209), .B2(new_n218), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(new_n247), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n247), .ZN(new_n264));
  INV_X1    g078(.A(new_n260), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT70), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n267), .A3(new_n253), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n255), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n228), .A2(new_n243), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n247), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n258), .B1(new_n272), .B2(KEYINPUT28), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n254), .A2(new_n269), .ZN(new_n274));
  AOI21_X1  g088(.A(G902), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n187), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n264), .A2(new_n259), .A3(new_n265), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n257), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n262), .A2(new_n259), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT71), .B(new_n254), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n247), .A2(KEYINPUT68), .A3(new_n253), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT68), .B1(new_n247), .B2(new_n253), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT31), .B1(new_n286), .B2(new_n244), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n247), .A2(new_n253), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n283), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n246), .B1(new_n219), .B2(new_n229), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n282), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n253), .B1(new_n263), .B2(new_n267), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT72), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n254), .B1(new_n280), .B2(new_n281), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n244), .A2(KEYINPUT31), .A3(new_n283), .A4(new_n290), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n301), .A2(new_n302), .A3(new_n305), .A4(new_n282), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n298), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G472), .A2(G902), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n278), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n308), .ZN(new_n310));
  AOI211_X1 g124(.A(KEYINPUT32), .B(new_n310), .C1(new_n298), .C2(new_n306), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n277), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT24), .B(G110), .Z(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT73), .ZN(new_n314));
  XNOR2_X1  g128(.A(G119), .B(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT74), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n237), .A2(G128), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT23), .B1(new_n213), .B2(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(KEYINPUT75), .B2(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G110), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT76), .Z(new_n325));
  INV_X1    g139(.A(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G125), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n330), .B2(new_n326), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(G146), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n317), .A2(new_n325), .A3(new_n333), .ZN(new_n334));
  OAI22_X1  g148(.A1(new_n314), .A2(new_n315), .B1(new_n323), .B2(G110), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n331), .A2(new_n214), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n329), .A2(new_n214), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G137), .ZN(new_n340));
  INV_X1    g154(.A(G221), .ZN(new_n341));
  INV_X1    g155(.A(G234), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n341), .A2(new_n342), .A3(G953), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n340), .B(new_n343), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G902), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n334), .A2(new_n338), .A3(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n346), .A2(KEYINPUT25), .A3(new_n347), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G217), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(G234), .B2(new_n347), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n346), .A2(new_n348), .ZN(new_n358));
  INV_X1    g172(.A(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n347), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT77), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n356), .A2(new_n357), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n359), .B1(new_n351), .B2(new_n352), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT78), .B1(new_n365), .B2(new_n362), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT9), .B(G234), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n341), .B1(new_n370), .B2(new_n347), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n216), .B(new_n188), .Z(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT79), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G104), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G107), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n374), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n381), .A2(new_n382), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n379), .A2(KEYINPUT81), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n384), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n379), .A2(KEYINPUT81), .ZN(new_n389));
  OAI21_X1  g203(.A(G101), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n372), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n217), .B1(new_n386), .B2(new_n390), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n222), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT12), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(KEYINPUT12), .B(new_n222), .C1(new_n392), .C2(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n392), .A2(KEYINPUT10), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n391), .A2(KEYINPUT82), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n386), .B2(new_n390), .ZN(new_n402));
  OAI211_X1 g216(.A(KEYINPUT10), .B(new_n217), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n385), .A2(new_n384), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n379), .B1(new_n374), .B2(new_n376), .ZN(new_n405));
  OAI21_X1  g219(.A(G101), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n406), .A2(KEYINPUT4), .ZN(new_n407));
  INV_X1    g221(.A(new_n406), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT80), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n410));
  OAI211_X1 g224(.A(KEYINPUT4), .B(new_n386), .C1(new_n406), .C2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n223), .B(new_n407), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n222), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n399), .A2(new_n403), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n398), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G110), .B(G140), .ZN(new_n416));
  INV_X1    g230(.A(G953), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n417), .A2(G227), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n416), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n399), .A2(new_n403), .A3(new_n412), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n222), .ZN(new_n422));
  INV_X1    g236(.A(new_n419), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n414), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(G469), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(G469), .A2(G902), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n398), .A2(new_n414), .A3(new_n423), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n423), .B1(new_n422), .B2(new_n414), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n428), .B(new_n347), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n371), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n426), .A3(new_n425), .ZN(new_n435));
  INV_X1    g249(.A(new_n371), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n223), .A2(G125), .ZN(new_n441));
  INV_X1    g255(.A(G125), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n217), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G224), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G953), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n444), .B(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n243), .B(new_n407), .C1(new_n409), .C2(new_n411), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n232), .A2(KEYINPUT5), .ZN(new_n450));
  INV_X1    g264(.A(new_n236), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n450), .B(G113), .C1(KEYINPUT5), .C2(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n452), .A2(new_n233), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n400), .B2(new_n402), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n454), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n455), .A2(KEYINPUT86), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n456), .A2(KEYINPUT6), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(KEYINPUT6), .A3(new_n458), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n448), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G210), .B1(G237), .B2(G902), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT7), .B(new_n447), .C1(new_n444), .C2(KEYINPUT87), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n447), .A2(KEYINPUT87), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n447), .A2(KEYINPUT7), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n441), .A2(new_n443), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n453), .A2(new_n391), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n455), .B(KEYINPUT8), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n453), .B2(new_n391), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n464), .B(new_n467), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n456), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n462), .A2(new_n347), .A3(new_n463), .A4(new_n473), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n474), .A2(KEYINPUT88), .ZN(new_n475));
  INV_X1    g289(.A(new_n463), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n347), .ZN(new_n477));
  INV_X1    g291(.A(new_n448), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n456), .A2(KEYINPUT6), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n457), .A2(new_n458), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n478), .B1(new_n481), .B2(new_n460), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n476), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT88), .A3(new_n474), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT84), .Z(new_n486));
  XOR2_X1   g300(.A(new_n486), .B(KEYINPUT85), .Z(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n235), .A2(G122), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n491), .B(KEYINPUT94), .Z(new_n492));
  NOR2_X1   g306(.A1(new_n235), .A2(G122), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n489), .B2(new_n490), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n378), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n489), .A2(new_n493), .A3(G107), .ZN(new_n496));
  XNOR2_X1  g310(.A(G128), .B(G143), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n193), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n498), .B2(KEYINPUT93), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(KEYINPUT93), .B2(new_n498), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g315(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n502));
  INV_X1    g316(.A(G143), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(G128), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n497), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(G134), .C1(new_n505), .C2(new_n502), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n489), .A2(new_n493), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n378), .ZN(new_n508));
  OAI221_X1 g322(.A(new_n506), .B1(G134), .B2(new_n505), .C1(new_n508), .C2(new_n496), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n369), .A2(new_n354), .A3(G953), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n501), .A2(KEYINPUT95), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n509), .B(new_n510), .C1(new_n495), .C2(new_n500), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n509), .B1(new_n495), .B2(new_n500), .ZN(new_n515));
  INV_X1    g329(.A(new_n510), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n347), .ZN(new_n519));
  INV_X1    g333(.A(G478), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n519), .B(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n249), .A2(G143), .A3(G214), .ZN(new_n524));
  AOI21_X1  g338(.A(G143), .B1(new_n249), .B2(G214), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT17), .B(G131), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  INV_X1    g341(.A(G131), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n332), .B(new_n526), .C1(new_n529), .C2(KEYINPUT17), .ZN(new_n530));
  OAI211_X1 g344(.A(KEYINPUT18), .B(G131), .C1(new_n524), .C2(new_n525), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT89), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n330), .A2(G146), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT18), .A2(G131), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n337), .A2(new_n533), .B1(new_n527), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n383), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n329), .B(KEYINPUT19), .Z(new_n541));
  OAI211_X1 g355(.A(new_n529), .B(new_n336), .C1(G146), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n539), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n536), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(G475), .A2(G902), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n523), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n540), .A2(KEYINPUT90), .A3(new_n544), .A4(new_n546), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(KEYINPUT20), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n537), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n543), .A2(KEYINPUT91), .ZN(new_n552));
  AOI21_X1  g366(.A(G902), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G475), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n523), .B(new_n556), .C1(new_n545), .C2(new_n547), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n550), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n522), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G952), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n560), .A2(KEYINPUT96), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(KEYINPUT96), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n417), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(G234), .B2(G237), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n566), .B(KEYINPUT97), .Z(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT98), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n564), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n559), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n440), .A2(new_n488), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n312), .A2(new_n368), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT99), .B(G101), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(G3));
  NOR2_X1   g390(.A1(new_n440), .A2(new_n367), .ZN(new_n577));
  INV_X1    g391(.A(new_n306), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n296), .A2(KEYINPUT71), .B1(new_n303), .B2(new_n304), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n302), .B1(new_n579), .B2(new_n301), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n347), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(KEYINPUT100), .A3(G472), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n307), .A2(new_n308), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n298), .B2(new_n306), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n584), .B1(new_n585), .B2(new_n187), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n577), .A2(new_n582), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n486), .B1(new_n483), .B2(new_n474), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n519), .A2(new_n520), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n518), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n517), .A2(KEYINPUT33), .A3(new_n512), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n347), .A2(G478), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n590), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n558), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n570), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n587), .A2(new_n589), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT34), .B(G104), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  INV_X1    g416(.A(new_n558), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n522), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n589), .A2(new_n604), .A3(new_n570), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n587), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G107), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  AND3_X1   g424(.A1(new_n435), .A2(KEYINPUT83), .A3(new_n436), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT83), .B1(new_n435), .B2(new_n436), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n488), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n582), .A2(new_n586), .A3(new_n613), .A4(new_n583), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n345), .A2(KEYINPUT36), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n339), .B(new_n615), .Z(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n361), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n365), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n559), .A3(new_n571), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT37), .B(G110), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G12));
  NAND3_X1  g437(.A1(new_n434), .A2(new_n439), .A3(new_n619), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT102), .B(G900), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n567), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n564), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n603), .A2(new_n522), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n588), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n312), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT103), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n312), .A2(new_n634), .A3(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  NAND2_X1  g451(.A1(new_n475), .A2(new_n484), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n522), .A2(new_n558), .ZN(new_n641));
  INV_X1    g455(.A(new_n486), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n641), .A2(new_n642), .A3(new_n618), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n611), .A2(new_n612), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n627), .B(KEYINPUT39), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n640), .B(new_n643), .C1(new_n646), .C2(KEYINPUT40), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(KEYINPUT40), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n583), .A2(KEYINPUT32), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n307), .A2(new_n278), .A3(new_n308), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n272), .A2(new_n254), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT105), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n244), .B2(new_n286), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n347), .B1(new_n654), .B2(new_n655), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G143), .ZN(G45));
  INV_X1    g475(.A(new_n624), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n596), .A2(new_n558), .A3(new_n628), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT107), .A3(new_n588), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n589), .B2(new_n663), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n312), .A2(new_n662), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  INV_X1    g483(.A(new_n431), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n429), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n347), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G469), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n436), .A3(new_n432), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n599), .A2(new_n589), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n312), .A2(new_n368), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT41), .B(G113), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NOR2_X1   g492(.A1(new_n606), .A2(new_n674), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n312), .A3(new_n368), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n679), .A2(new_n312), .A3(KEYINPUT108), .A4(new_n368), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  NOR2_X1   g499(.A1(new_n674), .A2(new_n589), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n620), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n312), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n581), .A2(new_n691), .A3(G472), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT109), .B1(new_n585), .B2(new_n187), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n356), .A2(new_n363), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT110), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n273), .A2(new_n253), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n310), .B1(new_n698), .B2(new_n305), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n641), .A2(new_n588), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n570), .A3(new_n674), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n694), .A2(new_n696), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  AOI21_X1  g518(.A(new_n699), .B1(new_n692), .B2(new_n693), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n687), .A2(new_n663), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n619), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  NAND2_X1  g522(.A1(new_n638), .A2(new_n642), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n710));
  NOR4_X1   g524(.A1(new_n709), .A2(new_n710), .A3(new_n437), .A4(new_n663), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n312), .A2(new_n696), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n312), .A2(new_n711), .A3(KEYINPUT111), .A4(new_n696), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n709), .A2(new_n437), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n312), .A2(new_n368), .A3(new_n664), .A4(new_n716), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n714), .A2(new_n715), .B1(new_n710), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n528), .ZN(G33));
  NAND4_X1  g533(.A1(new_n312), .A2(new_n368), .A3(new_n629), .A4(new_n716), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G134), .ZN(G36));
  NAND3_X1  g535(.A1(new_n582), .A2(new_n586), .A3(new_n583), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n603), .A2(new_n596), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT43), .Z(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n619), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n420), .A2(new_n424), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n420), .A2(KEYINPUT45), .A3(new_n424), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(G469), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n426), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n426), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n432), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n436), .ZN(new_n740));
  INV_X1    g554(.A(new_n645), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n729), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n709), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n739), .A2(KEYINPUT112), .A3(new_n436), .A4(new_n645), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n727), .A2(new_n728), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n195), .ZN(G39));
  AOI21_X1  g561(.A(new_n276), .B1(new_n649), .B2(new_n650), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n368), .A2(new_n709), .A3(new_n663), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n739), .A2(KEYINPUT47), .A3(new_n436), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT47), .B1(new_n739), .B2(new_n436), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n748), .B(new_n749), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n327), .ZN(G42));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n694), .A2(new_n696), .A3(new_n700), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n724), .A2(new_n564), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n640), .A2(new_n642), .A3(new_n674), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(KEYINPUT50), .A3(new_n758), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT116), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n766), .A3(new_n763), .ZN(new_n767));
  INV_X1    g581(.A(new_n659), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n709), .A2(new_n674), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n769), .A2(new_n368), .A3(new_n564), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n596), .A2(new_n558), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n758), .A2(new_n619), .A3(new_n705), .A4(new_n769), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n740), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n673), .A2(new_n371), .A3(new_n432), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n750), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n743), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(KEYINPUT115), .A3(new_n757), .A4(new_n758), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n757), .A2(new_n758), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n783), .B2(new_n779), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n765), .A2(new_n767), .A3(new_n774), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n758), .A2(new_n312), .A3(new_n696), .A4(new_n769), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n757), .A2(new_n686), .A3(new_n758), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n768), .A2(new_n770), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n597), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n563), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n780), .A2(new_n757), .A3(new_n758), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n764), .A2(KEYINPUT51), .A3(new_n774), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n756), .B1(new_n788), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n786), .A2(new_n787), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT118), .A3(new_n799), .A4(new_n797), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n312), .A2(new_n634), .A3(new_n631), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n634), .B1(new_n312), .B2(new_n631), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n668), .B(new_n707), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n701), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n619), .A2(new_n627), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n659), .A2(new_n433), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n806), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n665), .A2(new_n644), .A3(new_n667), .A4(new_n619), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n748), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n633), .B2(new_n635), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(KEYINPUT52), .A3(new_n707), .A4(new_n812), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n709), .A2(new_n437), .A3(new_n663), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n694), .A2(new_n619), .A3(new_n700), .A4(new_n820), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n709), .A2(new_n522), .A3(new_n558), .A4(new_n627), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n312), .A2(new_n662), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n720), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n714), .A2(new_n715), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n717), .A2(new_n710), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n703), .A2(new_n676), .A3(new_n689), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n682), .B2(new_n683), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n488), .A2(new_n604), .A3(new_n570), .ZN(new_n830));
  OAI22_X1  g644(.A1(new_n587), .A2(new_n830), .B1(new_n614), .B2(new_n620), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n368), .A2(new_n598), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n574), .B1(new_n614), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n832), .B2(new_n831), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n827), .A2(new_n829), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n805), .B1(new_n819), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n828), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n827), .A2(new_n684), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n814), .A2(new_n818), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n836), .A2(new_n833), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n838), .A2(new_n843), .A3(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n804), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(G952), .A2(G953), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n673), .A2(new_n432), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT49), .Z(new_n851));
  INV_X1    g665(.A(new_n487), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n723), .A2(new_n852), .A3(new_n371), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n696), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(new_n640), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n848), .A2(new_n849), .B1(new_n659), .B2(new_n855), .ZN(G75));
  NOR2_X1   g670(.A1(new_n417), .A2(G952), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n347), .B1(new_n838), .B2(new_n843), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n859), .B2(G210), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n481), .A2(new_n460), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT119), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT55), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(new_n478), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n858), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n837), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n867), .B2(new_n841), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n819), .A2(new_n837), .A3(new_n805), .ZN(new_n869));
  OAI21_X1  g683(.A(G902), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n859), .A2(KEYINPUT120), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n476), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n864), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n866), .B1(new_n875), .B2(new_n877), .ZN(G51));
  INV_X1    g692(.A(new_n734), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n426), .B(KEYINPUT57), .Z(new_n881));
  NAND3_X1  g695(.A1(new_n846), .A2(new_n847), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n671), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n857), .B1(new_n880), .B2(new_n883), .ZN(G54));
  AND2_X1   g698(.A1(KEYINPUT58), .A2(G475), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n872), .A2(new_n873), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n545), .ZN(new_n887));
  INV_X1    g701(.A(new_n545), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n872), .A2(new_n888), .A3(new_n873), .A4(new_n885), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n887), .A2(new_n858), .A3(new_n889), .ZN(G60));
  NAND2_X1  g704(.A1(G478), .A2(G902), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT59), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n846), .A2(new_n847), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n893), .A2(new_n594), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n594), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n857), .ZN(G63));
  XOR2_X1   g710(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n897));
  NAND2_X1  g711(.A1(G217), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT60), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n838), .B2(new_n843), .ZN(new_n900));
  INV_X1    g714(.A(new_n358), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n858), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n616), .B(new_n899), .C1(new_n838), .C2(new_n843), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n897), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT123), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n902), .A2(new_n903), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT61), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n908), .B(new_n897), .C1(new_n902), .C2(new_n903), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(G66));
  OAI21_X1  g724(.A(G953), .B1(new_n569), .B2(new_n445), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT124), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n842), .A2(new_n829), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n862), .B1(G898), .B2(new_n417), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G69));
  AOI21_X1  g730(.A(new_n417), .B1(G227), .B2(G900), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n230), .B(KEYINPUT125), .Z(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(new_n541), .Z(new_n919));
  NAND3_X1  g733(.A1(new_n742), .A2(new_n810), .A3(new_n744), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n312), .A2(new_n696), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT126), .ZN(new_n923));
  INV_X1    g737(.A(new_n754), .ZN(new_n924));
  INV_X1    g738(.A(new_n718), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .A4(new_n720), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n746), .A2(new_n809), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n417), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n417), .A2(G900), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT127), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(KEYINPUT127), .A3(new_n930), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n919), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n919), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n312), .A2(new_n368), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n604), .A2(new_n597), .ZN(new_n937));
  NOR4_X1   g751(.A1(new_n936), .A2(new_n646), .A3(new_n709), .A4(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n746), .A2(new_n754), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n660), .A2(new_n817), .A3(new_n707), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n935), .B1(new_n943), .B2(new_n417), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n917), .B1(new_n934), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n933), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n935), .B1(new_n946), .B2(new_n931), .ZN(new_n947));
  INV_X1    g761(.A(new_n917), .ZN(new_n948));
  INV_X1    g762(.A(new_n944), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n950), .ZN(G72));
  INV_X1    g765(.A(new_n248), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n913), .A2(new_n941), .A3(new_n942), .A4(new_n939), .ZN(new_n953));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  AOI211_X1 g769(.A(new_n254), .B(new_n952), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n955), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n926), .A2(new_n927), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(new_n913), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n952), .A2(new_n254), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n858), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n286), .A2(new_n244), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n957), .B1(new_n255), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n956), .B(new_n961), .C1(new_n844), .C2(new_n963), .ZN(G57));
endmodule


