//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OR2_X1    g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT65), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n202), .A2(new_n203), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n215), .A2(new_n216), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n223), .B1(new_n216), .B2(new_n215), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT66), .B(G238), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT67), .B(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI22_X1  g0027(.A1(new_n203), .A2(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n213), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n224), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  INV_X1    g0044(.A(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT68), .B(G107), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n217), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n218), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT69), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n257), .A2(G77), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n260), .A2(new_n261), .B1(new_n218), .B2(G68), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n254), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT11), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n267));
  OR3_X1    g0067(.A1(new_n267), .A2(KEYINPUT12), .A3(G68), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT12), .B1(new_n267), .B2(G68), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n254), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n268), .A2(new_n269), .B1(new_n272), .B2(G68), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n263), .B2(new_n264), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(G1), .B(G13), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n278), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n280), .B1(new_n285), .B2(G238), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n287), .A2(new_n289), .A3(G232), .A4(G1698), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n287), .A2(new_n289), .A3(G226), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G97), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT72), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n294), .B2(new_n296), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n286), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT13), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n286), .C1(new_n297), .C2(new_n298), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n277), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n302), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n305), .A2(G169), .A3(new_n304), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n276), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n310), .B(new_n275), .C1(new_n311), .C2(new_n305), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT74), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT3), .B(G33), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G222), .A3(new_n291), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(G1698), .ZN(new_n317));
  INV_X1    g0117(.A(G223), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n316), .B1(new_n226), .B2(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n296), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n280), .B1(new_n285), .B2(G226), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n254), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT8), .B(G58), .Z(new_n324));
  AOI22_X1  g0124(.A1(new_n257), .A2(new_n324), .B1(G150), .B2(new_n259), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n204), .A2(G20), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n272), .A2(G50), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G50), .B2(new_n267), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n322), .A2(G169), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n322), .A2(new_n306), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n320), .A2(G190), .A3(new_n321), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n322), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT71), .B1(new_n327), .B2(new_n329), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT9), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n327), .A2(KEYINPUT71), .A3(new_n329), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n327), .A2(KEYINPUT71), .A3(new_n329), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT9), .B1(new_n342), .B2(new_n337), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n336), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT10), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(KEYINPUT9), .A3(new_n337), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n336), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n332), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n353), .A2(KEYINPUT77), .A3(new_n271), .ZN(new_n354));
  INV_X1    g0154(.A(new_n267), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n354), .A2(new_n254), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT77), .B1(new_n353), .B2(new_n271), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n356), .A2(new_n357), .B1(new_n355), .B2(new_n353), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT76), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT76), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(G58), .A3(G68), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n363), .A3(new_n220), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n288), .A2(G33), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n368));
  OAI211_X1 g0168(.A(KEYINPUT7), .B(new_n218), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT75), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n315), .B2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n287), .A2(new_n289), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT75), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT7), .A4(new_n218), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n370), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n366), .B1(new_n376), .B2(G68), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n323), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n203), .B1(new_n372), .B2(new_n369), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n366), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n359), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n315), .A2(G226), .A3(G1698), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n287), .A2(new_n289), .A3(G223), .A4(new_n291), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n296), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n280), .B1(new_n285), .B2(G232), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n387), .A2(G179), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n277), .B1(new_n387), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n352), .B1(new_n382), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n375), .A2(new_n372), .ZN(new_n393));
  AOI21_X1  g0193(.A(G20), .B1(new_n287), .B2(new_n289), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n374), .B1(new_n394), .B2(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n365), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n254), .A3(new_n381), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n391), .B1(new_n398), .B2(new_n358), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT18), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n387), .A2(G190), .A3(new_n388), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n334), .B1(new_n387), .B2(new_n388), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(new_n403), .A3(new_n358), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT17), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n398), .A2(new_n403), .A3(new_n406), .A4(new_n358), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n392), .A2(new_n400), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n324), .A2(new_n259), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT15), .B(G87), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n409), .B1(new_n218), .B2(new_n226), .C1(new_n255), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n254), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n272), .A2(G77), .B1(new_n226), .B2(new_n355), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n284), .A2(new_n227), .B1(new_n279), .B2(new_n278), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n315), .A2(G232), .A3(new_n291), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n416), .B1(new_n208), .B2(new_n315), .C1(new_n317), .C2(new_n225), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n415), .B1(new_n417), .B2(new_n296), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n414), .B1(G169), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT70), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n306), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT70), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n414), .B(new_n422), .C1(G169), .C2(new_n418), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n414), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n418), .A2(G190), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n334), .C2(new_n418), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n351), .A2(new_n408), .A3(new_n424), .A4(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n314), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n287), .A2(new_n289), .A3(G250), .A4(new_n291), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n287), .A2(new_n289), .A3(G257), .A4(G1698), .ZN(new_n431));
  INV_X1    g0231(.A(G294), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n430), .B(new_n431), .C1(new_n281), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n296), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n266), .A2(G45), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(KEYINPUT79), .A3(G274), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT5), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G41), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n441), .A2(new_n438), .A3(new_n443), .A4(G274), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n296), .B1(new_n437), .B2(new_n438), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G264), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n434), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n277), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n433), .A2(new_n296), .B1(new_n448), .B2(G264), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n306), .A3(new_n447), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n287), .A2(new_n289), .A3(new_n218), .A4(G87), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n315), .A2(new_n218), .A3(G87), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G116), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n218), .B2(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n208), .A2(KEYINPUT23), .A3(G20), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n457), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT24), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n457), .A2(new_n460), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(KEYINPUT84), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(KEYINPUT84), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n254), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT25), .B1(new_n355), .B2(new_n208), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n208), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n266), .A2(G33), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n267), .A2(new_n478), .A3(new_n217), .A4(new_n253), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n476), .A2(new_n477), .B1(new_n480), .B2(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n454), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n481), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n470), .A2(KEYINPUT84), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n472), .A3(new_n468), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n254), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n450), .A2(new_n334), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G190), .B2(new_n450), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n482), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n267), .A2(G116), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n245), .B2(new_n479), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT78), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n207), .ZN(new_n495));
  NAND2_X1  g0295(.A1(KEYINPUT78), .A2(G97), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n281), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n218), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n253), .A2(new_n217), .B1(G20), .B2(new_n245), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n501), .A2(KEYINPUT20), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT20), .B1(new_n501), .B2(new_n502), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n493), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G303), .B1(new_n367), .B2(new_n368), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n287), .A2(new_n289), .A3(G257), .A4(new_n291), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n287), .A2(new_n289), .A3(G264), .A4(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n296), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n448), .A2(G270), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n447), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n512), .A3(G169), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT20), .ZN(new_n516));
  AND2_X1   g0316(.A1(KEYINPUT78), .A2(G97), .ZN(new_n517));
  NOR2_X1   g0317(.A1(KEYINPUT78), .A2(G97), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n499), .B1(new_n519), .B2(new_n281), .ZN(new_n520));
  INV_X1    g0320(.A(new_n502), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n501), .A2(KEYINPUT20), .A3(new_n502), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n277), .B1(new_n524), .B2(new_n493), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(KEYINPUT21), .A3(new_n512), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n510), .A2(new_n511), .A3(new_n447), .A4(G179), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(KEYINPUT82), .A3(new_n505), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT82), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n492), .B1(new_n522), .B2(new_n523), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n515), .A2(new_n526), .A3(new_n529), .A4(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n512), .A2(G200), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n512), .A2(new_n311), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n534), .A2(new_n535), .A3(new_n505), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n287), .A2(new_n289), .A3(G244), .A4(new_n291), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n315), .A2(KEYINPUT4), .A3(G244), .A4(new_n291), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n315), .A2(G250), .A3(G1698), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n498), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n296), .ZN(new_n544));
  AOI22_X1  g0344(.A1(G257), .A2(new_n448), .B1(new_n439), .B2(new_n446), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n277), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n306), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n208), .A2(KEYINPUT6), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n549), .A2(new_n517), .A3(new_n518), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT6), .B1(new_n209), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(G20), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n259), .A2(G77), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n208), .B1(new_n372), .B2(new_n369), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n254), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n267), .A2(G97), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n480), .B2(G97), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n547), .A2(new_n548), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n546), .A2(G200), .ZN(new_n562));
  INV_X1    g0362(.A(new_n559), .ZN(new_n563));
  INV_X1    g0363(.A(new_n369), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT7), .B1(new_n373), .B2(new_n218), .ZN(new_n565));
  OAI21_X1  g0365(.A(G107), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  INV_X1    g0367(.A(new_n551), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n495), .A2(KEYINPUT6), .A3(new_n208), .A4(new_n496), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n563), .B1(new_n574), .B2(new_n254), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n544), .A2(new_n545), .A3(G190), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n562), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g0377(.A(KEYINPUT15), .B(G87), .Z(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(new_n267), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  XNOR2_X1  g0380(.A(KEYINPUT78), .B(G97), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n255), .ZN(new_n582));
  NOR2_X1   g0382(.A1(G87), .A2(G107), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n517), .B2(new_n518), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n218), .B1(new_n293), .B2(new_n580), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n315), .A2(new_n218), .A3(G68), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n579), .B1(new_n588), .B2(new_n254), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n578), .B(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n480), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n287), .A2(new_n289), .A3(G244), .A4(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n287), .A2(new_n289), .A3(G238), .A4(new_n291), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(new_n461), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n296), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n436), .A2(G250), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n296), .A2(new_n597), .B1(new_n279), .B2(new_n436), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n277), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n595), .B2(new_n296), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n306), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n592), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(G200), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n596), .A2(G190), .A3(new_n599), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT81), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n480), .A2(new_n607), .A3(G87), .ZN(new_n608));
  INV_X1    g0408(.A(G87), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT81), .B1(new_n479), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n605), .A2(new_n589), .A3(new_n606), .A4(new_n611), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n561), .A2(new_n577), .A3(new_n604), .A4(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n429), .A2(new_n489), .A3(new_n537), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(G372));
  NAND3_X1  g0415(.A1(new_n606), .A2(new_n589), .A3(new_n611), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT86), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n600), .B2(G200), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n600), .A2(new_n617), .A3(G200), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n589), .A2(new_n591), .B1(new_n306), .B2(new_n602), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n600), .A2(new_n622), .A3(new_n277), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT85), .B1(new_n602), .B2(G169), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n488), .A2(new_n474), .A3(new_n481), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n561), .A4(new_n577), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n533), .A2(new_n482), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n561), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n626), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n625), .A2(new_n621), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n546), .A2(new_n277), .B1(new_n557), .B2(new_n559), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(new_n548), .A3(new_n604), .A4(new_n612), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n429), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n332), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n405), .A2(new_n407), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n312), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n309), .B2(new_n424), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n392), .A2(new_n400), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n349), .B1(new_n348), .B2(new_n336), .ZN(new_n648));
  AOI211_X1 g0448(.A(KEYINPUT10), .B(new_n335), .C1(new_n346), .C2(new_n347), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n641), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n640), .A2(new_n652), .ZN(G369));
  AND2_X1   g0453(.A1(new_n218), .A2(G13), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n266), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G343), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n505), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT87), .ZN(new_n663));
  MUX2_X1   g0463(.A(new_n533), .B(new_n537), .S(new_n663), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n489), .B1(new_n486), .B2(new_n660), .ZN(new_n667));
  INV_X1    g0467(.A(new_n482), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n660), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n533), .A2(new_n660), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n489), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n668), .B2(new_n661), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n671), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n214), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n581), .A2(new_n245), .A3(new_n583), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n678), .A2(new_n266), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n678), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n221), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT88), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT29), .B1(new_n639), .B2(new_n660), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT89), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n628), .B2(new_n629), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT21), .B1(new_n525), .B2(new_n512), .ZN(new_n688));
  AND4_X1   g0488(.A1(KEYINPUT21), .A2(new_n505), .A3(G169), .A4(new_n512), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n529), .A2(new_n532), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n690), .B(new_n691), .C1(new_n486), .C2(new_n454), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n588), .A2(new_n254), .ZN(new_n693));
  INV_X1    g0493(.A(new_n579), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n693), .A2(new_n611), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT86), .B1(new_n602), .B2(new_n334), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n695), .A2(new_n606), .A3(new_n620), .A4(new_n696), .ZN(new_n697));
  AND4_X1   g0497(.A1(new_n561), .A2(new_n577), .A3(new_n634), .A4(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n692), .A2(KEYINPUT89), .A3(new_n698), .A4(new_n627), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n631), .B1(new_n626), .B2(new_n632), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n634), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n687), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n660), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT90), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT90), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n706), .A3(new_n660), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n685), .B1(new_n708), .B2(KEYINPUT29), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n512), .A2(new_n306), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n450), .A3(new_n546), .A4(new_n600), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n544), .A2(new_n545), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n452), .A2(new_n602), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(new_n528), .A4(KEYINPUT30), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n544), .A2(new_n452), .A3(new_n545), .A4(new_n602), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n527), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n711), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n661), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(KEYINPUT31), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n489), .A2(new_n613), .A3(new_n537), .A4(new_n660), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n719), .A2(KEYINPUT31), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n709), .B1(G330), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n684), .B1(new_n724), .B2(G1), .ZN(G364));
  AOI21_X1  g0525(.A(new_n266), .B1(new_n654), .B2(G45), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n678), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n664), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n311), .A2(G20), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n735), .A2(G179), .A3(new_n334), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G107), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n218), .A2(new_n311), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n306), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n306), .A2(new_n334), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n744), .A2(G87), .B1(new_n747), .B2(G50), .ZN(new_n748));
  NOR4_X1   g0548(.A1(new_n218), .A2(new_n306), .A3(new_n311), .A4(G200), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n735), .A2(new_n306), .A3(new_n334), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n749), .A2(G58), .B1(new_n750), .B2(G68), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n741), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n735), .A2(G179), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G159), .ZN(new_n755));
  OR3_X1    g0555(.A1(new_n754), .A2(KEYINPUT32), .A3(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n311), .A2(G179), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n218), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G97), .ZN(new_n760));
  INV_X1    g0560(.A(new_n226), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n735), .A2(new_n306), .A3(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n373), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT32), .B1(new_n754), .B2(new_n755), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n756), .A2(new_n760), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n749), .A2(G322), .B1(new_n753), .B2(G329), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n315), .B1(new_n747), .B2(G326), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT33), .B(G317), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G311), .A2(new_n762), .B1(new_n750), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n759), .A2(G294), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n766), .A2(new_n767), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n743), .A2(KEYINPUT93), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n743), .A2(KEYINPUT93), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G303), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n774), .A2(new_n775), .B1(new_n739), .B2(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n752), .A2(new_n765), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n217), .B1(G20), .B2(new_n277), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n677), .A2(new_n315), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n251), .A2(G45), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n780), .B(new_n781), .C1(G45), .C2(new_n221), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n677), .A2(new_n373), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n783), .A2(G355), .B1(new_n245), .B2(new_n677), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n732), .A2(new_n779), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n778), .A2(new_n779), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n729), .B1(new_n734), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n665), .A2(KEYINPUT91), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n664), .A2(G330), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n728), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT94), .ZN(G396));
  NAND2_X1  g0594(.A1(new_n639), .A2(new_n660), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n425), .A2(new_n660), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n419), .A2(KEYINPUT70), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n423), .A2(new_n421), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n427), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n420), .A2(new_n421), .A3(new_n796), .A4(new_n423), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n660), .B(new_n802), .C1(new_n630), .C2(new_n638), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n723), .A2(G330), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n729), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT98), .B1(new_n806), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n806), .A2(KEYINPUT98), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G77), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n779), .A2(new_n730), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT95), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n729), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n740), .A2(G87), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n208), .B2(new_n774), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n749), .A2(G294), .B1(new_n753), .B2(G311), .ZN(new_n820));
  INV_X1    g0620(.A(new_n762), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n245), .B2(new_n821), .C1(new_n775), .C2(new_n746), .ZN(new_n822));
  INV_X1    g0622(.A(new_n750), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT96), .B(G283), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n760), .B(new_n373), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n819), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n747), .A2(G137), .B1(new_n762), .B2(G159), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n749), .A2(G143), .B1(new_n750), .B2(G150), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT34), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n315), .B1(new_n758), .B2(new_n202), .C1(new_n754), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n740), .B2(G68), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n833), .B(new_n836), .C1(new_n261), .C2(new_n774), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n829), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n779), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n817), .B1(new_n731), .B2(new_n802), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n812), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  NAND2_X1  g0643(.A1(new_n721), .A2(new_n722), .ZN(new_n844));
  INV_X1    g0644(.A(new_n720), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT106), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT106), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n723), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n429), .A2(new_n850), .A3(G330), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n398), .A2(new_n358), .ZN(new_n853));
  INV_X1    g0653(.A(new_n391), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n659), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n404), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT104), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n855), .A2(new_n856), .A3(new_n860), .A4(new_n404), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n398), .A2(new_n403), .A3(new_n358), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n399), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n864), .A2(KEYINPUT104), .A3(new_n860), .A4(new_n856), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n408), .B2(new_n856), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n852), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n645), .A2(new_n642), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n396), .A2(new_n365), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n379), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n359), .B1(new_n378), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT102), .B1(new_n871), .B2(new_n658), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n397), .A2(new_n254), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n377), .A2(KEYINPUT16), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n358), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT102), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n876), .A3(new_n659), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n875), .A2(new_n854), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n872), .A2(new_n877), .A3(new_n404), .A4(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(new_n861), .ZN(new_n883));
  OAI211_X1 g0683(.A(KEYINPUT38), .B(new_n879), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n867), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n276), .A2(new_n661), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n309), .A2(new_n312), .A3(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n276), .B(new_n661), .C1(new_n307), .C2(new_n308), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n803), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n850), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n802), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n847), .B2(new_n849), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n883), .B1(KEYINPUT37), .B2(new_n881), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n645), .A2(new_n642), .B1(new_n877), .B2(new_n872), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n852), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT40), .B1(new_n896), .B2(new_n884), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n890), .A2(KEYINPUT40), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(G330), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n851), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT107), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n867), .A2(new_n884), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n848), .B1(new_n844), .B2(new_n845), .ZN(new_n903));
  AOI211_X1 g0703(.A(KEYINPUT106), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n889), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT40), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n893), .A2(new_n897), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n429), .A3(new_n850), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n646), .A2(new_n658), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT101), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n420), .A2(new_n421), .A3(new_n423), .A4(new_n660), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT100), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n805), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(new_n805), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n891), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n896), .A2(new_n884), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n911), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT103), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(KEYINPUT103), .B(new_n911), .C1(new_n917), .C2(new_n918), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n867), .A2(new_n884), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n918), .B2(new_n923), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n309), .A2(new_n661), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n910), .B(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n709), .A2(new_n931), .A3(new_n429), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n703), .A2(new_n706), .A3(new_n660), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n706), .B1(new_n703), .B2(new_n660), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT29), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n685), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n429), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT105), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n651), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n930), .A2(new_n940), .B1(new_n266), .B2(new_n654), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n930), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n572), .B(KEYINPUT99), .Z(new_n943));
  INV_X1    g0743(.A(KEYINPUT35), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(G116), .A4(new_n219), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT36), .Z(new_n948));
  NAND4_X1  g0748(.A1(new_n222), .A2(new_n761), .A3(new_n363), .A4(new_n361), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n201), .A2(G68), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n266), .B(G13), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n942), .A2(new_n948), .A3(new_n951), .ZN(G367));
  INV_X1    g0752(.A(new_n780), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n242), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n786), .B1(new_n214), .B2(new_n410), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n728), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n373), .B1(new_n758), .B2(new_n208), .C1(new_n823), .C2(new_n432), .ZN(new_n957));
  INV_X1    g0757(.A(new_n749), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n958), .A2(new_n775), .B1(new_n754), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(G311), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n821), .A2(new_n825), .B1(new_n746), .B2(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n957), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n581), .B2(new_n739), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n245), .ZN(new_n965));
  INV_X1    g0765(.A(new_n774), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(G116), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n965), .B1(new_n967), .B2(KEYINPUT46), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n740), .A2(new_n761), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n373), .B1(new_n747), .B2(G143), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G137), .A2(new_n753), .B1(new_n750), .B2(G159), .ZN(new_n971));
  INV_X1    g0771(.A(new_n201), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n744), .A2(G58), .B1(new_n762), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n759), .A2(G68), .ZN(new_n975));
  INV_X1    g0775(.A(G150), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n976), .B2(new_n958), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT110), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n964), .A2(new_n968), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT47), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n840), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n956), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n626), .B1(new_n695), .B2(new_n660), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n634), .A2(new_n695), .A3(new_n660), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n983), .B1(new_n986), .B2(new_n733), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n561), .B(new_n577), .C1(new_n575), .C2(new_n660), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT108), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n632), .A2(new_n661), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n675), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT44), .Z(new_n993));
  NOR2_X1   g0793(.A1(new_n991), .A2(new_n675), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n671), .ZN(new_n997));
  INV_X1    g0797(.A(new_n674), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n669), .A2(new_n673), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT109), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n1000), .B2(new_n998), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(new_n665), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n724), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n724), .B1(new_n997), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n678), .B(KEYINPUT41), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n727), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n989), .A2(new_n674), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT42), .Z(new_n1010));
  OR2_X1    g0810(.A1(new_n989), .A2(new_n668), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n661), .B1(new_n1011), .B2(new_n561), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1008), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n991), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n671), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1015), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n987), .B1(new_n1007), .B2(new_n1018), .ZN(G387));
  OR2_X1    g0819(.A1(new_n669), .A2(new_n733), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n747), .A2(G322), .B1(new_n762), .B2(G303), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n961), .B2(new_n823), .C1(new_n959), .C2(new_n958), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n432), .B2(new_n743), .C1(new_n758), .C2(new_n825), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n1025));
  XNOR2_X1  g0825(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n315), .B1(new_n753), .B2(G326), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n245), .C2(new_n739), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n744), .A2(new_n761), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n353), .B2(new_n823), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n373), .B(new_n1030), .C1(G150), .C2(new_n753), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n958), .A2(new_n261), .B1(new_n746), .B2(new_n755), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G68), .B2(new_n762), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n740), .A2(G97), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n590), .A2(new_n759), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n840), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n953), .B1(new_n239), .B2(G45), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n679), .B2(new_n783), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n324), .A2(new_n261), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n440), .B1(new_n203), .B2(new_n813), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1041), .A2(new_n679), .A3(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1039), .A2(new_n1043), .B1(G107), .B2(new_n214), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n729), .B(new_n1037), .C1(new_n786), .C2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1003), .A2(new_n727), .B1(new_n1020), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1004), .A2(new_n678), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1003), .A2(new_n724), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT112), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(KEYINPUT112), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(G393));
  AND2_X1   g0852(.A1(new_n1003), .A2(new_n724), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n996), .B(new_n670), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n997), .A2(new_n1004), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n678), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1054), .A2(new_n727), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n953), .A2(new_n248), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n786), .B1(new_n214), .B2(new_n581), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n728), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n958), .A2(new_n755), .B1(new_n746), .B2(new_n976), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT51), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n818), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n753), .A2(G143), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n203), .B2(new_n743), .C1(new_n821), .C2(new_n353), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n315), .B1(new_n758), .B2(new_n813), .C1(new_n823), .C2(new_n201), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1069));
  NOR4_X1   g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT113), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n373), .B1(new_n825), .B2(new_n743), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G294), .A2(new_n762), .B1(new_n753), .B2(G322), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n775), .B2(new_n823), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(G116), .C2(new_n759), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n958), .A2(new_n961), .B1(new_n746), .B2(new_n959), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT52), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n741), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1071), .A2(KEYINPUT113), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1072), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1061), .B1(new_n1083), .B2(new_n779), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1016), .B2(new_n733), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1057), .A2(new_n1058), .A3(new_n1085), .ZN(G390));
  INV_X1    g0886(.A(KEYINPUT114), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n803), .B1(new_n705), .B2(new_n707), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n913), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n802), .B1(new_n933), .B2(new_n934), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(KEYINPUT114), .A3(new_n913), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n891), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n902), .A2(new_n927), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n925), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n917), .A2(new_n926), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n892), .A2(new_n807), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1095), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1093), .A2(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n850), .A2(G330), .A3(new_n889), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT115), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1103), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(KEYINPUT115), .A3(new_n1101), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n850), .A2(G330), .A3(new_n802), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n891), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1099), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n915), .A2(new_n916), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1113), .B1(new_n807), .B2(new_n803), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1103), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1120), .A2(new_n939), .A3(KEYINPUT116), .A4(new_n851), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT116), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n931), .B1(new_n709), .B2(new_n429), .ZN(new_n1123));
  AND4_X1   g0923(.A1(new_n931), .A2(new_n935), .A3(new_n429), .A4(new_n936), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n652), .B(new_n851), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1118), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1122), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1106), .A2(new_n1110), .A3(new_n1128), .ZN(new_n1129));
  AOI221_X4 g0929(.A(new_n1099), .B1(new_n1096), .B2(new_n1097), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1103), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n681), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n729), .B1(new_n353), .B2(new_n816), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n373), .B1(new_n753), .B2(G125), .ZN(new_n1137));
  INV_X1    g0937(.A(G128), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n746), .C1(new_n834), .C2(new_n958), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n744), .A2(G150), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1140), .A2(KEYINPUT53), .B1(G159), .B2(new_n759), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(KEYINPUT53), .B2(new_n1140), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1139), .B(new_n1142), .C1(new_n972), .C2(new_n740), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT117), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1145), .A2(new_n762), .B1(G137), .B2(new_n750), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT118), .Z(new_n1147));
  OAI221_X1 g0947(.A(new_n373), .B1(new_n758), .B2(new_n813), .C1(new_n823), .C2(new_n208), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n821), .A2(new_n581), .B1(new_n754), .B2(new_n432), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n958), .A2(new_n245), .B1(new_n746), .B2(new_n776), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G87), .A2(new_n966), .B1(new_n740), .B2(G68), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1143), .A2(new_n1147), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1136), .B1(new_n840), .B2(new_n1153), .C1(new_n925), .C2(new_n731), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n1104), .B2(new_n726), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT119), .B1(new_n1135), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT119), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1158), .B(new_n1155), .C1(new_n1129), .C2(new_n1134), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1157), .A2(new_n1159), .ZN(G378));
  NOR3_X1   g0960(.A1(new_n338), .A2(new_n340), .A3(new_n658), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n650), .B2(new_n332), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1161), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n351), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n908), .B2(G330), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n899), .B(new_n1168), .C1(new_n906), .C2(new_n907), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n929), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1168), .B1(new_n898), .B2(new_n899), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n919), .A2(new_n920), .B1(new_n925), .B2(new_n927), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n907), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT40), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n893), .B2(new_n885), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1169), .B(G330), .C1(new_n1175), .C2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1173), .A2(new_n922), .A3(new_n1174), .A4(new_n1178), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1172), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1109), .A2(new_n1101), .A3(new_n1133), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1125), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(KEYINPUT121), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n681), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT121), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT57), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1125), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1186), .B(new_n1187), .C1(new_n1188), .C2(new_n1180), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1184), .A2(new_n1185), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n728), .B1(new_n972), .B2(new_n815), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n590), .A2(new_n762), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n202), .B2(new_n739), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n749), .A2(G107), .B1(new_n750), .B2(G97), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n245), .B2(new_n746), .C1(new_n776), .C2(new_n754), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n975), .A2(new_n1029), .A3(new_n282), .A4(new_n373), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n373), .A2(new_n282), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G50), .B1(new_n281), .B2(new_n282), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1197), .A2(KEYINPUT58), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n747), .A2(G125), .B1(G132), .B2(new_n750), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n749), .A2(G128), .B1(new_n762), .B2(G137), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1145), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1203), .B1(new_n976), .B2(new_n758), .C1(new_n743), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n755), .C2(new_n739), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1200), .B1(KEYINPUT58), .B2(new_n1197), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1191), .B1(new_n1210), .B2(new_n779), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n1169), .B2(new_n731), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT120), .Z(new_n1213));
  INV_X1    g1013(.A(new_n1180), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n727), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1190), .A2(new_n1215), .ZN(G375));
  NAND2_X1  g1016(.A1(new_n1113), .A2(new_n730), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n728), .B1(G68), .B2(new_n815), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n315), .B1(new_n746), .B2(new_n834), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n749), .A2(G137), .B1(new_n762), .B2(G150), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1138), .B2(new_n754), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G50), .C2(new_n759), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G159), .A2(new_n966), .B1(new_n740), .B2(G58), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n823), .C2(new_n1204), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n774), .A2(new_n207), .B1(new_n775), .B2(new_n754), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT122), .Z(new_n1226));
  NAND2_X1  g1026(.A1(new_n740), .A2(G77), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n821), .A2(new_n208), .B1(new_n823), .B2(new_n245), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G283), .B2(new_n749), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n315), .B1(new_n747), .B2(G294), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1229), .A3(new_n1035), .A4(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1224), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1218), .B1(new_n1232), .B2(new_n779), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1120), .A2(new_n727), .B1(new_n1217), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1128), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1006), .B1(new_n1182), .B2(new_n1120), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(G381));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G375), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1190), .A2(KEYINPUT124), .A3(new_n1215), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT123), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1135), .B2(new_n1156), .ZN(new_n1242));
  AOI211_X1 g1042(.A(KEYINPUT123), .B(new_n1155), .C1(new_n1129), .C2(new_n1134), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1239), .A2(new_n1240), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G396), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1050), .A2(new_n1246), .A3(new_n1051), .ZN(new_n1247));
  OR4_X1    g1047(.A1(G384), .A2(new_n1247), .A3(G387), .A4(G390), .ZN(new_n1248));
  OR3_X1    g1048(.A1(new_n1245), .A2(G381), .A3(new_n1248), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  NAND2_X1  g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1247), .ZN(new_n1252));
  INV_X1    g1052(.A(G390), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(G387), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G390), .B(new_n987), .C1(new_n1007), .C2(new_n1018), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1251), .A2(new_n1247), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  INV_X1    g1060(.A(G213), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(G343), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1190), .B(new_n1215), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1006), .A3(new_n1214), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT125), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1183), .A2(new_n1267), .A3(new_n1006), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1215), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1262), .B1(new_n1263), .B2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1133), .A2(new_n681), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1182), .B2(new_n1120), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1125), .A2(KEYINPUT60), .A3(new_n1126), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(G384), .A3(new_n1234), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1276), .B2(new_n1234), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1262), .A2(G2897), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1280), .B(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1259), .B(new_n1260), .C1(new_n1271), .C2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1280), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1262), .B(new_n1285), .C1(new_n1263), .C2(new_n1270), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT63), .B1(new_n1286), .B2(KEYINPUT126), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1271), .A2(new_n1280), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1284), .A2(new_n1287), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1271), .A2(new_n1293), .A3(new_n1280), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1260), .B1(new_n1271), .B2(new_n1282), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1271), .B2(new_n1280), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1292), .B1(new_n1297), .B2(new_n1259), .ZN(G405));
  NAND2_X1  g1098(.A1(new_n1244), .A2(G375), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT127), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1263), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1299), .A2(KEYINPUT127), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1258), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1251), .A2(new_n1255), .A3(new_n1247), .A4(new_n1254), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1285), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1280), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1303), .B(new_n1308), .ZN(G402));
endmodule


