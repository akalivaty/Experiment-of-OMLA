//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n210), .B(new_n214), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G13), .A3(G20), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n207), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g0050(.A1(new_n250), .A2(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n245), .A2(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(KEYINPUT67), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G50), .ZN(new_n255));
  OR2_X1    g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G150), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n208), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n208), .B1(new_n201), .B2(new_n255), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n249), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n263), .A2(KEYINPUT66), .B1(new_n255), .B2(new_n247), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n256), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT9), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n256), .A2(new_n264), .A3(new_n268), .A4(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G222), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G77), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G223), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n273), .B1(new_n274), .B2(new_n271), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n245), .B1(G41), .B2(G45), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n281), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(G226), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G200), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n279), .A2(G190), .A3(new_n285), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n270), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(KEYINPUT68), .A3(new_n288), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT10), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n290), .B(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n279), .A2(new_n297), .A3(new_n285), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n266), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n259), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n247), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n254), .B2(new_n302), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n248), .A2(new_n207), .ZN(new_n305));
  INV_X1    g0105(.A(G68), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT7), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n271), .B2(G20), .ZN(new_n308));
  INV_X1    g0108(.A(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n306), .B1(new_n308), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G58), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n306), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n317), .B2(new_n201), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n257), .A2(G159), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n305), .B1(new_n321), .B2(KEYINPUT16), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT7), .B1(new_n313), .B2(new_n208), .ZN(new_n323));
  AOI211_X1 g0123(.A(new_n307), .B(G20), .C1(new_n310), .C2(new_n312), .ZN(new_n324));
  OAI21_X1  g0124(.A(G68), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n320), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT71), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(KEYINPUT71), .B(new_n328), .C1(new_n315), .C2(new_n320), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n322), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT72), .B(new_n322), .C1(new_n329), .C2(new_n331), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n304), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n271), .A2(new_n272), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n337), .A2(new_n276), .B1(new_n309), .B2(new_n216), .ZN(new_n338));
  INV_X1    g0138(.A(G226), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n275), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n278), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n282), .B1(G232), .B2(new_n284), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT73), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n341), .A2(KEYINPUT73), .A3(new_n342), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n343), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n347), .A2(new_n295), .B1(new_n297), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT18), .B1(new_n336), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n304), .ZN(new_n352));
  INV_X1    g0152(.A(new_n335), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n328), .B1(new_n315), .B2(new_n320), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT71), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n330), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT72), .B1(new_n357), .B2(new_n322), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n352), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n349), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n341), .A2(KEYINPUT73), .A3(new_n342), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT73), .B1(new_n341), .B2(new_n342), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n348), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n352), .C1(new_n353), .C2(new_n358), .ZN(new_n369));
  NAND2_X1  g0169(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n336), .B2(new_n368), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n351), .B(new_n361), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n250), .A2(G77), .A3(new_n252), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G77), .B2(new_n246), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n302), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n260), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n381), .B2(new_n249), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n284), .A2(G244), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n271), .A2(G232), .A3(new_n272), .ZN(new_n385));
  INV_X1    g0185(.A(G107), .ZN(new_n386));
  INV_X1    g0186(.A(G238), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n385), .B1(new_n386), .B2(new_n271), .C1(new_n275), .C2(new_n387), .ZN(new_n388));
  AOI211_X1 g0188(.A(new_n282), .B(new_n384), .C1(new_n388), .C2(new_n278), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n383), .B1(new_n389), .B2(G169), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n389), .A2(new_n297), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(G190), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n382), .C1(new_n362), .C2(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n301), .A2(new_n376), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n398));
  AND3_X1   g0198(.A1(KEYINPUT69), .A2(G33), .A3(G97), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT69), .B1(G33), .B2(G97), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n398), .B(new_n401), .C1(new_n337), .C2(new_n339), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n278), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n282), .B1(G238), .B2(new_n284), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT70), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT13), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n408), .A3(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n403), .A2(KEYINPUT70), .A3(new_n408), .A4(new_n404), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(G169), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT14), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n410), .A2(new_n411), .A3(new_n414), .A4(G169), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(G179), .A3(new_n409), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n247), .A2(new_n306), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT12), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n306), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n274), .B2(new_n260), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n250), .A2(G68), .A3(new_n252), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT11), .B1(new_n421), .B2(new_n249), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n410), .A2(new_n411), .A3(G200), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n366), .B1(new_n405), .B2(KEYINPUT13), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n428), .B2(new_n409), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n417), .A2(new_n426), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n397), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n271), .A2(new_n208), .A3(G87), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT22), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT24), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT23), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n208), .B2(G107), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n386), .A2(KEYINPUT23), .A3(G20), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G116), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n437), .A2(new_n438), .B1(new_n440), .B2(new_n208), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n434), .A2(new_n435), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n435), .B1(new_n434), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n249), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n245), .A2(G33), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n305), .A2(new_n246), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n386), .B1(KEYINPUT81), .B2(KEYINPUT25), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(new_n246), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n247), .A2(KEYINPUT81), .A3(KEYINPUT25), .A4(new_n386), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n446), .A2(G107), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(G250), .A2(G1698), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n219), .B2(G1698), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(new_n271), .B1(G33), .B2(G294), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(KEYINPUT82), .A3(new_n278), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n245), .B(G45), .C1(new_n458), .C2(KEYINPUT5), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT76), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n459), .A2(new_n460), .B1(KEYINPUT5), .B2(new_n458), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(KEYINPUT76), .C1(KEYINPUT5), .C2(new_n458), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n278), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G264), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT82), .ZN(new_n467));
  OAI211_X1 g0267(.A(G1), .B(G13), .C1(new_n309), .C2(new_n458), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n455), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n461), .A2(G274), .A3(new_n468), .A4(new_n464), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n457), .A2(new_n466), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT83), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(G169), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n456), .A2(new_n278), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n466), .A2(new_n474), .A3(new_n470), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n297), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n472), .B1(new_n471), .B2(G169), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n452), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n466), .A2(new_n474), .A3(new_n470), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n479), .A2(G200), .B1(new_n471), .B2(G190), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(new_n444), .A3(new_n451), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n248), .A2(new_n207), .B1(G20), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n208), .C1(G33), .C2(new_n218), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT20), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT78), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n246), .B2(G116), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n247), .A2(KEYINPUT78), .A3(new_n483), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n446), .A2(G116), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n295), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n271), .A2(G264), .A3(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n313), .A2(G303), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n337), .C2(new_n219), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n278), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n465), .A2(G270), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n470), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT21), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n297), .B1(new_n497), .B2(new_n278), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n250), .A2(G116), .A3(new_n445), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n492), .A2(new_n491), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n487), .A2(new_n488), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT20), .B1(new_n484), .B2(new_n486), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n503), .A2(new_n508), .A3(new_n470), .A4(new_n499), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT79), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n499), .A2(new_n470), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(KEYINPUT79), .A3(new_n508), .A4(new_n503), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n494), .A2(new_n500), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT21), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(KEYINPUT80), .B(KEYINPUT21), .C1(new_n494), .C2(new_n500), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n502), .B(new_n514), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n500), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G190), .ZN(new_n522));
  INV_X1    g0322(.A(new_n508), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n500), .A2(G200), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n271), .A2(G244), .A3(G1698), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(new_n439), .C1(new_n337), .C2(new_n387), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n278), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n463), .A2(new_n280), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n217), .B1(new_n462), .B2(G1), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n468), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(G190), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT77), .ZN(new_n535));
  INV_X1    g0335(.A(new_n533), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n529), .B2(new_n278), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT77), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(G190), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n537), .A2(new_n362), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT19), .B1(new_n399), .B2(new_n400), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n542), .A2(new_n208), .B1(new_n216), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n271), .A2(new_n208), .A3(G68), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n260), .B2(new_n218), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n249), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n380), .A2(new_n247), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n446), .A2(G87), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n541), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n537), .A2(G169), .ZN(new_n554));
  AOI211_X1 g0354(.A(G179), .B(new_n536), .C1(new_n529), .C2(new_n278), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n446), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n549), .B(new_n550), .C1(new_n380), .C2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n540), .A2(new_n553), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT6), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n218), .A2(new_n386), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(new_n543), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n386), .A2(KEYINPUT75), .A3(KEYINPUT6), .A4(G97), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT75), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT6), .A2(G97), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n568));
  OAI21_X1  g0368(.A(G107), .B1(new_n323), .B2(new_n324), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n249), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n246), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n446), .B2(G97), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n271), .A2(G244), .A3(new_n272), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n485), .B(new_n575), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n577), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n468), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n465), .A2(G257), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n470), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n295), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n580), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n278), .B1(new_n585), .B2(new_n578), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(new_n297), .A3(new_n470), .A4(new_n582), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n574), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(G200), .B1(new_n581), .B2(new_n583), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n586), .A2(G190), .A3(new_n470), .A4(new_n582), .ZN(new_n590));
  INV_X1    g0390(.A(new_n573), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n570), .B2(new_n249), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n559), .A2(new_n588), .A3(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n432), .A2(new_n482), .A3(new_n527), .A4(new_n594), .ZN(G372));
  NAND2_X1  g0395(.A1(new_n351), .A2(new_n361), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n372), .A2(new_n375), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n427), .A2(new_n429), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n417), .A2(new_n426), .B1(new_n599), .B2(new_n392), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n299), .B1(new_n601), .B2(new_n294), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n556), .A2(new_n558), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT84), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n481), .A2(new_n559), .A3(new_n588), .A4(new_n593), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT80), .B1(new_n501), .B2(KEYINPUT21), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n516), .A2(new_n515), .A3(new_n517), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n511), .A2(new_n513), .B1(new_n501), .B2(KEYINPUT21), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n478), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n604), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT26), .ZN(new_n612));
  INV_X1    g0412(.A(new_n588), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n559), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n540), .A2(new_n553), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n603), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n588), .ZN(new_n617));
  XNOR2_X1  g0417(.A(KEYINPUT85), .B(KEYINPUT26), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n602), .B1(new_n431), .B2(new_n621), .ZN(G369));
  INV_X1    g0422(.A(G330), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n245), .A2(new_n208), .A3(G13), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G213), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n520), .A2(new_n508), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n508), .A2(new_n629), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n608), .A2(new_n609), .A3(new_n525), .A4(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n623), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n452), .A2(new_n629), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n478), .A2(new_n481), .A3(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n452), .B(new_n629), .C1(new_n476), .C2(new_n477), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n629), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n452), .B(new_n639), .C1(new_n476), .C2(new_n477), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n629), .B1(new_n608), .B2(new_n609), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n482), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n638), .A2(new_n643), .ZN(G399));
  INV_X1    g0444(.A(new_n212), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G41), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR4_X1   g0447(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G1), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n205), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT28), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n616), .A2(KEYINPUT26), .A3(new_n588), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n618), .B1(new_n613), .B2(new_n559), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n629), .B1(new_n611), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT29), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI211_X1 g0457(.A(KEYINPUT29), .B(new_n629), .C1(new_n611), .C2(new_n619), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n537), .A2(new_n466), .A3(new_n474), .A4(new_n470), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n503), .A2(new_n499), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n586), .A2(new_n470), .A3(new_n582), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT30), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n537), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n475), .A2(new_n666), .A3(new_n297), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n664), .A2(new_n667), .A3(new_n521), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT87), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n479), .A2(G179), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n500), .A3(new_n663), .A4(new_n666), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT87), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n663), .A2(new_n660), .A3(new_n661), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n671), .B(new_n672), .C1(KEYINPUT30), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT30), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n669), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n639), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n671), .B1(new_n673), .B2(KEYINPUT30), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n673), .A2(KEYINPUT30), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n629), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n482), .A2(new_n527), .A3(new_n594), .A4(new_n639), .ZN(new_n686));
  OAI21_X1  g0486(.A(G330), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n659), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n651), .B1(new_n689), .B2(G1), .ZN(G364));
  NAND2_X1  g0490(.A1(new_n630), .A2(new_n632), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT88), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(G13), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G20), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n245), .B1(new_n696), .B2(G45), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n646), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n693), .A2(new_n694), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n271), .A2(new_n212), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT89), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(G355), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n703), .B2(G355), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(G116), .B2(new_n212), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n313), .A2(new_n212), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT90), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n462), .B2(new_n206), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n240), .A2(new_n462), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n706), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n207), .B1(G20), .B2(new_n295), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n699), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G179), .A2(G200), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n208), .B1(new_n720), .B2(G190), .ZN(new_n721));
  INV_X1    g0521(.A(G294), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n208), .A2(new_n297), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G190), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n362), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(KEYINPUT93), .B(G326), .Z(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n725), .A2(G200), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n723), .B(new_n729), .C1(G322), .C2(new_n730), .ZN(new_n731));
  OR3_X1    g0531(.A1(new_n362), .A2(KEYINPUT91), .A3(G179), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT91), .B1(new_n362), .B2(G179), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n208), .A2(G190), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G283), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n208), .A2(new_n366), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(new_n733), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G303), .ZN(new_n741));
  XOR2_X1   g0541(.A(KEYINPUT33), .B(G317), .Z(new_n742));
  NAND3_X1  g0542(.A1(new_n734), .A2(G179), .A3(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n724), .A2(new_n366), .A3(new_n362), .ZN(new_n745));
  INV_X1    g0545(.A(G311), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n313), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n734), .A2(new_n720), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n744), .B(new_n747), .C1(G329), .C2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n731), .A2(new_n737), .A3(new_n741), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n730), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n316), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n749), .A2(G159), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n727), .A2(new_n255), .B1(new_n754), .B2(KEYINPUT32), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n753), .B(new_n755), .C1(KEYINPUT32), .C2(new_n754), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n740), .A2(G87), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n271), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT92), .ZN(new_n759));
  INV_X1    g0559(.A(new_n721), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G97), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n761), .B1(new_n306), .B2(new_n743), .C1(new_n274), .C2(new_n745), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(G107), .B2(new_n736), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n756), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n758), .A2(KEYINPUT92), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n751), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n719), .B1(new_n766), .B2(new_n716), .ZN(new_n767));
  INV_X1    g0567(.A(new_n715), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n691), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n701), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(G396));
  OAI21_X1  g0571(.A(new_n395), .B1(new_n382), .B2(new_n639), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n393), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n392), .A2(new_n639), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(new_n621), .B2(new_n629), .ZN(new_n776));
  INV_X1    g0576(.A(new_n775), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n620), .A2(new_n639), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n699), .B1(new_n779), .B2(new_n687), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n687), .B2(new_n779), .ZN(new_n781));
  INV_X1    g0581(.A(new_n745), .ZN(new_n782));
  INV_X1    g0582(.A(new_n743), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G159), .A2(new_n782), .B1(new_n783), .B2(G150), .ZN(new_n784));
  INV_X1    g0584(.A(G137), .ZN(new_n785));
  INV_X1    g0585(.A(G143), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n784), .B1(new_n785), .B2(new_n727), .C1(new_n786), .C2(new_n752), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n736), .A2(G68), .ZN(new_n790));
  INV_X1    g0590(.A(G132), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n271), .B1(new_n721), .B2(new_n316), .C1(new_n791), .C2(new_n748), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(G50), .B2(new_n740), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n787), .A2(new_n788), .ZN(new_n795));
  INV_X1    g0595(.A(G303), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n761), .B1(new_n752), .B2(new_n722), .C1(new_n796), .C2(new_n727), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n736), .A2(G87), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n740), .A2(G107), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n271), .B1(new_n782), .B2(G116), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n783), .A2(G283), .B1(new_n749), .B2(G311), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n794), .A2(new_n795), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n716), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n716), .A2(new_n713), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n700), .B1(new_n274), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n804), .B(new_n806), .C1(new_n777), .C2(new_n714), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n781), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G384));
  NAND4_X1  g0609(.A1(new_n482), .A2(new_n527), .A3(new_n594), .A4(new_n639), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n682), .A2(new_n677), .ZN(new_n811));
  OAI211_X1 g0611(.A(KEYINPUT31), .B(new_n629), .C1(new_n680), .C2(new_n681), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n426), .A2(new_n629), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT94), .Z(new_n815));
  OR2_X1    g0615(.A1(new_n430), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n430), .A2(new_n815), .ZN(new_n817));
  AND4_X1   g0617(.A1(new_n777), .A2(new_n813), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n359), .A2(new_n349), .ZN(new_n819));
  INV_X1    g0619(.A(new_n627), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n359), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT37), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n819), .A2(new_n821), .A3(new_n822), .A4(new_n369), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n322), .A2(new_n354), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n352), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n349), .B2(new_n820), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n369), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n627), .B1(new_n824), .B2(new_n352), .ZN(new_n830));
  AOI22_X1  g0630(.A1(KEYINPUT95), .A2(new_n829), .B1(new_n376), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT95), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n823), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT38), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n829), .A2(KEYINPUT95), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n376), .A2(new_n830), .ZN(new_n836));
  AND4_X1   g0636(.A1(KEYINPUT38), .A2(new_n835), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n818), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(KEYINPUT98), .B(KEYINPUT40), .Z(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT38), .A4(new_n833), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT97), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n831), .A2(KEYINPUT97), .A3(KEYINPUT38), .A4(new_n833), .ZN(new_n845));
  INV_X1    g0645(.A(new_n821), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n376), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n819), .A2(new_n821), .A3(new_n369), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n823), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n844), .A2(new_n845), .A3(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n818), .A2(KEYINPUT40), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n841), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n432), .A2(new_n813), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT99), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n623), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n862), .A2(KEYINPUT100), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n862), .A2(KEYINPUT100), .B1(new_n858), .B2(new_n860), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n417), .A2(new_n426), .A3(new_n639), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT39), .B1(new_n851), .B2(new_n852), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n844), .A2(new_n868), .A3(new_n845), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT39), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n835), .A2(new_n836), .A3(new_n833), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n852), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n872), .B2(new_n842), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n867), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n816), .A2(new_n817), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n774), .B2(new_n778), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n834), .B2(new_n837), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n597), .A2(new_n820), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(KEYINPUT96), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT96), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n430), .A2(new_n815), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n430), .A2(new_n815), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n629), .B(new_n775), .C1(new_n611), .C2(new_n619), .ZN(new_n885));
  INV_X1    g0685(.A(new_n774), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n872), .B2(new_n842), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n881), .B1(new_n888), .B2(new_n878), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n874), .A2(new_n880), .A3(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n397), .B(new_n430), .C1(new_n657), .C2(new_n658), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n602), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n890), .B(new_n892), .Z(new_n893));
  OR2_X1    g0693(.A1(new_n865), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n865), .A2(new_n893), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n894), .B(new_n895), .C1(new_n245), .C2(new_n696), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(G116), .A3(new_n209), .A4(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT36), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n205), .A2(new_n274), .A3(new_n317), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n306), .A2(G50), .ZN(new_n902));
  OAI211_X1 g0702(.A(G1), .B(new_n695), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n896), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT101), .Z(G367));
  INV_X1    g0705(.A(new_n604), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n552), .A2(new_n629), .ZN(new_n907));
  MUX2_X1   g0707(.A(new_n906), .B(new_n616), .S(new_n907), .Z(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n715), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n721), .A2(new_n306), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n271), .B1(new_n748), .B2(new_n785), .C1(new_n727), .C2(new_n786), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n910), .B(new_n911), .C1(G150), .C2(new_n730), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n735), .A2(new_n274), .ZN(new_n913));
  INV_X1    g0713(.A(G159), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n745), .A2(new_n255), .B1(new_n743), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT108), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n740), .A2(G58), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n912), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n739), .A2(new_n483), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT46), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n727), .A2(new_n746), .B1(new_n721), .B2(new_n386), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(G303), .B2(new_n730), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n736), .A2(G97), .ZN(new_n925));
  INV_X1    g0725(.A(G317), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n743), .A2(new_n722), .B1(new_n748), .B2(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n271), .B(new_n927), .C1(G283), .C2(new_n782), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n920), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT47), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n716), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n232), .A2(new_n708), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n933), .B(new_n717), .C1(new_n212), .C2(new_n380), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n909), .A2(new_n932), .A3(new_n699), .A4(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT102), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n574), .A2(new_n629), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n588), .A2(new_n593), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n574), .A2(new_n584), .A3(new_n587), .A4(new_n629), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n938), .A2(new_n936), .A3(new_n939), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n944));
  NAND3_X1  g0744(.A1(new_n643), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n944), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n938), .A2(new_n939), .A3(new_n936), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n940), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n520), .A2(new_n478), .A3(new_n481), .A4(new_n639), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n640), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n946), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT44), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT44), .B1(new_n948), .B2(new_n950), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n945), .B(new_n951), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n638), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT105), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n945), .A2(new_n951), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT44), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n643), .B2(new_n943), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n957), .A2(new_n961), .A3(new_n962), .A4(new_n638), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n638), .B1(new_n957), .B2(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n605), .A2(new_n610), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n654), .A3(new_n906), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n639), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT29), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n520), .A2(new_n639), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n635), .A2(new_n970), .A3(new_n636), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n694), .A2(new_n949), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n949), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n633), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n620), .A2(new_n656), .A3(new_n639), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n969), .A2(new_n975), .A3(new_n976), .A4(new_n687), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n965), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n964), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT106), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT106), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n964), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n688), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n646), .B(KEYINPUT41), .Z(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT107), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n964), .A2(new_n978), .A3(new_n981), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n981), .B1(new_n964), .B2(new_n978), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n689), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT107), .ZN(new_n989));
  INV_X1    g0789(.A(new_n984), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n698), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n948), .A2(new_n478), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n629), .B1(new_n993), .B2(new_n588), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n482), .B(new_n642), .C1(new_n947), .C2(new_n940), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT43), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n994), .A2(new_n996), .B1(new_n997), .B2(new_n908), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n908), .A2(new_n997), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n998), .B(new_n999), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n638), .A2(new_n948), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1000), .B1(KEYINPUT103), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(KEYINPUT103), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n935), .B1(new_n992), .B2(new_n1005), .ZN(G387));
  NAND3_X1  g0806(.A1(new_n635), .A2(new_n636), .A3(new_n715), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n702), .A2(new_n648), .B1(G107), .B2(new_n212), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n236), .A2(G45), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n648), .B(new_n462), .C1(new_n306), .C2(new_n274), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT50), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n259), .B2(G50), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n302), .A2(KEYINPUT50), .A3(new_n255), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n709), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1008), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n699), .B1(new_n1016), .B2(new_n718), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n728), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n271), .B1(new_n1018), .B2(new_n749), .ZN(new_n1019));
  INV_X1    g0819(.A(G283), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n739), .A2(new_n722), .B1(new_n1020), .B2(new_n721), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G303), .A2(new_n782), .B1(new_n783), .B2(G311), .ZN(new_n1022));
  XOR2_X1   g0822(.A(KEYINPUT109), .B(G322), .Z(new_n1023));
  OAI221_X1 g0823(.A(new_n1022), .B1(new_n926), .B2(new_n752), .C1(new_n727), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1019), .B1(new_n483), .B2(new_n735), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n721), .A2(new_n380), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n752), .B2(new_n255), .C1(new_n914), .C2(new_n727), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G68), .A2(new_n782), .B1(new_n783), .B2(new_n302), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n740), .A2(G77), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n313), .B1(new_n749), .B2(G150), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n925), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1029), .A2(new_n1030), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT110), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n716), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n1037), .B2(KEYINPUT110), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1017), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1007), .A2(new_n1041), .B1(new_n975), .B2(new_n698), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n689), .A2(new_n975), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n646), .A3(new_n977), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  NAND2_X1  g0847(.A1(new_n954), .A2(new_n955), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT112), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n964), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n647), .B1(new_n1050), .B2(new_n977), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n986), .B2(new_n987), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n698), .A3(new_n964), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n708), .A2(new_n243), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n718), .B1(G97), .B2(new_n645), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n700), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n798), .B1(new_n306), .B2(new_n739), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n721), .A2(new_n274), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n271), .B1(new_n745), .B2(new_n259), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n743), .A2(new_n255), .B1(new_n748), .B2(new_n786), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G150), .A2(new_n726), .B1(new_n730), .B2(G159), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT51), .Z(new_n1063));
  AOI22_X1  g0863(.A1(G311), .A2(new_n730), .B1(new_n726), .B2(G317), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT52), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n1020), .A2(new_n739), .B1(new_n735), .B2(new_n386), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1023), .A2(new_n748), .B1(new_n743), .B2(new_n796), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n313), .B1(new_n745), .B2(new_n722), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n721), .A2(new_n483), .ZN(new_n1069));
  NOR4_X1   g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1061), .A2(new_n1063), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1056), .B1(new_n1039), .B2(new_n1071), .C1(new_n943), .C2(new_n768), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1052), .A2(new_n1053), .A3(new_n1072), .ZN(G390));
  OAI21_X1  g0873(.A(KEYINPUT39), .B1(new_n834), .B2(new_n837), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n844), .A2(new_n868), .A3(new_n845), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n887), .A2(new_n866), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n886), .B1(new_n655), .B2(new_n773), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(new_n875), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n866), .B(KEYINPUT113), .Z(new_n1080));
  NAND3_X1  g0880(.A1(new_n854), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n813), .A2(G330), .A3(new_n777), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1083), .A2(new_n875), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n676), .A2(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n623), .B1(new_n1086), .B2(new_n810), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n884), .A2(new_n1087), .A3(new_n777), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1077), .A2(new_n1088), .A3(new_n1081), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n778), .A2(new_n774), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1087), .A2(new_n777), .B1(new_n817), .B2(new_n816), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1083), .A2(new_n875), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1093), .A3(new_n1078), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n397), .A2(G330), .A3(new_n430), .A4(new_n813), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n891), .A2(new_n602), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1085), .A2(new_n1089), .A3(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1095), .A2(new_n1098), .A3(KEYINPUT114), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT114), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1077), .A2(new_n1088), .A3(new_n1081), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1084), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n646), .B(new_n1101), .C1(new_n1105), .C2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1074), .A2(new_n1075), .A3(new_n713), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n805), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n699), .B1(new_n1112), .B2(new_n302), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n727), .A2(new_n1020), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1058), .B(new_n1114), .C1(G116), .C2(new_n730), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n745), .A2(new_n218), .B1(new_n743), .B2(new_n386), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n271), .B(new_n1116), .C1(G294), .C2(new_n749), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1115), .A2(new_n757), .A3(new_n790), .A4(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n752), .A2(new_n791), .B1(new_n721), .B2(new_n914), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G128), .B2(new_n726), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n736), .A2(G50), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n313), .B1(new_n782), .B2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n783), .A2(G137), .B1(new_n749), .B2(G125), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1120), .A2(new_n1121), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G150), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n739), .A2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1118), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1113), .B1(new_n1131), .B2(new_n716), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT116), .Z(new_n1133));
  AOI22_X1  g0933(.A1(new_n1109), .A2(new_n698), .B1(new_n1111), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1110), .A2(new_n1134), .ZN(G378));
  NAND2_X1  g0935(.A1(new_n266), .A2(new_n820), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT55), .Z(new_n1137));
  NAND2_X1  g0937(.A1(new_n301), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1137), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n294), .A2(new_n300), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1139), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AND4_X1   g0946(.A1(G330), .A2(new_n841), .A3(new_n856), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n623), .B1(new_n838), .B2(new_n840), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1148), .B2(new_n856), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n890), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n856), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n884), .A2(new_n777), .A3(new_n813), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n872), .B2(new_n842), .ZN(new_n1153));
  OAI21_X1  g0953(.A(G330), .B1(new_n1153), .B2(new_n839), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1145), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n889), .A2(new_n880), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n841), .A2(new_n856), .A3(G330), .A4(new_n1146), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n874), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1145), .A2(new_n713), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n699), .B1(new_n1112), .B2(G50), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n727), .A2(new_n483), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n910), .B(new_n1162), .C1(G107), .C2(new_n730), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n736), .A2(G58), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT118), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n458), .B(new_n313), .C1(new_n745), .C2(new_n380), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n743), .A2(new_n218), .B1(new_n748), .B2(new_n1020), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1163), .A2(new_n1034), .A3(new_n1165), .A4(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT58), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(G33), .A2(G41), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT117), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1172), .B(new_n255), .C1(G41), .C2(new_n271), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n745), .A2(new_n785), .B1(new_n743), .B2(new_n791), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G125), .B2(new_n726), .ZN(new_n1175));
  OR3_X1    g0975(.A1(new_n739), .A2(KEYINPUT119), .A3(new_n1122), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT119), .B1(new_n739), .B2(new_n1122), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n730), .A2(G128), .B1(G150), .B2(new_n760), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1172), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT120), .B(G124), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1181), .B1(new_n748), .B2(new_n1182), .C1(new_n914), .C2(new_n735), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT121), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1170), .B(new_n1173), .C1(new_n1180), .C2(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT122), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1039), .B1(new_n1187), .B2(KEYINPUT122), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1161), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1159), .A2(new_n698), .B1(new_n1160), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1101), .A2(new_n1098), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1159), .A2(new_n1192), .A3(KEYINPUT57), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n646), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT57), .B1(new_n1159), .B2(new_n1192), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1191), .B1(new_n1194), .B2(new_n1195), .ZN(G375));
  NAND2_X1  g0996(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1104), .A2(new_n990), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n700), .B1(new_n306), .B2(new_n805), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n783), .A2(new_n1123), .B1(new_n749), .B2(G128), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1200), .B(new_n271), .C1(new_n1127), .C2(new_n745), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G132), .A2(new_n726), .B1(new_n730), .B2(G137), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n255), .B2(new_n721), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(G159), .C2(new_n740), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n271), .B1(new_n749), .B2(G303), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n386), .B2(new_n745), .C1(new_n483), .C2(new_n743), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n913), .B(new_n1206), .C1(G97), .C2(new_n740), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1031), .B1(new_n752), .B2(new_n1020), .C1(new_n722), .C2(new_n727), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1204), .A2(new_n1165), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1199), .B1(new_n1039), .B2(new_n1210), .C1(new_n884), .C2(new_n714), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n1096), .B2(new_n697), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1198), .A2(new_n1213), .ZN(G381));
  INV_X1    g1014(.A(G390), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1213), .A4(new_n1198), .ZN(new_n1217));
  OR4_X1    g1017(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1217), .ZN(G407));
  NOR3_X1   g1018(.A1(new_n1147), .A2(new_n890), .A3(new_n1149), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1157), .A2(new_n1155), .B1(new_n1156), .B2(new_n874), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n698), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1160), .A2(new_n1190), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1159), .A2(new_n1192), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT57), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n647), .B1(new_n1227), .B2(new_n1192), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1223), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(G378), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n628), .A2(G213), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(G407), .A2(G213), .A3(new_n1233), .ZN(G409));
  OAI211_X1 g1034(.A(G378), .B(new_n1191), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1159), .A2(new_n1192), .A3(new_n990), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1191), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1230), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT60), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n646), .B1(new_n1240), .B2(new_n1197), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1240), .B2(new_n1197), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n808), .B1(new_n1242), .B2(new_n1212), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1240), .A2(new_n1197), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G384), .B(new_n1213), .C1(new_n1244), .C2(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1239), .A2(new_n1231), .A3(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT124), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT63), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1239), .A2(KEYINPUT124), .A3(new_n1231), .A4(new_n1247), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(new_n1215), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(G393), .B(new_n770), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G390), .B(new_n935), .C1(new_n992), .C2(new_n1005), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1254), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n989), .B1(new_n988), .B2(new_n990), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n697), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1003), .B(new_n1004), .Z(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1265), .A2(KEYINPUT125), .A3(new_n935), .A4(G390), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1260), .A2(new_n1266), .A3(new_n1254), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1267), .A2(KEYINPUT126), .A3(new_n1255), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1267), .B2(new_n1255), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1258), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1239), .A2(new_n1231), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1232), .A2(G2897), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1243), .A2(new_n1245), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1232), .B(new_n1246), .C1(new_n1235), .C2(new_n1238), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT63), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1253), .A2(new_n1270), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1258), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1267), .A2(new_n1255), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1267), .A2(KEYINPUT126), .A3(new_n1255), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1280), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1191), .B2(new_n1236), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1229), .B2(G378), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1275), .B1(new_n1287), .B2(new_n1232), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1249), .B1(new_n1290), .B2(KEYINPUT62), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1288), .B(new_n1289), .C1(new_n1277), .C2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT62), .B1(new_n1252), .B2(new_n1290), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1285), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1279), .A2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1230), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1235), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1247), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1235), .A3(new_n1246), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1285), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1270), .A2(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1301), .A2(new_n1303), .ZN(G402));
endmodule


