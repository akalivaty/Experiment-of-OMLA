

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U556 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  NOR2_X1 U557 ( .A1(n533), .A2(n532), .ZN(G164) );
  NAND2_X1 U558 ( .A1(n658), .A2(n969), .ZN(n651) );
  AND2_X1 U559 ( .A1(n637), .A2(n636), .ZN(n658) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n617) );
  BUF_X1 U561 ( .A(n593), .Z(n594) );
  INV_X1 U562 ( .A(G2105), .ZN(n529) );
  NOR2_X4 U563 ( .A1(G651), .A2(G543), .ZN(n643) );
  AND2_X2 U564 ( .A1(n633), .A2(n632), .ZN(n678) );
  NAND2_X1 U565 ( .A1(n879), .A2(G138), .ZN(n528) );
  NOR2_X1 U566 ( .A1(n721), .A2(n733), .ZN(n523) );
  INV_X1 U567 ( .A(KEYINPUT105), .ZN(n694) );
  XNOR2_X1 U568 ( .A(n695), .B(n694), .ZN(n701) );
  AND2_X1 U569 ( .A1(n617), .A2(n616), .ZN(n632) );
  NAND2_X1 U570 ( .A1(n803), .A2(G66), .ZN(n645) );
  XNOR2_X1 U571 ( .A(n623), .B(KEYINPUT13), .ZN(n624) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n524) );
  XNOR2_X1 U573 ( .A(KEYINPUT15), .B(KEYINPUT75), .ZN(n649) );
  INV_X1 U574 ( .A(KEYINPUT1), .ZN(n540) );
  XNOR2_X1 U575 ( .A(n625), .B(n624), .ZN(n628) );
  NOR2_X1 U576 ( .A1(n628), .A2(n627), .ZN(n630) );
  XNOR2_X1 U577 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n767) );
  NAND2_X1 U578 ( .A1(n630), .A2(n629), .ZN(n977) );
  XNOR2_X2 U579 ( .A(n525), .B(n524), .ZN(n879) );
  AND2_X1 U580 ( .A1(G2104), .A2(n529), .ZN(n526) );
  XNOR2_X1 U581 ( .A(n526), .B(KEYINPUT64), .ZN(n593) );
  NAND2_X1 U582 ( .A1(G102), .A2(n593), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n533) );
  NOR2_X2 U584 ( .A1(G2104), .A2(n529), .ZN(n874) );
  NAND2_X1 U585 ( .A1(G126), .A2(n874), .ZN(n531) );
  AND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n875) );
  NAND2_X1 U587 ( .A1(G114), .A2(n875), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .ZN(n638) );
  AND2_X1 U590 ( .A1(n638), .A2(G651), .ZN(n802) );
  NAND2_X1 U591 ( .A1(G72), .A2(n802), .ZN(n535) );
  NAND2_X1 U592 ( .A1(G85), .A2(n643), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n535), .A2(n534), .ZN(n538) );
  INV_X1 U594 ( .A(n638), .ZN(n574) );
  NOR2_X2 U595 ( .A1(G651), .A2(n574), .ZN(n806) );
  NAND2_X1 U596 ( .A1(G47), .A2(n806), .ZN(n536) );
  XOR2_X1 U597 ( .A(KEYINPUT66), .B(n536), .Z(n537) );
  NOR2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n543) );
  INV_X1 U599 ( .A(G651), .ZN(n539) );
  NOR2_X1 U600 ( .A1(G543), .A2(n539), .ZN(n541) );
  XNOR2_X2 U601 ( .A(n541), .B(n540), .ZN(n803) );
  NAND2_X1 U602 ( .A1(n803), .A2(G60), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U604 ( .A(KEYINPUT67), .B(n544), .Z(G290) );
  NAND2_X1 U605 ( .A1(G64), .A2(n803), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G52), .A2(n806), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G77), .A2(n802), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G90), .A2(n643), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U612 ( .A1(n551), .A2(n550), .ZN(G171) );
  INV_X1 U613 ( .A(G171), .ZN(G301) );
  NAND2_X1 U614 ( .A1(G63), .A2(n803), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G51), .A2(n806), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U617 ( .A(KEYINPUT6), .B(n554), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n643), .A2(G89), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G76), .A2(n802), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U622 ( .A(n558), .B(KEYINPUT5), .Z(n559) );
  NOR2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT7), .B(n561), .Z(n562) );
  XNOR2_X1 U625 ( .A(KEYINPUT76), .B(n562), .ZN(G168) );
  XOR2_X1 U626 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U627 ( .A1(G62), .A2(n803), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G50), .A2(n806), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT81), .B(n565), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G75), .A2(n802), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G88), .A2(n643), .ZN(n566) );
  AND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(G303) );
  NAND2_X1 U635 ( .A1(G49), .A2(n806), .ZN(n571) );
  NAND2_X1 U636 ( .A1(G74), .A2(G651), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT79), .B(n572), .Z(n573) );
  NOR2_X1 U639 ( .A1(n803), .A2(n573), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(G87), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(G288) );
  NAND2_X1 U642 ( .A1(G86), .A2(n643), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G61), .A2(n803), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT80), .B(n579), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n802), .A2(G73), .ZN(n580) );
  XOR2_X1 U647 ( .A(KEYINPUT2), .B(n580), .Z(n581) );
  NOR2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n806), .A2(G48), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(G305) );
  NAND2_X1 U651 ( .A1(n593), .A2(G101), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n586), .B(KEYINPUT65), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n587), .B(KEYINPUT23), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G125), .A2(n874), .ZN(n588) );
  AND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n633) );
  NAND2_X1 U656 ( .A1(G137), .A2(n879), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G113), .A2(n875), .ZN(n590) );
  AND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n769) );
  AND2_X1 U659 ( .A1(n769), .A2(G40), .ZN(n616) );
  NAND2_X1 U660 ( .A1(n633), .A2(n616), .ZN(n592) );
  NOR2_X1 U661 ( .A1(n617), .A2(n592), .ZN(n763) );
  XNOR2_X1 U662 ( .A(KEYINPUT94), .B(n763), .ZN(n613) );
  XOR2_X1 U663 ( .A(KEYINPUT38), .B(KEYINPUT93), .Z(n596) );
  NAND2_X1 U664 ( .A1(G105), .A2(n594), .ZN(n595) );
  XNOR2_X1 U665 ( .A(n596), .B(n595), .ZN(n603) );
  NAND2_X1 U666 ( .A1(G141), .A2(n879), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G129), .A2(n874), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n875), .A2(G117), .ZN(n599) );
  XOR2_X1 U670 ( .A(KEYINPUT92), .B(n599), .Z(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n860) );
  NAND2_X1 U673 ( .A1(G1996), .A2(n860), .ZN(n612) );
  NAND2_X1 U674 ( .A1(n875), .A2(G107), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G95), .A2(n594), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U677 ( .A1(G119), .A2(n874), .ZN(n606) );
  XNOR2_X1 U678 ( .A(KEYINPUT91), .B(n606), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n879), .A2(G131), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n856) );
  NAND2_X1 U682 ( .A1(G1991), .A2(n856), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n1009) );
  NAND2_X1 U684 ( .A1(n613), .A2(n1009), .ZN(n753) );
  XNOR2_X1 U685 ( .A(G1986), .B(G290), .ZN(n986) );
  NAND2_X1 U686 ( .A1(n986), .A2(n763), .ZN(n614) );
  XOR2_X1 U687 ( .A(KEYINPUT87), .B(n614), .Z(n615) );
  NAND2_X1 U688 ( .A1(n753), .A2(n615), .ZN(n737) );
  NAND2_X1 U689 ( .A1(n633), .A2(n632), .ZN(n696) );
  AND2_X1 U690 ( .A1(n696), .A2(G1341), .ZN(n631) );
  XOR2_X1 U691 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n619) );
  NAND2_X1 U692 ( .A1(G81), .A2(n643), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n620), .B(KEYINPUT70), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G68), .A2(n802), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n625) );
  INV_X1 U697 ( .A(KEYINPUT72), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n803), .A2(G56), .ZN(n626) );
  XOR2_X1 U699 ( .A(KEYINPUT14), .B(n626), .Z(n627) );
  NAND2_X1 U700 ( .A1(n806), .A2(G43), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n631), .A2(n977), .ZN(n637) );
  NAND2_X1 U702 ( .A1(n678), .A2(G1996), .ZN(n635) );
  XOR2_X1 U703 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n634) );
  XNOR2_X1 U704 ( .A(n635), .B(n634), .ZN(n636) );
  AND2_X1 U705 ( .A1(G79), .A2(G651), .ZN(n639) );
  NAND2_X1 U706 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U707 ( .A(KEYINPUT74), .B(n640), .Z(n642) );
  AND2_X1 U708 ( .A1(G54), .A2(n806), .ZN(n641) );
  NOR2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n648) );
  NAND2_X1 U710 ( .A1(G92), .A2(n643), .ZN(n644) );
  NAND2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n646), .B(KEYINPUT73), .ZN(n647) );
  AND2_X1 U713 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X2 U714 ( .A(n650), .B(n649), .ZN(n969) );
  XNOR2_X1 U715 ( .A(KEYINPUT98), .B(n651), .ZN(n656) );
  NAND2_X1 U716 ( .A1(G1348), .A2(n696), .ZN(n653) );
  NAND2_X1 U717 ( .A1(G2067), .A2(n678), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U719 ( .A(KEYINPUT99), .B(n654), .Z(n655) );
  AND2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U721 ( .A(n657), .B(KEYINPUT100), .ZN(n660) );
  NOR2_X1 U722 ( .A1(n969), .A2(n658), .ZN(n659) );
  NOR2_X1 U723 ( .A1(n660), .A2(n659), .ZN(n671) );
  NAND2_X1 U724 ( .A1(G65), .A2(n803), .ZN(n662) );
  NAND2_X1 U725 ( .A1(G53), .A2(n806), .ZN(n661) );
  NAND2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U727 ( .A1(G78), .A2(n802), .ZN(n664) );
  NAND2_X1 U728 ( .A1(G91), .A2(n643), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n984) );
  NAND2_X1 U731 ( .A1(n678), .A2(G2072), .ZN(n667) );
  XNOR2_X1 U732 ( .A(n667), .B(KEYINPUT27), .ZN(n669) );
  XOR2_X1 U733 ( .A(KEYINPUT96), .B(G1956), .Z(n942) );
  NOR2_X1 U734 ( .A1(n678), .A2(n942), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n673) );
  AND2_X1 U736 ( .A1(n984), .A2(n673), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT101), .ZN(n676) );
  NOR2_X1 U739 ( .A1(n984), .A2(n673), .ZN(n674) );
  XOR2_X1 U740 ( .A(KEYINPUT28), .B(n674), .Z(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n677), .B(KEYINPUT29), .ZN(n682) );
  XOR2_X1 U743 ( .A(KEYINPUT25), .B(G2078), .Z(n927) );
  NOR2_X1 U744 ( .A1(n927), .A2(n696), .ZN(n680) );
  XOR2_X1 U745 ( .A(KEYINPUT95), .B(G1961), .Z(n951) );
  NOR2_X1 U746 ( .A1(n678), .A2(n951), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n687) );
  NOR2_X1 U748 ( .A1(G301), .A2(n687), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n692) );
  NOR2_X1 U750 ( .A1(G2084), .A2(n696), .ZN(n708) );
  NAND2_X1 U751 ( .A1(G8), .A2(n696), .ZN(n733) );
  NOR2_X1 U752 ( .A1(G1966), .A2(n733), .ZN(n706) );
  NOR2_X1 U753 ( .A1(n708), .A2(n706), .ZN(n683) );
  NAND2_X1 U754 ( .A1(G8), .A2(n683), .ZN(n684) );
  XNOR2_X1 U755 ( .A(KEYINPUT30), .B(n684), .ZN(n685) );
  NOR2_X1 U756 ( .A1(G168), .A2(n685), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT102), .ZN(n689) );
  AND2_X1 U758 ( .A1(n687), .A2(G301), .ZN(n688) );
  NOR2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U760 ( .A(n690), .B(KEYINPUT31), .ZN(n691) );
  NOR2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U762 ( .A(n693), .B(KEYINPUT103), .ZN(n704) );
  NAND2_X1 U763 ( .A1(n704), .A2(G286), .ZN(n695) );
  NOR2_X1 U764 ( .A1(G1971), .A2(n733), .ZN(n698) );
  NOR2_X1 U765 ( .A1(G2090), .A2(n696), .ZN(n697) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G303), .A2(n699), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n702), .A2(G8), .ZN(n703) );
  XNOR2_X1 U770 ( .A(n703), .B(KEYINPUT32), .ZN(n712) );
  INV_X1 U771 ( .A(n704), .ZN(n705) );
  NOR2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U773 ( .A(n707), .B(KEYINPUT104), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n708), .A2(G8), .ZN(n709) );
  NAND2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n720) );
  NOR2_X1 U777 ( .A1(G2090), .A2(G303), .ZN(n713) );
  XNOR2_X1 U778 ( .A(n713), .B(KEYINPUT106), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n714), .A2(G8), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n720), .A2(n715), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n716), .A2(n733), .ZN(n730) );
  NOR2_X1 U782 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NOR2_X1 U783 ( .A1(G1971), .A2(G303), .ZN(n991) );
  NOR2_X1 U784 ( .A1(n965), .A2(n991), .ZN(n718) );
  INV_X1 U785 ( .A(KEYINPUT33), .ZN(n717) );
  AND2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n728) );
  NAND2_X1 U788 ( .A1(G1976), .A2(G288), .ZN(n967) );
  INV_X1 U789 ( .A(n967), .ZN(n721) );
  NOR2_X1 U790 ( .A1(KEYINPUT33), .A2(n523), .ZN(n726) );
  XOR2_X1 U791 ( .A(G1981), .B(G305), .Z(n972) );
  INV_X1 U792 ( .A(n972), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n965), .A2(KEYINPUT33), .ZN(n722) );
  NOR2_X1 U794 ( .A1(n722), .A2(n733), .ZN(n723) );
  OR2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U796 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U797 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n735) );
  NOR2_X1 U799 ( .A1(G1981), .A2(G305), .ZN(n731) );
  XOR2_X1 U800 ( .A(n731), .B(KEYINPUT24), .Z(n732) );
  NOR2_X1 U801 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U802 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U803 ( .A1(n737), .A2(n736), .ZN(n750) );
  XNOR2_X1 U804 ( .A(G2067), .B(KEYINPUT37), .ZN(n738) );
  XOR2_X1 U805 ( .A(n738), .B(KEYINPUT88), .Z(n760) );
  NAND2_X1 U806 ( .A1(n879), .A2(G140), .ZN(n740) );
  NAND2_X1 U807 ( .A1(G104), .A2(n594), .ZN(n739) );
  NAND2_X1 U808 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U809 ( .A(KEYINPUT34), .B(n741), .ZN(n747) );
  NAND2_X1 U810 ( .A1(G128), .A2(n874), .ZN(n743) );
  NAND2_X1 U811 ( .A1(G116), .A2(n875), .ZN(n742) );
  NAND2_X1 U812 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U813 ( .A(KEYINPUT35), .B(n744), .ZN(n745) );
  XNOR2_X1 U814 ( .A(KEYINPUT89), .B(n745), .ZN(n746) );
  NOR2_X1 U815 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U816 ( .A(n748), .B(KEYINPUT36), .ZN(n749) );
  XOR2_X1 U817 ( .A(n749), .B(KEYINPUT90), .Z(n888) );
  AND2_X1 U818 ( .A1(n760), .A2(n888), .ZN(n1021) );
  NAND2_X1 U819 ( .A1(n763), .A2(n1021), .ZN(n759) );
  NAND2_X1 U820 ( .A1(n750), .A2(n759), .ZN(n766) );
  NOR2_X1 U821 ( .A1(G1986), .A2(G290), .ZN(n751) );
  NOR2_X1 U822 ( .A1(G1991), .A2(n856), .ZN(n1002) );
  NOR2_X1 U823 ( .A1(n751), .A2(n1002), .ZN(n752) );
  XNOR2_X1 U824 ( .A(KEYINPUT107), .B(n752), .ZN(n754) );
  NAND2_X1 U825 ( .A1(n754), .A2(n753), .ZN(n755) );
  OR2_X1 U826 ( .A1(n860), .A2(G1996), .ZN(n1003) );
  NAND2_X1 U827 ( .A1(n755), .A2(n1003), .ZN(n757) );
  XOR2_X1 U828 ( .A(KEYINPUT108), .B(KEYINPUT39), .Z(n756) );
  XNOR2_X1 U829 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U830 ( .A1(n759), .A2(n758), .ZN(n762) );
  NOR2_X1 U831 ( .A1(n888), .A2(n760), .ZN(n761) );
  XNOR2_X1 U832 ( .A(n761), .B(KEYINPUT109), .ZN(n1018) );
  NAND2_X1 U833 ( .A1(n762), .A2(n1018), .ZN(n764) );
  NAND2_X1 U834 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U835 ( .A1(n766), .A2(n765), .ZN(n768) );
  XNOR2_X1 U836 ( .A(n768), .B(n767), .ZN(G329) );
  AND2_X1 U837 ( .A1(n633), .A2(n769), .ZN(G160) );
  XOR2_X1 U838 ( .A(G2446), .B(G2451), .Z(n771) );
  XNOR2_X1 U839 ( .A(G2454), .B(KEYINPUT111), .ZN(n770) );
  XNOR2_X1 U840 ( .A(n771), .B(n770), .ZN(n778) );
  XOR2_X1 U841 ( .A(G2438), .B(G2430), .Z(n773) );
  XNOR2_X1 U842 ( .A(G2435), .B(G2443), .ZN(n772) );
  XNOR2_X1 U843 ( .A(n773), .B(n772), .ZN(n774) );
  XOR2_X1 U844 ( .A(n774), .B(G2427), .Z(n776) );
  XNOR2_X1 U845 ( .A(G1341), .B(G1348), .ZN(n775) );
  XNOR2_X1 U846 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U847 ( .A(n778), .B(n777), .ZN(n779) );
  AND2_X1 U848 ( .A1(n779), .A2(G14), .ZN(G401) );
  AND2_X1 U849 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U850 ( .A(G132), .ZN(G219) );
  INV_X1 U851 ( .A(G82), .ZN(G220) );
  INV_X1 U852 ( .A(G57), .ZN(G237) );
  NAND2_X1 U853 ( .A1(G7), .A2(G661), .ZN(n780) );
  XNOR2_X1 U854 ( .A(n780), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U855 ( .A(G223), .B(KEYINPUT69), .ZN(n842) );
  NAND2_X1 U856 ( .A1(n842), .A2(G567), .ZN(n781) );
  XOR2_X1 U857 ( .A(KEYINPUT11), .B(n781), .Z(G234) );
  INV_X1 U858 ( .A(G860), .ZN(n786) );
  OR2_X1 U859 ( .A1(n977), .A2(n786), .ZN(G153) );
  NAND2_X1 U860 ( .A1(G868), .A2(G301), .ZN(n783) );
  OR2_X1 U861 ( .A1(n969), .A2(G868), .ZN(n782) );
  NAND2_X1 U862 ( .A1(n783), .A2(n782), .ZN(G284) );
  XOR2_X1 U863 ( .A(KEYINPUT68), .B(n984), .Z(G299) );
  NAND2_X1 U864 ( .A1(G868), .A2(G286), .ZN(n785) );
  INV_X1 U865 ( .A(G868), .ZN(n825) );
  NAND2_X1 U866 ( .A1(G299), .A2(n825), .ZN(n784) );
  NAND2_X1 U867 ( .A1(n785), .A2(n784), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n786), .A2(G559), .ZN(n787) );
  NAND2_X1 U869 ( .A1(n787), .A2(n969), .ZN(n788) );
  XNOR2_X1 U870 ( .A(n788), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U871 ( .A1(G868), .A2(n977), .ZN(n791) );
  NAND2_X1 U872 ( .A1(G868), .A2(n969), .ZN(n789) );
  NOR2_X1 U873 ( .A1(G559), .A2(n789), .ZN(n790) );
  NOR2_X1 U874 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U875 ( .A1(G123), .A2(n874), .ZN(n792) );
  XNOR2_X1 U876 ( .A(n792), .B(KEYINPUT18), .ZN(n795) );
  NAND2_X1 U877 ( .A1(n594), .A2(G99), .ZN(n793) );
  XOR2_X1 U878 ( .A(KEYINPUT77), .B(n793), .Z(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U880 ( .A1(G135), .A2(n879), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G111), .A2(n875), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n1001) );
  XNOR2_X1 U884 ( .A(G2096), .B(n1001), .ZN(n801) );
  INV_X1 U885 ( .A(G2100), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n800), .ZN(G156) );
  NAND2_X1 U887 ( .A1(G80), .A2(n802), .ZN(n805) );
  NAND2_X1 U888 ( .A1(G67), .A2(n803), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n805), .A2(n804), .ZN(n810) );
  NAND2_X1 U890 ( .A1(G93), .A2(n643), .ZN(n808) );
  NAND2_X1 U891 ( .A1(G55), .A2(n806), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n808), .A2(n807), .ZN(n809) );
  OR2_X1 U893 ( .A1(n810), .A2(n809), .ZN(n824) );
  NAND2_X1 U894 ( .A1(G559), .A2(n969), .ZN(n811) );
  XOR2_X1 U895 ( .A(n977), .B(n811), .Z(n821) );
  XOR2_X1 U896 ( .A(n821), .B(KEYINPUT78), .Z(n812) );
  NOR2_X1 U897 ( .A1(G860), .A2(n812), .ZN(n813) );
  XOR2_X1 U898 ( .A(n824), .B(n813), .Z(G145) );
  INV_X1 U899 ( .A(G303), .ZN(G166) );
  XOR2_X1 U900 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n815) );
  XNOR2_X1 U901 ( .A(G299), .B(KEYINPUT19), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n815), .B(n814), .ZN(n816) );
  XOR2_X1 U903 ( .A(n824), .B(n816), .Z(n818) );
  XNOR2_X1 U904 ( .A(G290), .B(G166), .ZN(n817) );
  XNOR2_X1 U905 ( .A(n818), .B(n817), .ZN(n819) );
  XNOR2_X1 U906 ( .A(n819), .B(G305), .ZN(n820) );
  XNOR2_X1 U907 ( .A(n820), .B(G288), .ZN(n891) );
  XNOR2_X1 U908 ( .A(n891), .B(n821), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n822), .A2(G868), .ZN(n823) );
  XNOR2_X1 U910 ( .A(n823), .B(KEYINPUT84), .ZN(n827) );
  NAND2_X1 U911 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U912 ( .A1(n827), .A2(n826), .ZN(G295) );
  NAND2_X1 U913 ( .A1(G2084), .A2(G2078), .ZN(n828) );
  XNOR2_X1 U914 ( .A(n828), .B(KEYINPUT85), .ZN(n829) );
  XNOR2_X1 U915 ( .A(n829), .B(KEYINPUT20), .ZN(n830) );
  NAND2_X1 U916 ( .A1(n830), .A2(G2090), .ZN(n831) );
  XNOR2_X1 U917 ( .A(KEYINPUT21), .B(n831), .ZN(n832) );
  NAND2_X1 U918 ( .A1(n832), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U919 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U920 ( .A1(G120), .A2(G108), .ZN(n833) );
  NOR2_X1 U921 ( .A1(G237), .A2(n833), .ZN(n834) );
  NAND2_X1 U922 ( .A1(G69), .A2(n834), .ZN(n847) );
  NAND2_X1 U923 ( .A1(n847), .A2(G567), .ZN(n840) );
  NOR2_X1 U924 ( .A1(G220), .A2(G219), .ZN(n835) );
  XOR2_X1 U925 ( .A(KEYINPUT22), .B(n835), .Z(n836) );
  NOR2_X1 U926 ( .A1(G218), .A2(n836), .ZN(n837) );
  NAND2_X1 U927 ( .A1(G96), .A2(n837), .ZN(n846) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n846), .ZN(n838) );
  XNOR2_X1 U929 ( .A(KEYINPUT86), .B(n838), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n923) );
  NAND2_X1 U931 ( .A1(G483), .A2(G661), .ZN(n841) );
  NOR2_X1 U932 ( .A1(n923), .A2(n841), .ZN(n845) );
  NAND2_X1 U933 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U936 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n845), .A2(n844), .ZN(G188) );
  XOR2_X1 U939 ( .A(G108), .B(KEYINPUT122), .Z(G238) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  NOR2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  NAND2_X1 U945 ( .A1(G124), .A2(n874), .ZN(n848) );
  XOR2_X1 U946 ( .A(KEYINPUT44), .B(n848), .Z(n849) );
  XNOR2_X1 U947 ( .A(n849), .B(KEYINPUT115), .ZN(n851) );
  NAND2_X1 U948 ( .A1(G100), .A2(n594), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U950 ( .A1(G136), .A2(n879), .ZN(n853) );
  NAND2_X1 U951 ( .A1(G112), .A2(n875), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U953 ( .A1(n855), .A2(n854), .ZN(G162) );
  XNOR2_X1 U954 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n856), .B(KEYINPUT117), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n859), .B(n1001), .Z(n862) );
  XOR2_X1 U958 ( .A(G160), .B(n860), .Z(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U960 ( .A(n863), .B(G162), .Z(n873) );
  NAND2_X1 U961 ( .A1(n879), .A2(G139), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G103), .A2(n594), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U964 ( .A1(G127), .A2(n874), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G115), .A2(n875), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U969 ( .A(KEYINPUT118), .B(n871), .Z(n1012) );
  XNOR2_X1 U970 ( .A(G164), .B(n1012), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n886) );
  NAND2_X1 U972 ( .A1(G130), .A2(n874), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G118), .A2(n875), .ZN(n876) );
  NAND2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U975 ( .A1(G106), .A2(n594), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n878), .B(KEYINPUT116), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G142), .A2(n879), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U979 ( .A(n882), .B(KEYINPUT45), .Z(n883) );
  NOR2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U981 ( .A(n886), .B(n885), .Z(n887) );
  XOR2_X1 U982 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U983 ( .A1(G37), .A2(n889), .ZN(n890) );
  XOR2_X1 U984 ( .A(KEYINPUT119), .B(n890), .Z(G395) );
  XNOR2_X1 U985 ( .A(n977), .B(n891), .ZN(n893) );
  XNOR2_X1 U986 ( .A(G171), .B(n969), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U988 ( .A(n894), .B(G286), .ZN(n895) );
  NOR2_X1 U989 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U990 ( .A(KEYINPUT41), .B(G1981), .Z(n897) );
  XNOR2_X1 U991 ( .A(G1961), .B(G1956), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U993 ( .A(n898), .B(KEYINPUT114), .Z(n900) );
  XNOR2_X1 U994 ( .A(G1996), .B(G1991), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U996 ( .A(G1976), .B(G1971), .Z(n902) );
  XNOR2_X1 U997 ( .A(G1986), .B(G1966), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1000 ( .A(KEYINPUT113), .B(G2474), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(G229) );
  XOR2_X1 U1002 ( .A(G2096), .B(KEYINPUT43), .Z(n908) );
  XNOR2_X1 U1003 ( .A(G2090), .B(G2678), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1005 ( .A(n909), .B(KEYINPUT112), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G2067), .B(G2072), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1008 ( .A(KEYINPUT42), .B(G2100), .Z(n913) );
  XNOR2_X1 U1009 ( .A(G2084), .B(G2078), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(G227) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G397), .A2(n917), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n923), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n918), .B(KEYINPUT120), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G395), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT121), .B(n922), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(n923), .ZN(G319) );
  INV_X1 U1022 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1023 ( .A(G2067), .B(G26), .Z(n924) );
  NAND2_X1 U1024 ( .A1(n924), .A2(G28), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(G1996), .B(G32), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(G33), .B(G2072), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(G1991), .B(G25), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(G27), .B(n927), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT53), .B(n934), .Z(n937) );
  XOR2_X1 U1034 ( .A(G34), .B(KEYINPUT54), .Z(n935) );
  XNOR2_X1 U1035 ( .A(G2084), .B(n935), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G35), .B(G2090), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1039 ( .A(KEYINPUT55), .B(n940), .Z(n941) );
  NOR2_X1 U1040 ( .A1(G29), .A2(n941), .ZN(n999) );
  XNOR2_X1 U1041 ( .A(n942), .B(G20), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(G1981), .B(G6), .ZN(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1046 ( .A(KEYINPUT59), .B(G1348), .Z(n947) );
  XNOR2_X1 U1047 ( .A(G4), .B(n947), .ZN(n948) );
  NOR2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n950), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(n951), .B(G5), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(G23), .B(G1976), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n959) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n960), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1061 ( .A(KEYINPUT61), .B(n963), .Z(n964) );
  NOR2_X1 U1062 ( .A1(G16), .A2(n964), .ZN(n996) );
  XOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .Z(n993) );
  INV_X1 U1064 ( .A(n965), .ZN(n966) );
  NAND2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1066 ( .A(KEYINPUT124), .B(n968), .Z(n971) );
  XNOR2_X1 U1067 ( .A(n969), .B(G1348), .ZN(n970) );
  NAND2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n983) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(KEYINPUT57), .B(n974), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G171), .B(G1961), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n975) );
  NAND2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n977), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n984), .B(G1956), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n985), .B(KEYINPUT123), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1085 ( .A(KEYINPUT125), .B(n994), .Z(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(G11), .A2(n997), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(n1000), .B(KEYINPUT126), .ZN(n1027) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1011) );
  XNOR2_X1 U1091 ( .A(G160), .B(G2084), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G2090), .B(G162), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(KEYINPUT51), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XOR2_X1 U1098 ( .A(G164), .B(G2078), .Z(n1014) );
  XNOR2_X1 U1099 ( .A(G2072), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(KEYINPUT50), .B(n1015), .Z(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(KEYINPUT52), .B(n1022), .ZN(n1024) );
  INV_X1 U1106 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(G29), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

