//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT74), .B(KEYINPUT23), .Z(new_n196));
  OAI211_X1 g010(.A(new_n190), .B(new_n195), .C1(new_n196), .C2(new_n188), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n197), .B2(G110), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .A4(KEYINPUT16), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT16), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT75), .B1(new_n201), .B2(KEYINPUT16), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n199), .B(new_n205), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n206), .B(KEYINPUT75), .C1(KEYINPUT16), .C2(new_n201), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n199), .B1(new_n211), .B2(new_n205), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n198), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n191), .A2(new_n192), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n197), .B2(G110), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n201), .A2(new_n203), .A3(new_n199), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n221), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n213), .A2(new_n219), .A3(new_n224), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n230), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G217), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(G234), .B2(new_n227), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n226), .A2(new_n228), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n237), .A2(G902), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n243));
  INV_X1    g057(.A(G237), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n222), .A3(G210), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT27), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G101), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n248), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT67), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT67), .B1(new_n249), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(G116), .B(G119), .Z(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n254), .A2(KEYINPUT66), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT2), .B(G113), .Z(new_n258));
  XNOR2_X1  g072(.A(G116), .B(G119), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI22_X1  g074(.A1(new_n256), .A2(new_n260), .B1(new_n259), .B2(new_n258), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  XNOR2_X1  g076(.A(G143), .B(G146), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT0), .B(G128), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n199), .A2(G143), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G146), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n273), .A3(KEYINPUT64), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n265), .A2(new_n267), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT11), .A3(G134), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G137), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n281));
  INV_X1    g095(.A(G131), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n278), .B2(G137), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n280), .A2(new_n281), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n277), .A3(new_n282), .A4(new_n279), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT65), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n277), .A3(new_n279), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G131), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n275), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT1), .B1(new_n269), .B2(G146), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n271), .A2(G128), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n268), .B(new_n270), .C1(KEYINPUT1), .C2(new_n187), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n278), .A2(G137), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n276), .A2(G134), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n285), .B2(new_n287), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n261), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT68), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n288), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT66), .B1(new_n254), .B2(new_n255), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n258), .A2(new_n257), .A3(new_n259), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n304), .A2(new_n305), .B1(new_n254), .B2(new_n255), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n285), .A2(new_n287), .B1(G131), .B2(new_n289), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n303), .B(new_n306), .C1(new_n307), .C2(new_n275), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n300), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n286), .A2(KEYINPUT65), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n286), .A2(KEYINPUT65), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n290), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n275), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n303), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT68), .A3(new_n261), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n309), .A2(KEYINPUT28), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n308), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n253), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT30), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n314), .B2(new_n303), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n291), .A2(new_n299), .A3(KEYINPUT30), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n261), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n249), .A2(new_n250), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n308), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n314), .A2(new_n321), .A3(new_n303), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT30), .B1(new_n291), .B2(new_n299), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n306), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n308), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT31), .A3(new_n326), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n320), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n243), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n253), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n309), .A2(KEYINPUT28), .A3(new_n316), .ZN(new_n341));
  INV_X1    g155(.A(new_n319), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT31), .B1(new_n334), .B2(new_n326), .ZN(new_n344));
  NOR4_X1   g158(.A1(new_n332), .A2(new_n333), .A3(new_n328), .A4(new_n325), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT69), .A3(new_n337), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT32), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n339), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n338), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n319), .A2(new_n253), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n306), .B1(new_n314), .B2(new_n303), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n318), .B1(new_n356), .B2(KEYINPUT68), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n309), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT70), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n353), .B(new_n354), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n341), .A2(KEYINPUT70), .A3(new_n355), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT71), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n354), .A2(new_n353), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT70), .B1(new_n341), .B2(new_n355), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n358), .A2(new_n359), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n363), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n319), .B(KEYINPUT73), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT72), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n300), .A2(new_n369), .A3(new_n308), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n261), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n370), .A2(KEYINPUT28), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n325), .A2(new_n353), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n362), .A2(new_n367), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G472), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n242), .B1(new_n352), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT88), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n218), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n218), .A2(new_n380), .A3(new_n379), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n201), .A2(new_n203), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n382), .B(new_n383), .C1(new_n199), .C2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n199), .ZN(new_n386));
  INV_X1    g200(.A(new_n383), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(new_n381), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n244), .A2(new_n222), .A3(G214), .ZN(new_n390));
  OR3_X1    g204(.A1(new_n390), .A2(KEYINPUT86), .A3(new_n269), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT86), .B1(new_n390), .B2(new_n269), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n244), .A2(new_n222), .A3(KEYINPUT84), .A4(G214), .ZN(new_n396));
  AND4_X1   g210(.A1(KEYINPUT85), .A2(new_n395), .A3(new_n269), .A4(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(G143), .B1(new_n390), .B2(new_n394), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT85), .B1(new_n398), .B2(new_n396), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n393), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT18), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(new_n282), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI221_X1 g217(.A(new_n393), .B1(new_n401), .B2(new_n282), .C1(new_n397), .C2(new_n399), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n389), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(G131), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n282), .B(new_n393), .C1(new_n397), .C2(new_n399), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT17), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n209), .B(new_n217), .C1(new_n406), .C2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n405), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G113), .B(G122), .ZN(new_n413));
  INV_X1    g227(.A(G104), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n405), .B(new_n415), .C1(new_n409), .C2(new_n411), .ZN(new_n418));
  AOI21_X1  g232(.A(G902), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G475), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n405), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n384), .A2(KEYINPUT90), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT19), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n217), .B1(new_n425), .B2(G146), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n408), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n406), .A2(KEYINPUT89), .A3(new_n407), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT91), .B1(new_n430), .B2(new_n415), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT91), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n406), .A2(KEYINPUT89), .A3(new_n407), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT89), .B1(new_n406), .B2(new_n407), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n433), .A2(new_n434), .A3(new_n426), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n432), .B(new_n416), .C1(new_n435), .C2(new_n423), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n431), .A2(new_n436), .A3(new_n418), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n438));
  NOR2_X1   g252(.A1(G475), .A2(G902), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n438), .B1(new_n437), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n422), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G952), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G953), .ZN(new_n444));
  INV_X1    g258(.A(G234), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(new_n244), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT94), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(G902), .B(G953), .C1(new_n445), .C2(new_n244), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT95), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(G898), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT9), .B(G234), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n454), .A2(new_n236), .A3(G953), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT92), .B1(new_n187), .B2(G143), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n269), .A3(G128), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT13), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT93), .ZN(new_n463));
  INV_X1    g277(.A(new_n460), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n464), .A2(KEYINPUT13), .B1(new_n187), .B2(G143), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n278), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n460), .B1(G128), .B2(new_n269), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n467), .A2(G134), .ZN(new_n468));
  XOR2_X1   g282(.A(G116), .B(G122), .Z(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(G107), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n467), .B(new_n278), .ZN(new_n473));
  INV_X1    g287(.A(G107), .ZN(new_n474));
  INV_X1    g288(.A(G122), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G116), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n476), .B2(KEYINPUT14), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n469), .B(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n456), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  OAI221_X1 g294(.A(new_n455), .B1(new_n473), .B2(new_n478), .C1(new_n466), .C2(new_n471), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n227), .ZN(new_n483));
  INV_X1    g297(.A(G478), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n483), .B(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n442), .A2(new_n453), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G214), .B1(G237), .B2(G902), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n488), .B(KEYINPUT81), .Z(new_n489));
  OAI21_X1  g303(.A(G210), .B1(G237), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n293), .A2(new_n294), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n202), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n313), .B2(new_n202), .ZN(new_n494));
  INV_X1    g308(.A(G224), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(G953), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n494), .B(new_n496), .Z(new_n497));
  OR2_X1    g311(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n474), .A2(G104), .ZN(new_n499));
  AND2_X1   g313(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G101), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n414), .A2(G107), .ZN(new_n503));
  NOR2_X1   g317(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(G104), .A3(new_n474), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n499), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G101), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n304), .A2(new_n305), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT5), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n189), .A3(G116), .ZN(new_n512));
  OAI211_X1 g326(.A(G113), .B(new_n512), .C1(new_n254), .C2(new_n511), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n505), .A2(new_n503), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n414), .A2(G107), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n504), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n515), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT4), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n501), .A2(KEYINPUT78), .A3(new_n503), .A4(new_n505), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(G101), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n261), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n502), .B1(new_n526), .B2(new_n515), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n525), .B1(new_n527), .B2(new_n522), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n514), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT82), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT82), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(new_n514), .C1(new_n524), .C2(new_n528), .ZN(new_n532));
  XNOR2_X1  g346(.A(G110), .B(G122), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n514), .B(new_n533), .C1(new_n524), .C2(new_n528), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT6), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n533), .B1(new_n529), .B2(KEYINPUT82), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(KEYINPUT6), .A3(new_n532), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n497), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT7), .B1(new_n495), .B2(G953), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n494), .B(new_n542), .Z(new_n543));
  AND2_X1   g357(.A1(new_n510), .A2(new_n513), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n544), .A2(new_n509), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n514), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n533), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n536), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n227), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n491), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n497), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n539), .A2(KEYINPUT6), .A3(new_n532), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n539), .A2(new_n532), .B1(KEYINPUT6), .B2(new_n536), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n494), .B(new_n542), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n546), .B2(new_n547), .ZN(new_n558));
  AOI21_X1  g372(.A(G902), .B1(new_n558), .B2(new_n536), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n490), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n489), .B1(new_n552), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n520), .A2(G101), .A3(new_n522), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n313), .B(new_n523), .C1(new_n564), .C2(new_n525), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n506), .A2(new_n294), .A3(new_n293), .A4(new_n508), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n509), .A2(KEYINPUT10), .A3(new_n294), .A4(new_n293), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n565), .A2(new_n307), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n571));
  INV_X1    g385(.A(new_n566), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n506), .A2(new_n508), .B1(new_n294), .B2(new_n293), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n312), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n573), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n307), .B1(new_n575), .B2(new_n566), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n577));
  OAI21_X1  g391(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G140), .ZN(new_n579));
  INV_X1    g393(.A(G227), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G953), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n579), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n570), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n523), .A2(new_n313), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n568), .B(new_n569), .C1(new_n585), .C2(new_n528), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n312), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(new_n570), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n588), .B2(new_n583), .ZN(new_n589));
  INV_X1    g403(.A(G469), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n227), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n227), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n570), .A2(new_n578), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n582), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT80), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n583), .C1(new_n586), .C2(new_n312), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n587), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n570), .B2(new_n583), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n591), .B(new_n593), .C1(new_n590), .C2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G221), .B1(new_n454), .B2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n562), .A2(new_n563), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n378), .A2(new_n487), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  INV_X1    g420(.A(new_n453), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n561), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n484), .A2(new_n227), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n483), .B2(G478), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n456), .B2(KEYINPUT96), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n482), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n480), .A2(new_n481), .A3(new_n613), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n484), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n608), .A2(new_n442), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(G472), .B1(new_n336), .B2(G902), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n339), .A2(new_n620), .A3(new_n347), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n621), .A2(new_n603), .A3(new_n242), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  NAND3_X1  g439(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n626), .A2(KEYINPUT97), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n437), .A2(new_n439), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT20), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(KEYINPUT97), .A3(new_n626), .ZN(new_n630));
  OR3_X1    g444(.A1(new_n419), .A2(KEYINPUT98), .A3(new_n420), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT98), .B1(new_n419), .B2(new_n420), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n631), .A2(new_n486), .A3(new_n632), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n608), .A2(new_n627), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n622), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT99), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT35), .B(G107), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  INV_X1    g452(.A(new_n621), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n220), .B(KEYINPUT100), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n643), .A2(new_n240), .B1(new_n237), .B2(new_n235), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n604), .A2(new_n487), .A3(new_n639), .A4(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n448), .B1(new_n649), .B2(new_n451), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n633), .A2(new_n630), .A3(new_n627), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n377), .A2(new_n351), .A3(new_n349), .ZN(new_n654));
  INV_X1    g468(.A(new_n561), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n603), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n653), .A2(new_n654), .A3(new_n645), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  NAND2_X1  g472(.A1(new_n442), .A2(new_n486), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n489), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n661), .A3(new_n644), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n327), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n370), .A2(new_n340), .A3(new_n371), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n227), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n352), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n352), .A2(KEYINPUT101), .A3(new_n668), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n662), .A2(new_n663), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n552), .A2(new_n560), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT38), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n650), .B(KEYINPUT39), .Z(new_n678));
  NAND3_X1  g492(.A1(new_n601), .A2(new_n602), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n664), .A2(new_n673), .A3(new_n674), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  NAND3_X1  g499(.A1(new_n442), .A2(new_n618), .A3(new_n651), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n654), .A3(new_n645), .A4(new_n656), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NAND2_X1  g503(.A1(new_n589), .A2(new_n227), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(new_n602), .A3(new_n591), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n378), .A2(new_n619), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT41), .B(G113), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  NAND3_X1  g509(.A1(new_n634), .A2(new_n378), .A3(new_n692), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT103), .B(G116), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G18));
  NAND2_X1  g512(.A1(new_n692), .A2(new_n561), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n487), .A2(new_n654), .A3(new_n700), .A4(new_n645), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  NOR2_X1   g516(.A1(new_n659), .A2(new_n655), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n373), .A2(new_n253), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n344), .A2(new_n345), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n337), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n620), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n242), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n703), .A2(new_n607), .A3(new_n692), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  NAND3_X1  g524(.A1(new_n645), .A2(new_n620), .A3(new_n706), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n686), .A2(new_n699), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n202), .ZN(G27));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  INV_X1    g528(.A(new_n242), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n552), .A2(new_n560), .A3(new_n661), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n603), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n654), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n714), .B1(new_n718), .B2(new_n686), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n350), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT104), .B1(new_n336), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n348), .B1(new_n336), .B2(new_n338), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n346), .A2(new_n724), .A3(new_n350), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n722), .A2(new_n723), .A3(new_n725), .A4(KEYINPUT105), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n377), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n715), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT106), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n733), .A3(new_n715), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n687), .A2(KEYINPUT42), .A3(new_n717), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n720), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n282), .ZN(G33));
  NOR2_X1   g553(.A1(new_n718), .A2(new_n652), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT107), .B(G134), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G36));
  NOR2_X1   g556(.A1(new_n639), .A2(new_n644), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n421), .B1(new_n629), .B2(new_n626), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n744), .B2(new_n618), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n422), .B(new_n618), .C1(new_n440), .C2(new_n441), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n743), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n743), .B(KEYINPUT44), .C1(new_n745), .C2(new_n748), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n590), .B1(new_n600), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT45), .B(new_n595), .C1(new_n598), .C2(new_n599), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n592), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n591), .B1(new_n756), .B2(KEYINPUT46), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  AOI211_X1 g572(.A(new_n758), .B(new_n592), .C1(new_n754), .C2(new_n755), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n602), .B(new_n678), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n716), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n751), .A2(new_n752), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  OAI21_X1  g579(.A(new_n602), .B1(new_n757), .B2(new_n759), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT47), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n242), .A2(new_n552), .A3(new_n560), .A4(new_n661), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n377), .A2(new_n768), .A3(new_n351), .A4(new_n349), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n686), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n771), .B(new_n602), .C1(new_n757), .C2(new_n759), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n767), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  NAND3_X1  g588(.A1(new_n715), .A2(new_n602), .A3(new_n661), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n691), .A2(new_n591), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n775), .B(new_n746), .C1(KEYINPUT49), .C2(new_n776), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT109), .Z(new_n778));
  INV_X1    g592(.A(new_n673), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n776), .A2(KEYINPUT49), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n677), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n746), .B(new_n747), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n448), .ZN(new_n783));
  INV_X1    g597(.A(new_n711), .ZN(new_n784));
  INV_X1    g598(.A(new_n716), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n692), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n692), .A3(KEYINPUT116), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n783), .A2(KEYINPUT117), .A3(new_n784), .A4(new_n790), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n242), .B(new_n447), .C1(new_n788), .C2(new_n789), .ZN(new_n792));
  INV_X1    g606(.A(new_n618), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n744), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n792), .A2(new_n671), .A3(new_n672), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n691), .A2(new_n602), .A3(new_n591), .A4(new_n489), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT115), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(KEYINPUT115), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n677), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n448), .A3(new_n708), .A4(new_n782), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n762), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n782), .A2(new_n448), .A3(new_n806), .A4(new_n708), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n767), .A2(new_n772), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n602), .B2(new_n776), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n783), .A2(new_n784), .A3(new_n790), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n797), .A2(new_n805), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n816), .B2(new_n817), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n735), .A2(new_n783), .A3(new_n790), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n779), .A2(new_n442), .A3(new_n618), .A4(new_n792), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n783), .A2(new_n700), .A3(new_n708), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n444), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n819), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n645), .A2(new_n650), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n669), .A2(new_n656), .A3(new_n660), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n712), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n657), .A2(new_n828), .A3(new_n829), .A4(new_n688), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n654), .A2(new_n656), .A3(new_n645), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n712), .B1(new_n834), .B2(new_n653), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n688), .A4(new_n828), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n832), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n830), .A2(KEYINPUT112), .A3(new_n831), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n696), .A2(new_n605), .A3(new_n693), .A4(new_n709), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n442), .A2(new_n793), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n442), .B2(new_n486), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n562), .A2(new_n563), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n607), .A3(new_n622), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n646), .B(new_n701), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n734), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n733), .B1(new_n730), .B2(new_n715), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n719), .B1(new_n850), .B2(new_n736), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n687), .A2(new_n784), .A3(new_n717), .ZN(new_n852));
  INV_X1    g666(.A(new_n486), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n631), .A3(new_n632), .A4(new_n651), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n603), .A3(new_n716), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n630), .A2(new_n627), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n654), .A4(new_n645), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT110), .B1(new_n858), .B2(new_n740), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n378), .A2(new_n653), .A3(new_n717), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT110), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n852), .A3(new_n861), .A4(new_n857), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AND4_X1   g677(.A1(KEYINPUT53), .A2(new_n847), .A3(new_n851), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n832), .A2(new_n836), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n851), .A3(new_n863), .A4(new_n847), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n840), .A2(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n866), .A2(new_n867), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n847), .A2(new_n851), .A3(new_n863), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT111), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n847), .A2(new_n851), .A3(new_n863), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n840), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n871), .B1(new_n876), .B2(new_n867), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n826), .B(new_n870), .C1(new_n869), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n781), .B1(new_n879), .B2(new_n880), .ZN(G75));
  OAI21_X1  g695(.A(KEYINPUT118), .B1(new_n868), .B2(new_n227), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n866), .A2(new_n867), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n838), .A2(new_n839), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n847), .A2(new_n851), .A3(new_n863), .A4(KEYINPUT53), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n883), .B(G902), .C1(new_n884), .C2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n882), .A2(new_n491), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n554), .A2(new_n555), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n497), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n556), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT55), .ZN(new_n893));
  XOR2_X1   g707(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n443), .A2(G953), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT120), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(G210), .B(G902), .C1(new_n884), .C2(new_n887), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n902), .B2(new_n893), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n896), .A2(new_n903), .ZN(G51));
  XNOR2_X1  g718(.A(new_n592), .B(KEYINPUT57), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n884), .A2(new_n887), .A3(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n840), .A2(new_n864), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n866), .A2(new_n867), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n869), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n905), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n589), .B(KEYINPUT121), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n754), .A2(new_n755), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT122), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n882), .A2(new_n888), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n899), .B1(new_n912), .B2(new_n915), .ZN(G54));
  AND3_X1   g730(.A1(new_n437), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n882), .A2(new_n888), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n898), .ZN(new_n919));
  INV_X1    g733(.A(new_n437), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n882), .A2(new_n888), .A3(KEYINPUT58), .A4(G475), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G60));
  NAND2_X1  g736(.A1(new_n615), .A2(new_n616), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n609), .B(KEYINPUT59), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n906), .B2(new_n909), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n898), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n870), .B1(new_n877), .B2(new_n869), .ZN(new_n928));
  INV_X1    g742(.A(new_n924), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n923), .B2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n884), .B2(new_n887), .ZN(new_n935));
  INV_X1    g749(.A(new_n239), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n899), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n868), .A2(new_n933), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n643), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(KEYINPUT61), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n452), .B2(new_n495), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n847), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n890), .B1(G898), .B2(new_n222), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  INV_X1    g762(.A(new_n684), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n657), .A2(new_n829), .A3(new_n688), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT62), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n657), .A2(new_n688), .A3(new_n829), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n684), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n752), .A2(new_n763), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT44), .B1(new_n782), .B2(new_n743), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n773), .ZN(new_n958));
  INV_X1    g772(.A(new_n678), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n718), .A2(new_n843), .A3(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n951), .A2(new_n954), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n222), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n330), .A2(new_n331), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n425), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT123), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n649), .A2(new_n222), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n773), .A2(new_n860), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n760), .A2(new_n655), .A3(new_n659), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n848), .B2(new_n849), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n736), .B1(new_n732), .B2(new_n734), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n969), .B(new_n971), .C1(new_n972), .C2(new_n720), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n957), .B2(new_n950), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n952), .A2(new_n764), .A3(KEYINPUT124), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n965), .B(new_n968), .C1(new_n977), .C2(new_n222), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n967), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(G953), .B1(new_n580), .B2(new_n649), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G72));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n334), .B(KEYINPUT125), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n984), .A2(new_n326), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n975), .A2(new_n976), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n969), .A2(new_n971), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(new_n738), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n847), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  AOI21_X1  g805(.A(new_n985), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n983), .B1(new_n992), .B2(new_n899), .ZN(new_n993));
  INV_X1    g807(.A(new_n991), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n977), .B2(new_n847), .ZN(new_n995));
  OAI211_X1 g809(.A(KEYINPUT126), .B(new_n898), .C1(new_n995), .C2(new_n985), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n951), .A2(new_n847), .A3(new_n954), .A4(new_n961), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n991), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n326), .A3(new_n984), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n994), .B1(new_n327), .B2(new_n354), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n877), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n982), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n877), .A2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n993), .A2(new_n996), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1005), .A2(new_n1006), .A3(KEYINPUT127), .A4(new_n1000), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1004), .A2(new_n1007), .ZN(G57));
endmodule


