

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579;

  XNOR2_X1 U321 ( .A(n338), .B(n290), .ZN(n339) );
  XNOR2_X1 U322 ( .A(n356), .B(KEYINPUT96), .ZN(n495) );
  XNOR2_X1 U323 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U324 ( .A(n545), .B(KEYINPUT28), .Z(n511) );
  NOR2_X1 U325 ( .A1(n577), .A2(n409), .ZN(n289) );
  XOR2_X1 U326 ( .A(G29GAT), .B(KEYINPUT1), .Z(n290) );
  INV_X1 U327 ( .A(n534), .ZN(n409) );
  XOR2_X1 U328 ( .A(G1GAT), .B(G127GAT), .Z(n331) );
  AND2_X1 U329 ( .A1(n455), .A2(n289), .ZN(n411) );
  XOR2_X1 U330 ( .A(KEYINPUT38), .B(n449), .Z(n472) );
  XNOR2_X1 U331 ( .A(n450), .B(KEYINPUT40), .ZN(n451) );
  XNOR2_X1 U332 ( .A(n452), .B(n451), .ZN(G1330GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n292) );
  XNOR2_X1 U334 ( .A(G15GAT), .B(KEYINPUT86), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n309) );
  XOR2_X1 U336 ( .A(G71GAT), .B(G120GAT), .Z(n294) );
  XNOR2_X1 U337 ( .A(G183GAT), .B(G127GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U339 ( .A(n295), .B(KEYINPUT64), .Z(n297) );
  XOR2_X1 U340 ( .A(G113GAT), .B(KEYINPUT0), .Z(n335) );
  XNOR2_X1 U341 ( .A(n335), .B(G99GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U343 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n299) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U346 ( .A(n301), .B(n300), .Z(n307) );
  XNOR2_X1 U347 ( .A(G176GAT), .B(KEYINPUT18), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n302), .B(KEYINPUT17), .ZN(n303) );
  XOR2_X1 U349 ( .A(n303), .B(KEYINPUT19), .Z(n305) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G190GAT), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n354) );
  XOR2_X1 U352 ( .A(G43GAT), .B(G134GAT), .Z(n391) );
  XNOR2_X1 U353 ( .A(n354), .B(n391), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U355 ( .A(n309), .B(n308), .Z(n548) );
  XOR2_X1 U356 ( .A(n548), .B(KEYINPUT88), .Z(n359) );
  XOR2_X1 U357 ( .A(G50GAT), .B(G218GAT), .Z(n381) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n310), .B(KEYINPUT90), .ZN(n350) );
  XNOR2_X1 U360 ( .A(n381), .B(n350), .ZN(n311) );
  XOR2_X1 U361 ( .A(G106GAT), .B(G78GAT), .Z(n442) );
  XNOR2_X1 U362 ( .A(n311), .B(n442), .ZN(n317) );
  XOR2_X1 U363 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n313) );
  XNOR2_X1 U364 ( .A(G141GAT), .B(G162GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n332) );
  XOR2_X1 U366 ( .A(n332), .B(G148GAT), .Z(n315) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U369 ( .A(n317), .B(n316), .Z(n325) );
  XOR2_X1 U370 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n319) );
  XNOR2_X1 U371 ( .A(G204GAT), .B(G155GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U373 ( .A(KEYINPUT22), .B(G211GAT), .Z(n321) );
  XNOR2_X1 U374 ( .A(G22GAT), .B(KEYINPUT89), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n545) );
  XOR2_X1 U378 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n327) );
  XNOR2_X1 U379 ( .A(KEYINPUT5), .B(KEYINPUT92), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n342) );
  XOR2_X1 U381 ( .A(KEYINPUT4), .B(G57GAT), .Z(n329) );
  NAND2_X1 U382 ( .A1(G225GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U384 ( .A(n330), .B(KEYINPUT93), .Z(n334) );
  XOR2_X1 U385 ( .A(G155GAT), .B(n331), .Z(n396) );
  XNOR2_X1 U386 ( .A(n332), .B(n396), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n340) );
  XOR2_X1 U388 ( .A(G120GAT), .B(G148GAT), .Z(n431) );
  XOR2_X1 U389 ( .A(G85GAT), .B(n431), .Z(n337) );
  XNOR2_X1 U390 ( .A(G134GAT), .B(n335), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U392 ( .A(n342), .B(n341), .Z(n371) );
  XNOR2_X1 U393 ( .A(KEYINPUT94), .B(n371), .ZN(n543) );
  XOR2_X1 U394 ( .A(G218GAT), .B(G36GAT), .Z(n344) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n347) );
  XOR2_X1 U397 ( .A(KEYINPUT81), .B(G211GAT), .Z(n346) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G183GAT), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n404) );
  XOR2_X1 U400 ( .A(n347), .B(n404), .Z(n352) );
  XOR2_X1 U401 ( .A(G64GAT), .B(KEYINPUT77), .Z(n349) );
  XNOR2_X1 U402 ( .A(G204GAT), .B(G92GAT), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n445) );
  XNOR2_X1 U404 ( .A(n350), .B(n445), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n540) );
  XOR2_X1 U407 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n355) );
  XNOR2_X1 U408 ( .A(n540), .B(n355), .ZN(n366) );
  NOR2_X1 U409 ( .A1(n543), .A2(n366), .ZN(n356) );
  NAND2_X1 U410 ( .A1(n511), .A2(n495), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n357), .B(KEYINPUT97), .ZN(n358) );
  NAND2_X1 U412 ( .A1(n359), .A2(n358), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n360), .B(KEYINPUT98), .ZN(n373) );
  INV_X1 U414 ( .A(n548), .ZN(n490) );
  NOR2_X1 U415 ( .A1(n490), .A2(n540), .ZN(n361) );
  NOR2_X1 U416 ( .A1(n545), .A2(n361), .ZN(n362) );
  XNOR2_X1 U417 ( .A(KEYINPUT25), .B(n362), .ZN(n369) );
  XOR2_X1 U418 ( .A(KEYINPUT100), .B(KEYINPUT26), .Z(n364) );
  NAND2_X1 U419 ( .A1(n545), .A2(n490), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U421 ( .A(KEYINPUT99), .B(n365), .ZN(n564) );
  NOR2_X1 U422 ( .A1(n366), .A2(n564), .ZN(n367) );
  XNOR2_X1 U423 ( .A(KEYINPUT101), .B(n367), .ZN(n368) );
  NAND2_X1 U424 ( .A1(n369), .A2(n368), .ZN(n370) );
  NAND2_X1 U425 ( .A1(n371), .A2(n370), .ZN(n372) );
  NAND2_X1 U426 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U427 ( .A(KEYINPUT102), .B(n374), .ZN(n455) );
  XOR2_X1 U428 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n376) );
  XNOR2_X1 U429 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U431 ( .A(G99GAT), .B(G85GAT), .Z(n432) );
  XOR2_X1 U432 ( .A(n377), .B(n432), .Z(n383) );
  XOR2_X1 U433 ( .A(KEYINPUT8), .B(KEYINPUT71), .Z(n379) );
  XNOR2_X1 U434 ( .A(G36GAT), .B(G29GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U436 ( .A(KEYINPUT7), .B(n380), .Z(n428) );
  XNOR2_X1 U437 ( .A(n428), .B(n381), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U439 ( .A(G92GAT), .B(G106GAT), .Z(n385) );
  NAND2_X1 U440 ( .A1(G232GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U442 ( .A(n387), .B(n386), .Z(n393) );
  XOR2_X1 U443 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n389) );
  XNOR2_X1 U444 ( .A(G190GAT), .B(G162GAT), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n501) );
  XNOR2_X1 U448 ( .A(KEYINPUT36), .B(n501), .ZN(n577) );
  XOR2_X1 U449 ( .A(KEYINPUT13), .B(KEYINPUT73), .Z(n395) );
  XNOR2_X1 U450 ( .A(G71GAT), .B(G57GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n446) );
  XOR2_X1 U452 ( .A(n446), .B(n396), .Z(n408) );
  XOR2_X1 U453 ( .A(KEYINPUT82), .B(KEYINPUT15), .Z(n398) );
  XNOR2_X1 U454 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U456 ( .A(G64GAT), .B(G78GAT), .Z(n400) );
  NAND2_X1 U457 ( .A1(G231GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U459 ( .A(n402), .B(n401), .Z(n406) );
  XNOR2_X1 U460 ( .A(G15GAT), .B(G22GAT), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n403), .B(KEYINPUT72), .ZN(n423) );
  XNOR2_X1 U462 ( .A(n423), .B(n404), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n534) );
  INV_X1 U465 ( .A(KEYINPUT37), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n487) );
  XOR2_X1 U467 ( .A(KEYINPUT68), .B(G1GAT), .Z(n413) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(G197GAT), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U470 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U473 ( .A(n417), .B(n416), .Z(n422) );
  XOR2_X1 U474 ( .A(KEYINPUT29), .B(G8GAT), .Z(n419) );
  NAND2_X1 U475 ( .A1(G229GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U477 ( .A(KEYINPUT66), .B(n420), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U479 ( .A(G50GAT), .B(G43GAT), .Z(n425) );
  XNOR2_X1 U480 ( .A(G113GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U482 ( .A(n427), .B(n426), .Z(n430) );
  XNOR2_X1 U483 ( .A(G169GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n566) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U486 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U488 ( .A(KEYINPUT76), .B(KEYINPUT74), .Z(n436) );
  XNOR2_X1 U489 ( .A(KEYINPUT31), .B(KEYINPUT78), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U491 ( .A(n438), .B(n437), .Z(n444) );
  XOR2_X1 U492 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n440) );
  XNOR2_X1 U493 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U497 ( .A(n446), .B(n445), .Z(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n571) );
  AND2_X1 U499 ( .A1(n566), .A2(n571), .ZN(n458) );
  AND2_X1 U500 ( .A1(n487), .A2(n458), .ZN(n449) );
  NOR2_X1 U501 ( .A1(n472), .A2(n490), .ZN(n452) );
  INV_X1 U502 ( .A(G43GAT), .ZN(n450) );
  INV_X1 U503 ( .A(n501), .ZN(n561) );
  NOR2_X1 U504 ( .A1(n561), .A2(n534), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT83), .B(n453), .Z(n454) );
  XNOR2_X1 U506 ( .A(KEYINPUT16), .B(n454), .ZN(n456) );
  NAND2_X1 U507 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n457), .B(KEYINPUT103), .ZN(n474) );
  NAND2_X1 U509 ( .A1(n458), .A2(n474), .ZN(n465) );
  NOR2_X1 U510 ( .A1(n543), .A2(n465), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U513 ( .A(G1GAT), .B(n461), .Z(G1324GAT) );
  NOR2_X1 U514 ( .A1(n540), .A2(n465), .ZN(n462) );
  XOR2_X1 U515 ( .A(G8GAT), .B(n462), .Z(G1325GAT) );
  NOR2_X1 U516 ( .A1(n490), .A2(n465), .ZN(n464) );
  XNOR2_X1 U517 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n464), .B(n463), .ZN(G1326GAT) );
  NOR2_X1 U519 ( .A1(n511), .A2(n465), .ZN(n467) );
  XNOR2_X1 U520 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n467), .B(n466), .ZN(G1327GAT) );
  NOR2_X1 U522 ( .A1(n472), .A2(n543), .ZN(n469) );
  XNOR2_X1 U523 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n468) );
  XNOR2_X1 U524 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U525 ( .A(G29GAT), .B(n470), .ZN(G1328GAT) );
  NOR2_X1 U526 ( .A1(n472), .A2(n540), .ZN(n471) );
  XOR2_X1 U527 ( .A(G36GAT), .B(n471), .Z(G1329GAT) );
  NOR2_X1 U528 ( .A1(n511), .A2(n472), .ZN(n473) );
  XOR2_X1 U529 ( .A(G50GAT), .B(n473), .Z(G1331GAT) );
  XNOR2_X1 U530 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n478) );
  XOR2_X1 U531 ( .A(KEYINPUT41), .B(n571), .Z(n496) );
  NOR2_X1 U532 ( .A1(n566), .A2(n496), .ZN(n486) );
  NAND2_X1 U533 ( .A1(n474), .A2(n486), .ZN(n483) );
  NOR2_X1 U534 ( .A1(n543), .A2(n483), .ZN(n476) );
  XNOR2_X1 U535 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(G1332GAT) );
  NOR2_X1 U538 ( .A1(n540), .A2(n483), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(G1333GAT) );
  NOR2_X1 U541 ( .A1(n490), .A2(n483), .ZN(n481) );
  XOR2_X1 U542 ( .A(KEYINPUT110), .B(n481), .Z(n482) );
  XNOR2_X1 U543 ( .A(G71GAT), .B(n482), .ZN(G1334GAT) );
  NOR2_X1 U544 ( .A1(n511), .A2(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(G1335GAT) );
  NAND2_X1 U547 ( .A1(n487), .A2(n486), .ZN(n492) );
  NOR2_X1 U548 ( .A1(n543), .A2(n492), .ZN(n488) );
  XOR2_X1 U549 ( .A(G85GAT), .B(n488), .Z(G1336GAT) );
  NOR2_X1 U550 ( .A1(n540), .A2(n492), .ZN(n489) );
  XOR2_X1 U551 ( .A(G92GAT), .B(n489), .Z(G1337GAT) );
  NOR2_X1 U552 ( .A1(n490), .A2(n492), .ZN(n491) );
  XOR2_X1 U553 ( .A(G99GAT), .B(n491), .Z(G1338GAT) );
  NOR2_X1 U554 ( .A1(n511), .A2(n492), .ZN(n493) );
  XOR2_X1 U555 ( .A(KEYINPUT44), .B(n493), .Z(n494) );
  XNOR2_X1 U556 ( .A(G106GAT), .B(n494), .ZN(G1339GAT) );
  XOR2_X1 U557 ( .A(G113GAT), .B(KEYINPUT115), .Z(n515) );
  INV_X1 U558 ( .A(n495), .ZN(n509) );
  XOR2_X1 U559 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n498) );
  INV_X1 U560 ( .A(n496), .ZN(n554) );
  NAND2_X1 U561 ( .A1(n554), .A2(n566), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(KEYINPUT111), .B(n534), .ZN(n558) );
  NOR2_X1 U564 ( .A1(n499), .A2(n558), .ZN(n500) );
  NAND2_X1 U565 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(KEYINPUT47), .ZN(n507) );
  NOR2_X1 U567 ( .A1(n577), .A2(n534), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(KEYINPUT45), .ZN(n504) );
  NAND2_X1 U569 ( .A1(n504), .A2(n571), .ZN(n505) );
  NOR2_X1 U570 ( .A1(n505), .A2(n566), .ZN(n506) );
  NOR2_X1 U571 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT48), .B(n508), .ZN(n541) );
  NOR2_X1 U573 ( .A1(n509), .A2(n541), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n548), .A2(n524), .ZN(n510) );
  XNOR2_X1 U575 ( .A(KEYINPUT113), .B(n510), .ZN(n512) );
  NAND2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n513) );
  XOR2_X1 U577 ( .A(KEYINPUT114), .B(n513), .Z(n520) );
  NAND2_X1 U578 ( .A1(n566), .A2(n520), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1340GAT) );
  XOR2_X1 U580 ( .A(G120GAT), .B(KEYINPUT49), .Z(n517) );
  NAND2_X1 U581 ( .A1(n554), .A2(n520), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1341GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n558), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT50), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G127GAT), .B(n519), .ZN(G1342GAT) );
  XOR2_X1 U586 ( .A(G134GAT), .B(KEYINPUT51), .Z(n522) );
  NAND2_X1 U587 ( .A1(n520), .A2(n561), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1343GAT) );
  INV_X1 U589 ( .A(n564), .ZN(n523) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U591 ( .A(KEYINPUT116), .B(n525), .Z(n537) );
  NAND2_X1 U592 ( .A1(n537), .A2(n566), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT117), .B(KEYINPUT119), .Z(n528) );
  XNOR2_X1 U595 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U597 ( .A(n529), .B(KEYINPUT120), .Z(n531) );
  XNOR2_X1 U598 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n533) );
  NAND2_X1 U600 ( .A1(n537), .A2(n554), .ZN(n532) );
  XOR2_X1 U601 ( .A(n533), .B(n532), .Z(G1345GAT) );
  XOR2_X1 U602 ( .A(G155GAT), .B(KEYINPUT121), .Z(n536) );
  NAND2_X1 U603 ( .A1(n409), .A2(n537), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1346GAT) );
  NAND2_X1 U605 ( .A1(n537), .A2(n561), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n538), .B(KEYINPUT122), .ZN(n539) );
  XNOR2_X1 U607 ( .A(G162GAT), .B(n539), .ZN(G1347GAT) );
  NOR2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(KEYINPUT54), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n565) );
  NOR2_X1 U611 ( .A1(n545), .A2(n565), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT123), .B(KEYINPUT55), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n549) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT124), .B(n550), .Z(n560) );
  NAND2_X1 U616 ( .A1(n560), .A2(n566), .ZN(n553) );
  XOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT125), .Z(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT126), .B(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n560), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(n557), .ZN(G1349GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  XOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT127), .Z(n568) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n574), .A2(n566), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U636 ( .A(n574), .ZN(n576) );
  OR2_X1 U637 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n409), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(n578), .Z(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

