

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U549 ( .A(KEYINPUT74), .B(n588), .Z(n973) );
  INV_X1 U550 ( .A(KEYINPUT27), .ZN(n734) );
  XNOR2_X1 U551 ( .A(n734), .B(KEYINPUT101), .ZN(n735) );
  XNOR2_X1 U552 ( .A(n736), .B(n735), .ZN(n738) );
  INV_X1 U553 ( .A(KEYINPUT29), .ZN(n751) );
  NAND2_X1 U554 ( .A1(n724), .A2(n723), .ZN(n767) );
  INV_X1 U555 ( .A(KEYINPUT72), .ZN(n579) );
  XNOR2_X1 U556 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U557 ( .A(n582), .B(n581), .ZN(n583) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n724) );
  NOR2_X1 U559 ( .A1(G651), .A2(n639), .ZN(n650) );
  NOR2_X1 U560 ( .A1(G543), .A2(G651), .ZN(n515) );
  XNOR2_X1 U561 ( .A(n515), .B(KEYINPUT64), .ZN(n651) );
  NAND2_X1 U562 ( .A1(n651), .A2(G89), .ZN(n516) );
  XNOR2_X1 U563 ( .A(n516), .B(KEYINPUT78), .ZN(n517) );
  XNOR2_X1 U564 ( .A(n517), .B(KEYINPUT4), .ZN(n519) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n639) );
  INV_X1 U566 ( .A(G651), .ZN(n521) );
  NOR2_X2 U567 ( .A1(n639), .A2(n521), .ZN(n654) );
  NAND2_X1 U568 ( .A1(G76), .A2(n654), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U570 ( .A(n520), .B(KEYINPUT5), .ZN(n528) );
  NOR2_X1 U571 ( .A1(G543), .A2(n521), .ZN(n522) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n522), .Z(n655) );
  NAND2_X1 U573 ( .A1(n655), .A2(G63), .ZN(n523) );
  XOR2_X1 U574 ( .A(KEYINPUT79), .B(n523), .Z(n525) );
  NAND2_X1 U575 ( .A1(n650), .A2(G51), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT6), .B(n526), .Z(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U579 ( .A(n529), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U580 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U581 ( .A(G2105), .ZN(n533) );
  NOR2_X1 U582 ( .A1(G2104), .A2(n533), .ZN(n871) );
  NAND2_X1 U583 ( .A1(G126), .A2(n871), .ZN(n531) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n872) );
  NAND2_X1 U585 ( .A1(G114), .A2(n872), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U587 ( .A(KEYINPUT90), .B(n532), .ZN(n539) );
  AND2_X1 U588 ( .A1(n533), .A2(G2104), .ZN(n867) );
  NAND2_X1 U589 ( .A1(G102), .A2(n867), .ZN(n537) );
  NOR2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  XOR2_X1 U591 ( .A(n534), .B(KEYINPUT17), .Z(n535) );
  XNOR2_X1 U592 ( .A(KEYINPUT66), .B(n535), .ZN(n868) );
  NAND2_X1 U593 ( .A1(G138), .A2(n868), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U595 ( .A1(n539), .A2(n538), .ZN(G164) );
  NAND2_X1 U596 ( .A1(G101), .A2(n867), .ZN(n540) );
  XOR2_X1 U597 ( .A(KEYINPUT23), .B(n540), .Z(n543) );
  NAND2_X1 U598 ( .A1(G113), .A2(n872), .ZN(n541) );
  XOR2_X1 U599 ( .A(KEYINPUT65), .B(n541), .Z(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G125), .A2(n871), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G137), .A2(n868), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U604 ( .A1(n547), .A2(n546), .ZN(G160) );
  XOR2_X1 U605 ( .A(G2427), .B(G2435), .Z(n549) );
  XNOR2_X1 U606 ( .A(G2454), .B(G2443), .ZN(n548) );
  XNOR2_X1 U607 ( .A(n549), .B(n548), .ZN(n556) );
  XOR2_X1 U608 ( .A(G2451), .B(KEYINPUT105), .Z(n551) );
  XNOR2_X1 U609 ( .A(G2430), .B(G2438), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U611 ( .A(n552), .B(G2446), .Z(n554) );
  XNOR2_X1 U612 ( .A(G1348), .B(G1341), .ZN(n553) );
  XNOR2_X1 U613 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U614 ( .A(n556), .B(n555), .ZN(n557) );
  AND2_X1 U615 ( .A1(n557), .A2(G14), .ZN(G401) );
  NAND2_X1 U616 ( .A1(G52), .A2(n650), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G64), .A2(n655), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n564) );
  NAND2_X1 U619 ( .A1(n654), .A2(G77), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G90), .A2(n651), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U623 ( .A1(n564), .A2(n563), .ZN(G171) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U625 ( .A(G57), .ZN(G237) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  NAND2_X1 U628 ( .A1(G53), .A2(n650), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G65), .A2(n655), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n654), .A2(G78), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G91), .A2(n651), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n745) );
  INV_X1 U635 ( .A(n745), .ZN(G299) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n825) );
  NAND2_X1 U639 ( .A1(n825), .A2(G567), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(KEYINPUT11), .ZN(n573) );
  XNOR2_X1 U641 ( .A(KEYINPUT69), .B(n573), .ZN(G234) );
  XOR2_X1 U642 ( .A(G860), .B(KEYINPUT75), .Z(n602) );
  NAND2_X1 U643 ( .A1(n655), .A2(G56), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT14), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G81), .A2(n651), .ZN(n575) );
  XOR2_X1 U646 ( .A(n575), .B(KEYINPUT12), .Z(n578) );
  AND2_X1 U647 ( .A1(n654), .A2(G68), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT70), .ZN(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n580) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n585), .B(KEYINPUT73), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G43), .A2(n650), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n602), .A2(n973), .ZN(G153) );
  XOR2_X1 U656 ( .A(G171), .B(KEYINPUT76), .Z(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U658 ( .A1(G66), .A2(n655), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G79), .A2(n654), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G54), .A2(n650), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G92), .A2(n651), .ZN(n591) );
  XNOR2_X1 U663 ( .A(KEYINPUT77), .B(n591), .ZN(n592) );
  NOR2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n596), .B(KEYINPUT15), .ZN(n958) );
  INV_X1 U667 ( .A(n958), .ZN(n739) );
  INV_X1 U668 ( .A(G868), .ZN(n668) );
  NAND2_X1 U669 ( .A1(n739), .A2(n668), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(G284) );
  NOR2_X1 U671 ( .A1(G286), .A2(n668), .ZN(n600) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(G297) );
  INV_X1 U674 ( .A(G559), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n739), .A2(n603), .ZN(n604) );
  XOR2_X1 U677 ( .A(KEYINPUT16), .B(n604), .Z(G148) );
  NAND2_X1 U678 ( .A1(n958), .A2(G868), .ZN(n605) );
  NOR2_X1 U679 ( .A1(G559), .A2(n605), .ZN(n607) );
  AND2_X1 U680 ( .A1(n973), .A2(n668), .ZN(n606) );
  NOR2_X1 U681 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G123), .A2(n871), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT80), .ZN(n609) );
  XNOR2_X1 U684 ( .A(KEYINPUT18), .B(n609), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G99), .A2(n867), .ZN(n610) );
  XOR2_X1 U686 ( .A(KEYINPUT81), .B(n610), .Z(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G111), .A2(n872), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G135), .A2(n868), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n927) );
  XOR2_X1 U692 ( .A(n927), .B(G2096), .Z(n617) );
  NOR2_X1 U693 ( .A1(G2100), .A2(n617), .ZN(n618) );
  XOR2_X1 U694 ( .A(KEYINPUT82), .B(n618), .Z(G156) );
  NAND2_X1 U695 ( .A1(G559), .A2(n958), .ZN(n619) );
  XOR2_X1 U696 ( .A(n973), .B(n619), .Z(n666) );
  NOR2_X1 U697 ( .A1(G860), .A2(n666), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G55), .A2(n650), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G67), .A2(n655), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n654), .A2(G80), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G93), .A2(n651), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n669) );
  XNOR2_X1 U705 ( .A(n626), .B(n669), .ZN(G145) );
  NAND2_X1 U706 ( .A1(n655), .A2(G61), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G86), .A2(n651), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G73), .A2(n654), .ZN(n629) );
  XNOR2_X1 U710 ( .A(n629), .B(KEYINPUT83), .ZN(n630) );
  XNOR2_X1 U711 ( .A(n630), .B(KEYINPUT2), .ZN(n631) );
  NOR2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n633), .B(KEYINPUT84), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G48), .A2(n650), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G49), .A2(n650), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U719 ( .A1(n655), .A2(n638), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n639), .A2(G87), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n641), .A2(n640), .ZN(G288) );
  NAND2_X1 U722 ( .A1(n650), .A2(G47), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n654), .A2(G72), .ZN(n643) );
  NAND2_X1 U724 ( .A1(G85), .A2(n651), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U726 ( .A1(G60), .A2(n655), .ZN(n644) );
  XNOR2_X1 U727 ( .A(KEYINPUT67), .B(n644), .ZN(n645) );
  NOR2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(KEYINPUT68), .ZN(G290) );
  NAND2_X1 U731 ( .A1(n650), .A2(G50), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G88), .A2(n651), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n659) );
  NAND2_X1 U734 ( .A1(G75), .A2(n654), .ZN(n657) );
  NAND2_X1 U735 ( .A1(G62), .A2(n655), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U737 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n660), .B(KEYINPUT85), .ZN(G303) );
  INV_X1 U739 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U740 ( .A(G288), .B(KEYINPUT19), .ZN(n662) );
  XNOR2_X1 U741 ( .A(G290), .B(G166), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n669), .B(n663), .ZN(n664) );
  XNOR2_X1 U744 ( .A(n664), .B(G299), .ZN(n665) );
  XNOR2_X1 U745 ( .A(G305), .B(n665), .ZN(n898) );
  XNOR2_X1 U746 ( .A(n666), .B(n898), .ZN(n667) );
  NOR2_X1 U747 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U748 ( .A1(G868), .A2(n669), .ZN(n670) );
  NOR2_X1 U749 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U750 ( .A(KEYINPUT86), .B(n672), .Z(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U755 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U759 ( .A1(G218), .A2(n678), .ZN(n679) );
  XOR2_X1 U760 ( .A(KEYINPUT87), .B(n679), .Z(n680) );
  NAND2_X1 U761 ( .A1(G96), .A2(n680), .ZN(n830) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n830), .ZN(n685) );
  NAND2_X1 U763 ( .A1(G120), .A2(G69), .ZN(n681) );
  NOR2_X1 U764 ( .A1(G237), .A2(n681), .ZN(n682) );
  XNOR2_X1 U765 ( .A(KEYINPUT88), .B(n682), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n683), .A2(G108), .ZN(n829) );
  NAND2_X1 U767 ( .A1(G567), .A2(n829), .ZN(n684) );
  NAND2_X1 U768 ( .A1(n685), .A2(n684), .ZN(n901) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U770 ( .A1(n901), .A2(n686), .ZN(n828) );
  NAND2_X1 U771 ( .A1(G36), .A2(n828), .ZN(n687) );
  XOR2_X1 U772 ( .A(KEYINPUT89), .B(n687), .Z(G176) );
  XNOR2_X1 U773 ( .A(G1986), .B(G290), .ZN(n962) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n722) );
  NOR2_X1 U775 ( .A1(n724), .A2(n722), .ZN(n820) );
  NAND2_X1 U776 ( .A1(n962), .A2(n820), .ZN(n809) );
  XOR2_X1 U777 ( .A(n820), .B(KEYINPUT97), .Z(n707) );
  NAND2_X1 U778 ( .A1(G105), .A2(n867), .ZN(n688) );
  XOR2_X1 U779 ( .A(KEYINPUT38), .B(n688), .Z(n695) );
  NAND2_X1 U780 ( .A1(n872), .A2(G117), .ZN(n689) );
  XNOR2_X1 U781 ( .A(KEYINPUT95), .B(n689), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n871), .A2(G129), .ZN(n690) );
  XOR2_X1 U783 ( .A(KEYINPUT94), .B(n690), .Z(n691) );
  NOR2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U785 ( .A(KEYINPUT96), .B(n693), .Z(n694) );
  NOR2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U787 ( .A1(G141), .A2(n868), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n880) );
  NAND2_X1 U789 ( .A1(G1996), .A2(n880), .ZN(n706) );
  NAND2_X1 U790 ( .A1(G107), .A2(n872), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G131), .A2(n868), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U793 ( .A1(G119), .A2(n871), .ZN(n701) );
  NAND2_X1 U794 ( .A1(G95), .A2(n867), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U797 ( .A(n704), .B(KEYINPUT93), .ZN(n888) );
  NAND2_X1 U798 ( .A1(G1991), .A2(n888), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n928) );
  NAND2_X1 U800 ( .A1(n707), .A2(n928), .ZN(n708) );
  XOR2_X1 U801 ( .A(KEYINPUT98), .B(n708), .Z(n813) );
  XNOR2_X1 U802 ( .A(KEYINPUT99), .B(n813), .ZN(n720) );
  XNOR2_X1 U803 ( .A(KEYINPUT37), .B(G2067), .ZN(n818) );
  NAND2_X1 U804 ( .A1(n867), .A2(G104), .ZN(n709) );
  XOR2_X1 U805 ( .A(KEYINPUT91), .B(n709), .Z(n711) );
  NAND2_X1 U806 ( .A1(G140), .A2(n868), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n712), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n871), .A2(G128), .ZN(n713) );
  XNOR2_X1 U810 ( .A(n713), .B(KEYINPUT92), .ZN(n715) );
  NAND2_X1 U811 ( .A1(G116), .A2(n872), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U813 ( .A(KEYINPUT35), .B(n716), .Z(n717) );
  NOR2_X1 U814 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n719), .ZN(n892) );
  NOR2_X1 U816 ( .A1(n818), .A2(n892), .ZN(n940) );
  NAND2_X1 U817 ( .A1(n820), .A2(n940), .ZN(n816) );
  NAND2_X1 U818 ( .A1(n720), .A2(n816), .ZN(n721) );
  XNOR2_X1 U819 ( .A(n721), .B(KEYINPUT100), .ZN(n807) );
  INV_X1 U820 ( .A(n722), .ZN(n723) );
  NAND2_X1 U821 ( .A1(G8), .A2(n767), .ZN(n803) );
  INV_X1 U822 ( .A(n767), .ZN(n753) );
  NOR2_X1 U823 ( .A1(n753), .A2(G1348), .ZN(n726) );
  NOR2_X1 U824 ( .A1(G2067), .A2(n767), .ZN(n725) );
  NOR2_X1 U825 ( .A1(n726), .A2(n725), .ZN(n740) );
  NAND2_X1 U826 ( .A1(n739), .A2(n740), .ZN(n733) );
  NAND2_X1 U827 ( .A1(G1996), .A2(n753), .ZN(n727) );
  XNOR2_X1 U828 ( .A(n727), .B(KEYINPUT26), .ZN(n728) );
  NAND2_X1 U829 ( .A1(n728), .A2(n973), .ZN(n731) );
  NAND2_X1 U830 ( .A1(G1341), .A2(n767), .ZN(n729) );
  XNOR2_X1 U831 ( .A(KEYINPUT103), .B(n729), .ZN(n730) );
  NOR2_X1 U832 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U833 ( .A1(n733), .A2(n732), .ZN(n744) );
  NAND2_X1 U834 ( .A1(G2072), .A2(n753), .ZN(n736) );
  AND2_X1 U835 ( .A1(n767), .A2(G1956), .ZN(n737) );
  NOR2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n746) );
  AND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n742) );
  NOR2_X1 U838 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U840 ( .A1(n744), .A2(n743), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n746), .A2(n745), .ZN(n748) );
  XOR2_X1 U842 ( .A(KEYINPUT102), .B(KEYINPUT28), .Z(n747) );
  XNOR2_X1 U843 ( .A(n748), .B(n747), .ZN(n749) );
  NAND2_X1 U844 ( .A1(n750), .A2(n749), .ZN(n752) );
  XNOR2_X1 U845 ( .A(n752), .B(n751), .ZN(n757) );
  INV_X1 U846 ( .A(G1961), .ZN(n995) );
  NAND2_X1 U847 ( .A1(n767), .A2(n995), .ZN(n755) );
  XNOR2_X1 U848 ( .A(G2078), .B(KEYINPUT25), .ZN(n914) );
  NAND2_X1 U849 ( .A1(n753), .A2(n914), .ZN(n754) );
  NAND2_X1 U850 ( .A1(n755), .A2(n754), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n761), .A2(G171), .ZN(n756) );
  NAND2_X1 U852 ( .A1(n757), .A2(n756), .ZN(n766) );
  NOR2_X1 U853 ( .A1(G1966), .A2(n803), .ZN(n778) );
  NOR2_X1 U854 ( .A1(G2084), .A2(n767), .ZN(n775) );
  NOR2_X1 U855 ( .A1(n778), .A2(n775), .ZN(n758) );
  NAND2_X1 U856 ( .A1(G8), .A2(n758), .ZN(n759) );
  XNOR2_X1 U857 ( .A(KEYINPUT30), .B(n759), .ZN(n760) );
  NOR2_X1 U858 ( .A1(G168), .A2(n760), .ZN(n763) );
  NOR2_X1 U859 ( .A1(G171), .A2(n761), .ZN(n762) );
  NOR2_X1 U860 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U861 ( .A(KEYINPUT31), .B(n764), .Z(n765) );
  NAND2_X1 U862 ( .A1(n766), .A2(n765), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n776), .A2(G286), .ZN(n772) );
  NOR2_X1 U864 ( .A1(G1971), .A2(n803), .ZN(n769) );
  NOR2_X1 U865 ( .A1(G2090), .A2(n767), .ZN(n768) );
  NOR2_X1 U866 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U867 ( .A1(n770), .A2(G303), .ZN(n771) );
  NAND2_X1 U868 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U869 ( .A1(n773), .A2(G8), .ZN(n774) );
  XNOR2_X1 U870 ( .A(KEYINPUT32), .B(n774), .ZN(n793) );
  NAND2_X1 U871 ( .A1(G8), .A2(n775), .ZN(n780) );
  INV_X1 U872 ( .A(n776), .ZN(n777) );
  NOR2_X1 U873 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n794) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n966) );
  AND2_X1 U876 ( .A1(n794), .A2(n966), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n793), .A2(n781), .ZN(n785) );
  INV_X1 U878 ( .A(n966), .ZN(n783) );
  NOR2_X1 U879 ( .A1(G1976), .A2(G288), .ZN(n788) );
  NOR2_X1 U880 ( .A1(G1971), .A2(G303), .ZN(n782) );
  NOR2_X1 U881 ( .A1(n788), .A2(n782), .ZN(n967) );
  OR2_X1 U882 ( .A1(n783), .A2(n967), .ZN(n784) );
  AND2_X1 U883 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U884 ( .A1(n803), .A2(n786), .ZN(n787) );
  NOR2_X1 U885 ( .A1(KEYINPUT33), .A2(n787), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n788), .A2(KEYINPUT33), .ZN(n789) );
  NOR2_X1 U887 ( .A1(n789), .A2(n803), .ZN(n790) );
  NOR2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U889 ( .A(G1981), .B(G305), .Z(n955) );
  NAND2_X1 U890 ( .A1(n792), .A2(n955), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n797) );
  NOR2_X1 U892 ( .A1(G2090), .A2(G303), .ZN(n795) );
  NAND2_X1 U893 ( .A1(G8), .A2(n795), .ZN(n796) );
  NAND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U895 ( .A1(n798), .A2(n803), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n805) );
  NOR2_X1 U897 ( .A1(G1981), .A2(G305), .ZN(n801) );
  XOR2_X1 U898 ( .A(n801), .B(KEYINPUT24), .Z(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n823) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n880), .ZN(n933) );
  NOR2_X1 U904 ( .A1(n888), .A2(G1991), .ZN(n810) );
  XNOR2_X1 U905 ( .A(n810), .B(KEYINPUT104), .ZN(n929) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n929), .A2(n811), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n933), .A2(n814), .ZN(n815) );
  XNOR2_X1 U910 ( .A(KEYINPUT39), .B(n815), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n818), .A2(n892), .ZN(n937) );
  NAND2_X1 U913 ( .A1(n819), .A2(n937), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n824), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U919 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  NOR2_X1 U927 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U929 ( .A(G1991), .B(G2474), .ZN(n840) );
  XOR2_X1 U930 ( .A(G1981), .B(G1966), .Z(n832) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1986), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U933 ( .A(G1976), .B(G1971), .Z(n834) );
  XNOR2_X1 U934 ( .A(G1961), .B(G1956), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(G229) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2072), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n841), .B(KEYINPUT107), .ZN(n851) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(KEYINPUT43), .Z(n843) );
  XNOR2_X1 U943 ( .A(G2678), .B(G2096), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U945 ( .A(G2100), .B(G2090), .Z(n845) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2084), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U948 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U949 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G227) );
  NAND2_X1 U952 ( .A1(G124), .A2(n871), .ZN(n852) );
  XOR2_X1 U953 ( .A(KEYINPUT111), .B(n852), .Z(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G100), .A2(n867), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G112), .A2(n872), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G136), .A2(n868), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U960 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U961 ( .A1(G130), .A2(n871), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G118), .A2(n872), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G106), .A2(n867), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G142), .A2(n868), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U967 ( .A(KEYINPUT45), .B(n864), .Z(n865) );
  NOR2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n882) );
  NAND2_X1 U969 ( .A1(G103), .A2(n867), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G139), .A2(n868), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G127), .A2(n871), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G115), .A2(n872), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(n875), .ZN(n876) );
  XNOR2_X1 U976 ( .A(KEYINPUT113), .B(n876), .ZN(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n943) );
  XOR2_X1 U978 ( .A(G164), .B(n943), .Z(n879) );
  XNOR2_X1 U979 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(n882), .B(n881), .Z(n884) );
  XNOR2_X1 U981 ( .A(G160), .B(n927), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n894) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n886) );
  XNOR2_X1 U984 ( .A(G162), .B(KEYINPUT114), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(KEYINPUT46), .B(n887), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n888), .B(KEYINPUT115), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n973), .B(G286), .ZN(n897) );
  XNOR2_X1 U993 ( .A(G171), .B(n958), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U995 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U996 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U997 ( .A(KEYINPUT106), .B(n901), .Z(G319) );
  NOR2_X1 U998 ( .A1(G229), .A2(G227), .ZN(n902) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n902), .ZN(n903) );
  NOR2_X1 U1000 ( .A1(G401), .A2(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n904) );
  AND2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n906), .A2(G319), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1005 ( .A(G2090), .B(G35), .ZN(n919) );
  XNOR2_X1 U1006 ( .A(G2067), .B(G26), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(G33), .B(G2072), .ZN(n907) );
  NOR2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n913) );
  XOR2_X1 U1009 ( .A(G1991), .B(G25), .Z(n909) );
  NAND2_X1 U1010 ( .A1(n909), .A2(G28), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(G32), .B(G1996), .ZN(n910) );
  NOR2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n916) );
  XOR2_X1 U1014 ( .A(G27), .B(n914), .Z(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT53), .B(n917), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n922) );
  XOR2_X1 U1018 ( .A(G2084), .B(KEYINPUT54), .Z(n920) );
  XNOR2_X1 U1019 ( .A(G34), .B(n920), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT119), .B(n923), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G29), .A2(n924), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT55), .ZN(n953) );
  XOR2_X1 U1024 ( .A(G2084), .B(G160), .Z(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(n934), .B(KEYINPUT51), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT116), .B(n941), .ZN(n949) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT118), .B(n942), .ZN(n946) );
  XOR2_X1 U1037 ( .A(n943), .B(KEYINPUT117), .Z(n944) );
  XOR2_X1 U1038 ( .A(G2072), .B(n944), .Z(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT50), .B(n947), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(n950), .ZN(n951) );
  NAND2_X1 U1043 ( .A1(G29), .A2(n951), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n1010) );
  INV_X1 U1045 ( .A(G16), .ZN(n1005) );
  XOR2_X1 U1046 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n954) );
  XNOR2_X1 U1047 ( .A(n1005), .B(n954), .ZN(n979) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G168), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(KEYINPUT57), .ZN(n977) );
  XNOR2_X1 U1051 ( .A(G1348), .B(n958), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(G171), .B(G1961), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n972) );
  XNOR2_X1 U1055 ( .A(G299), .B(G1956), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(n963), .B(KEYINPUT121), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(G1971), .A2(G303), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(n970), .B(KEYINPUT122), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1063 ( .A(G1341), .B(n973), .Z(n974) );
  NOR2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1065 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1066 ( .A1(n979), .A2(n978), .ZN(n1007) );
  XOR2_X1 U1067 ( .A(G1986), .B(G24), .Z(n982) );
  XNOR2_X1 U1068 ( .A(G23), .B(KEYINPUT125), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n980), .B(G1976), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(n982), .A2(n981), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(G22), .B(G1971), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1073 ( .A(KEYINPUT58), .B(n985), .Z(n1002) );
  XOR2_X1 U1074 ( .A(G20), .B(G1956), .Z(n989) );
  XNOR2_X1 U1075 ( .A(G1341), .B(G19), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G6), .B(G1981), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n993) );
  XNOR2_X1 U1079 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(n990), .B(G4), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n991), .B(G1348), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n994), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(n995), .B(G5), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G21), .B(G1966), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(KEYINPUT124), .B(n1000), .Z(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(KEYINPUT61), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(n1008), .B(KEYINPUT126), .ZN(n1009) );
  NOR2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1095 ( .A1(n1011), .A2(G11), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1012), .B(KEYINPUT127), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(KEYINPUT62), .B(n1013), .ZN(G311) );
  INV_X1 U1098 ( .A(G311), .ZN(G150) );
endmodule

