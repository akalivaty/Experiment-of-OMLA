//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT68), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G218), .A3(G220), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT70), .Z(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT71), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI21_X1  g034(.A(KEYINPUT72), .B1(new_n454), .B2(G2106), .ZN(new_n460));
  AND3_X1   g035(.A1(new_n454), .A2(KEYINPUT72), .A3(G2106), .ZN(new_n461));
  AOI211_X1 g036(.A(new_n460), .B(new_n461), .C1(G567), .C2(new_n457), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT74), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n466), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(KEYINPUT73), .A2(G113), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n463), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n471), .A2(new_n472), .A3(new_n479), .ZN(G160));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n464), .A2(new_n465), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n463), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n484), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT75), .Z(G162));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n464), .B2(new_n465), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(KEYINPUT76), .B(new_n495), .C1(new_n464), .C2(new_n465), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n481), .A2(new_n503), .A3(G138), .A4(new_n463), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI211_X1 g084(.A(G50), .B(G543), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n511), .A2(new_n512), .B1(new_n508), .B2(new_n509), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(G62), .B1(new_n512), .B2(new_n511), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT77), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n518), .ZN(new_n525));
  OAI21_X1  g100(.A(G651), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT77), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(new_n529), .A3(G88), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n526), .A2(new_n527), .A3(new_n530), .A4(new_n510), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n520), .A2(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n529), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n512), .A2(new_n511), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n529), .A2(G89), .ZN(new_n539));
  NAND2_X1  g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n537), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n516), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n548), .B1(new_n547), .B2(new_n546), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n529), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n513), .ZN(new_n551));
  AOI22_X1  g126(.A1(G52), .A2(new_n550), .B1(new_n551), .B2(G90), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  AOI22_X1  g129(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n516), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n535), .A2(new_n557), .B1(new_n513), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT79), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n538), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(G651), .A2(new_n569), .B1(new_n551), .B2(G91), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n535), .C2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(KEYINPUT80), .B2(KEYINPUT9), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n550), .B(new_n575), .C1(KEYINPUT80), .C2(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n570), .A2(new_n574), .A3(new_n576), .ZN(G299));
  AND3_X1   g152(.A1(new_n520), .A2(KEYINPUT81), .A3(new_n531), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT81), .B1(new_n520), .B2(new_n531), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G303));
  NAND2_X1  g155(.A1(new_n550), .A2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n551), .A2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n538), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G73), .ZN(new_n587));
  INV_X1    g162(.A(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n551), .A2(G86), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n529), .A2(G48), .A3(G543), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(G47), .A2(new_n550), .B1(new_n551), .B2(G85), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n516), .B2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n551), .A2(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n550), .A2(KEYINPUT82), .ZN(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n535), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n538), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n601), .A2(new_n604), .B1(G651), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n597), .B1(new_n610), .B2(G868), .ZN(G284));
  XNOR2_X1  g186(.A(G284), .B(KEYINPUT83), .ZN(G321));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(G299), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(G168), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(new_n613), .B2(G168), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  OR2_X1    g193(.A1(new_n556), .A2(new_n559), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n613), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n609), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n481), .A2(new_n469), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT84), .B(G2100), .Z(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n483), .A2(G123), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n486), .A2(G135), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n463), .A2(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n628), .A2(new_n629), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT86), .Z(new_n653));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n650), .B2(new_n651), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(G401));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(G2100), .Z(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n635), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  INV_X1    g251(.A(new_n671), .ZN(new_n677));
  INV_X1    g252(.A(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n673), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n680), .C1(new_n677), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT89), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n683), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G35), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT98), .Z(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G162), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT29), .ZN(new_n695));
  INV_X1    g270(.A(G2090), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n486), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n483), .A2(G129), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT26), .Z(new_n701));
  NAND3_X1  g276(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT95), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT95), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G29), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(KEYINPUT96), .C1(G29), .C2(G32), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(KEYINPUT96), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G4), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n610), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT24), .ZN(new_n714));
  INV_X1    g289(.A(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G160), .B2(new_n691), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n713), .A2(G1348), .B1(G2084), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  NOR2_X1   g295(.A1(G171), .A2(new_n711), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G5), .B2(new_n711), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n719), .B1(G1348), .B2(new_n713), .C1(new_n720), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n711), .A2(G19), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n560), .B2(new_n711), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1341), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n691), .A2(G33), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n486), .A2(G139), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT25), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G127), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n463), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n727), .B1(new_n736), .B2(new_n691), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT94), .B(G2072), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n711), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n711), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G1966), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT31), .B(G11), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT97), .B(G28), .Z(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n744), .B2(KEYINPUT30), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT30), .B2(new_n744), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n743), .B(new_n746), .C1(new_n634), .C2(new_n691), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n741), .B2(G1966), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n726), .A2(new_n739), .A3(new_n742), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G164), .A2(new_n691), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G27), .B2(new_n691), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n691), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n483), .A2(G128), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n486), .A2(G140), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(new_n691), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n753), .A2(new_n754), .A3(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n723), .A2(new_n749), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n718), .A2(G2084), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n711), .A2(G20), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT23), .Z(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G299), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1956), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n768), .B(new_n773), .C1(new_n720), .C2(new_n722), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n697), .A2(new_n710), .A3(new_n767), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT99), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n711), .A2(G22), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT92), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n711), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT93), .Z(new_n780));
  INV_X1    g355(.A(G1971), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  MUX2_X1   g358(.A(G6), .B(G305), .S(G16), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT32), .B(G1981), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n711), .A2(G23), .ZN(new_n787));
  INV_X1    g362(.A(G288), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n711), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT33), .B(G1976), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT91), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n782), .A2(new_n783), .A3(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n691), .A2(G25), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n483), .A2(G119), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n486), .A2(G131), .ZN(new_n799));
  OR2_X1    g374(.A1(G95), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n691), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT90), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G1991), .Z(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  MUX2_X1   g384(.A(G24), .B(G290), .S(G16), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1986), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n795), .A2(new_n796), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT36), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n776), .A2(new_n814), .ZN(G311));
  NAND2_X1  g390(.A1(new_n776), .A2(new_n814), .ZN(G150));
  AOI22_X1  g391(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n516), .ZN(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n535), .A2(new_n819), .B1(new_n513), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT37), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n609), .A2(new_n617), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n818), .A2(new_n821), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n619), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n560), .A2(new_n822), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n828), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n823), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n825), .B1(new_n836), .B2(new_n837), .ZN(G145));
  NAND2_X1  g413(.A1(new_n705), .A2(new_n761), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n761), .B1(new_n703), .B2(new_n704), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(G164), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n703), .A2(new_n704), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(new_n762), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n506), .B1(new_n844), .B2(new_n840), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n736), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT102), .B1(new_n847), .B2(KEYINPUT101), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(KEYINPUT102), .B2(new_n847), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n842), .A2(new_n845), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n483), .A2(G130), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n463), .A2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G142), .B2(new_n486), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n625), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n803), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n634), .B(G160), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  INV_X1    g437(.A(new_n859), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n849), .A2(new_n863), .A3(new_n851), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n860), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT103), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n860), .A2(new_n867), .A3(new_n862), .A4(new_n864), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n862), .B1(new_n860), .B2(new_n864), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(G37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n621), .B(new_n833), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n609), .A2(G299), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n609), .A2(G299), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n621), .B(new_n832), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n876), .A2(KEYINPUT41), .A3(new_n877), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT41), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n874), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(G290), .B(G305), .Z(new_n886));
  NOR2_X1   g461(.A1(G166), .A2(new_n788), .ZN(new_n887));
  AOI21_X1  g462(.A(G288), .B1(new_n531), .B2(new_n520), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n886), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n879), .A2(new_n883), .A3(new_n874), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n885), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n892), .B1(new_n896), .B2(new_n884), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n897), .A3(G868), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT105), .B1(new_n829), .B2(new_n613), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n895), .A2(new_n897), .A3(KEYINPUT105), .A4(G868), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(G295));
  AND3_X1   g477(.A1(new_n900), .A2(KEYINPUT106), .A3(new_n901), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT106), .B1(new_n900), .B2(new_n901), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(G331));
  XNOR2_X1  g480(.A(new_n832), .B(G301), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G168), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n832), .B(G171), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G286), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n878), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n881), .A2(new_n882), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n907), .A3(new_n909), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n890), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n890), .B1(new_n912), .B2(new_n914), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT107), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(KEYINPUT43), .C1(new_n917), .C2(new_n918), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n915), .A2(new_n916), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n918), .A2(new_n925), .ZN(new_n926));
  AOI211_X1 g501(.A(KEYINPUT108), .B(new_n890), .C1(new_n912), .C2(new_n914), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n923), .B(new_n924), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n920), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n924), .B1(new_n917), .B2(new_n918), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n924), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT44), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n935), .ZN(G397));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n506), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n472), .ZN(new_n941));
  INV_X1    g516(.A(new_n479), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n941), .A2(new_n942), .A3(G40), .A4(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1996), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n761), .B(new_n764), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n843), .A2(G1996), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n803), .A2(new_n807), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n803), .A2(new_n807), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(G290), .B(G1986), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n945), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT116), .ZN(new_n957));
  AOI21_X1  g532(.A(G1384), .B1(new_n500), .B2(new_n505), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n957), .A3(new_n959), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n944), .B1(new_n938), .B2(KEYINPUT50), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n772), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT121), .ZN(new_n966));
  OR3_X1    g541(.A1(G299), .A2(new_n966), .A3(KEYINPUT57), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(KEYINPUT57), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n966), .A2(KEYINPUT57), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(G299), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n958), .A2(KEYINPUT45), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n939), .B(G1384), .C1(new_n500), .C2(new_n505), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n974), .A2(new_n975), .A3(new_n944), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT56), .B(G2072), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n965), .A2(new_n973), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n958), .A2(new_n959), .ZN(new_n980));
  AOI21_X1  g555(.A(G1348), .B1(new_n963), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n958), .A2(G160), .A3(G40), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(G2067), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n610), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G40), .ZN(new_n987));
  NOR4_X1   g562(.A1(new_n471), .A2(new_n472), .A3(new_n479), .A4(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n959), .B2(new_n958), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(new_n960), .ZN(new_n990));
  AOI21_X1  g565(.A(G1956), .B1(new_n990), .B2(new_n962), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n958), .A2(KEYINPUT45), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n940), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n977), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n972), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n986), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(KEYINPUT61), .A3(new_n979), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT122), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n981), .A2(new_n983), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n609), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n984), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n609), .A2(KEYINPUT60), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n1003), .A2(KEYINPUT60), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n996), .A2(new_n979), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT61), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n982), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT58), .B(G1341), .ZN(new_n1010));
  OAI22_X1  g585(.A1(new_n993), .A2(G1996), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n560), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT59), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1005), .A2(new_n1008), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n997), .B1(new_n1000), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT126), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n788), .A2(G1976), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  AOI211_X1 g594(.A(new_n1018), .B(new_n1019), .C1(new_n988), .C2(new_n958), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT111), .B1(new_n982), .B2(G8), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT112), .ZN(new_n1023));
  OAI21_X1  g598(.A(G8), .B1(new_n938), .B2(new_n944), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1018), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n982), .A2(KEYINPUT111), .A3(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1017), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(KEYINPUT52), .A3(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT113), .B(G86), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n528), .A2(new_n529), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n589), .B1(new_n528), .B2(G61), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n592), .B(new_n1032), .C1(new_n1033), .C2(new_n516), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n590), .A2(new_n591), .A3(new_n1036), .A4(new_n592), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1035), .A2(new_n1037), .A3(KEYINPUT49), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT49), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1040), .B(KEYINPUT114), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1027), .A2(new_n1017), .A3(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1030), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n578), .A2(new_n579), .A3(new_n1019), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n993), .A2(new_n781), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n961), .A2(new_n963), .A3(new_n696), .A4(new_n962), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT117), .B(new_n1054), .C1(new_n1057), .C2(new_n1019), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1019), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1053), .B1(G303), .B2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1051), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n578), .A2(new_n579), .A3(new_n1019), .A4(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1059), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n963), .A2(new_n696), .A3(new_n980), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1055), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G8), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1067), .B1(new_n1070), .B2(new_n1054), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1019), .B1(new_n1055), .B2(new_n1068), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(new_n1064), .A3(KEYINPUT110), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1049), .A2(new_n1066), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n938), .A2(KEYINPUT50), .ZN(new_n1076));
  AOI21_X1  g651(.A(G2084), .B1(new_n958), .B2(new_n959), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n988), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n976), .B2(G1966), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1078), .B1(new_n963), .B2(new_n1077), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G286), .A2(G8), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT51), .B1(new_n1083), .B2(KEYINPUT123), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1966), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n993), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G2084), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n980), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT118), .B1(new_n1090), .B2(new_n989), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1091), .A3(new_n1079), .ZN(new_n1092));
  OAI211_X1 g667(.A(G8), .B(new_n1084), .C1(new_n1092), .C2(G286), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1083), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1086), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n993), .A2(G2078), .B1(KEYINPUT124), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(KEYINPUT124), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n976), .A2(new_n752), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n963), .A2(new_n980), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n720), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(G301), .B(KEYINPUT54), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1104), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1097), .B1(new_n993), .B2(G2078), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1097), .A2(new_n987), .A3(G2078), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n941), .A2(new_n943), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n473), .A2(new_n478), .A3(KEYINPUT125), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n473), .A2(new_n478), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n463), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1109), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(new_n940), .A3(new_n992), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1106), .A2(new_n1107), .A3(new_n1102), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1105), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1096), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1016), .B1(new_n1075), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1094), .B1(new_n1092), .B2(G8), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1121), .A2(new_n1085), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1122), .B2(new_n1093), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1072), .A2(new_n1064), .A3(KEYINPUT110), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT110), .B1(new_n1072), .B2(new_n1064), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1030), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1123), .A2(new_n1128), .A3(KEYINPUT126), .A4(new_n1066), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1015), .A2(new_n1120), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G288), .A2(G1976), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1044), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT114), .B1(new_n1027), .B2(new_n1040), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(KEYINPUT115), .A3(new_n1037), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1131), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1037), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(new_n1140), .A3(new_n1027), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1049), .A2(new_n1126), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1103), .A2(G171), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1075), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1122), .B2(new_n1093), .ZN(new_n1147));
  AND4_X1   g722(.A1(new_n1146), .A2(new_n1086), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1143), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1130), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1082), .A2(G286), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1049), .A2(new_n1074), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1070), .A2(KEYINPUT120), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1054), .B1(new_n1072), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT63), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1049), .A2(new_n1066), .A3(new_n1074), .A4(new_n1152), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1159), .A2(KEYINPUT119), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n1159), .B2(KEYINPUT119), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n956), .B1(new_n1151), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G290), .A2(G1986), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n945), .A2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT48), .Z(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n954), .B2(new_n945), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n705), .A2(new_n948), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n945), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT127), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT46), .Z(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  OAI22_X1  g749(.A1(new_n950), .A2(new_n953), .B1(G2067), .B2(new_n761), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1167), .B(new_n1174), .C1(new_n945), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1163), .A2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g752(.A(G227), .ZN(new_n1179));
  NAND3_X1  g753(.A1(G319), .A2(new_n1179), .A3(new_n689), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n653), .B2(new_n655), .ZN(new_n1181));
  NAND3_X1  g755(.A1(new_n929), .A2(new_n872), .A3(new_n1181), .ZN(G225));
  INV_X1    g756(.A(G225), .ZN(G308));
endmodule


