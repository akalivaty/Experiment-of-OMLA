//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G148gat), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(new_n207), .B2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n207), .A2(G148gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n209), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n223), .B2(KEYINPUT2), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n211), .A2(new_n214), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT74), .B(G218gat), .Z(new_n227));
  OAI211_X1 g026(.A(G211gat), .B(new_n226), .C1(new_n227), .C2(KEYINPUT22), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(KEYINPUT22), .ZN(new_n229));
  INV_X1    g028(.A(G211gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G218gat), .ZN(new_n233));
  INV_X1    g032(.A(G218gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n228), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n225), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n224), .ZN(new_n241));
  XNOR2_X1  g040(.A(G141gat), .B(G148gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n214), .B1(new_n242), .B2(KEYINPUT2), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT29), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n236), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n205), .B1(new_n240), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT3), .B1(new_n236), .B2(new_n237), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT78), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI221_X1 g052(.A(new_n204), .B1(new_n236), .B2(new_n246), .C1(new_n249), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G22gat), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G78gat), .B(G106gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT31), .B(G50gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n257), .B1(new_n248), .B2(new_n254), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(KEYINPUT85), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT85), .A4(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(G113gat), .B2(G120gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(G113gat), .A2(G120gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n276), .A2(G134gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(G134gat), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n277), .A2(new_n278), .B1(new_n270), .B2(new_n272), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n225), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(new_n279), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT80), .B1(new_n244), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n251), .A2(new_n252), .A3(new_n283), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT39), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n289), .A2(KEYINPUT88), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n244), .A2(new_n283), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT4), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n282), .A2(new_n284), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(KEYINPUT4), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n251), .A2(KEYINPUT3), .A3(new_n252), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT79), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT79), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n251), .A2(new_n297), .A3(KEYINPUT3), .A4(new_n252), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n245), .A2(new_n280), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n286), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n289), .A2(KEYINPUT88), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n290), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT39), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT83), .ZN(new_n308));
  XOR2_X1   g107(.A(G57gat), .B(G85gat), .Z(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT87), .B1(new_n306), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n312), .B(KEYINPUT86), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(new_n305), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n303), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n319), .A2(KEYINPUT40), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n286), .A2(KEYINPUT4), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n285), .A2(new_n321), .B1(KEYINPUT4), .B2(new_n291), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT5), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n285), .A2(new_n287), .ZN(new_n325));
  INV_X1    g124(.A(new_n286), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT81), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n323), .A2(KEYINPUT81), .A3(new_n327), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n326), .A2(KEYINPUT5), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n294), .A2(new_n300), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n294), .A2(new_n300), .A3(KEYINPUT84), .A4(new_n332), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n316), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n319), .B2(KEYINPUT40), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n320), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n342));
  AND3_X1   g141(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT68), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G190gat), .ZN(new_n349));
  INV_X1    g148(.A(G183gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT65), .B1(new_n352), .B2(KEYINPUT23), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n354), .B(new_n355), .C1(G169gat), .C2(G176gat), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n345), .A2(new_n351), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT66), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G169gat), .ZN(new_n363));
  INV_X1    g162(.A(G176gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT23), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT67), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n365), .B(KEYINPUT67), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n357), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT64), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n343), .B(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n344), .B1(new_n350), .B2(new_n346), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n356), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n360), .A2(new_n361), .B1(KEYINPUT23), .B2(new_n352), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n371), .A2(KEYINPUT25), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n350), .A2(KEYINPUT27), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G183gat), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n347), .A2(new_n349), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT69), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(new_n363), .A3(new_n364), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(new_n391), .C1(new_n367), .C2(new_n368), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT70), .ZN(new_n393));
  NAND2_X1  g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n392), .B2(new_n394), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n387), .B(new_n388), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n380), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G226gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(new_n203), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n342), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n380), .B2(new_n397), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n371), .A2(KEYINPUT25), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n379), .A2(new_n375), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n397), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n237), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n403), .B1(new_n407), .B2(new_n402), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n236), .B(new_n401), .C1(new_n408), .C2(new_n342), .ZN(new_n409));
  INV_X1    g208(.A(new_n236), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n400), .B1(new_n406), .B2(new_n237), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(new_n403), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G64gat), .ZN(new_n415));
  INV_X1    g214(.A(G92gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT30), .A4(new_n417), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n409), .A2(new_n417), .A3(new_n412), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT76), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n421), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n268), .B1(new_n341), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n413), .A2(KEYINPUT37), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(KEYINPUT38), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT75), .B1(new_n411), .B2(new_n403), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n434), .A2(new_n401), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n435), .B2(new_n236), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n236), .B1(new_n434), .B2(new_n401), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT89), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n408), .A2(new_n236), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT90), .B1(new_n440), .B2(KEYINPUT37), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n437), .B2(KEYINPUT89), .ZN(new_n442));
  AOI211_X1 g241(.A(new_n433), .B(new_n236), .C1(new_n434), .C2(new_n401), .ZN(new_n443));
  OAI211_X1 g242(.A(KEYINPUT90), .B(KEYINPUT37), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n432), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n418), .A2(KEYINPUT38), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n446), .A2(new_n418), .B1(new_n413), .B2(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n323), .A2(KEYINPUT81), .A3(new_n327), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n335), .B(new_n336), .C1(new_n449), .C2(new_n328), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n312), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n450), .B2(new_n312), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n413), .B(KEYINPUT37), .Z(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  OAI221_X1 g254(.A(new_n451), .B1(new_n453), .B2(new_n338), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n430), .B1(new_n448), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n380), .A2(new_n280), .A3(new_n397), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n280), .B1(new_n380), .B2(new_n397), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT71), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI211_X1 g262(.A(KEYINPUT71), .B(new_n280), .C1(new_n380), .C2(new_n397), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G43gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G71gat), .B(G99gat), .ZN(new_n472));
  XOR2_X1   g271(.A(new_n471), .B(new_n472), .Z(new_n473));
  NAND3_X1  g272(.A1(new_n466), .A2(new_n468), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n406), .A2(new_n283), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n462), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n458), .A4(new_n460), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n473), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n465), .B(KEYINPUT32), .C1(new_n467), .C2(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n474), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n482), .B2(new_n474), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n485), .A2(KEYINPUT36), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(KEYINPUT36), .ZN(new_n487));
  INV_X1    g286(.A(new_n312), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n331), .B2(new_n337), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n451), .B1(new_n453), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n428), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n486), .A2(new_n487), .B1(new_n268), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n457), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n451), .B1(new_n453), .B2(new_n338), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT35), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n494), .A2(new_n495), .A3(new_n267), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n485), .A2(KEYINPUT91), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n483), .B2(new_n484), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n496), .A2(new_n428), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT92), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n474), .A2(new_n482), .ZN(new_n502));
  INV_X1    g301(.A(new_n480), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n474), .A2(new_n480), .A3(new_n482), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n267), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n501), .B(KEYINPUT35), .C1(new_n491), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n485), .A2(new_n428), .A3(new_n490), .A4(new_n267), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n501), .B1(new_n509), .B2(KEYINPUT35), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n500), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n493), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G113gat), .B(G141gat), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT94), .ZN(new_n514));
  XOR2_X1   g313(.A(G169gat), .B(G197gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(KEYINPUT12), .Z(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g320(.A1(G29gat), .A2(G36gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT96), .Z(new_n523));
  NOR2_X1   g322(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n524));
  NOR2_X1   g323(.A1(G29gat), .A2(G36gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT14), .ZN(new_n526));
  OR4_X1    g325(.A1(new_n521), .A2(new_n523), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n526), .A2(KEYINPUT95), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n522), .B1(new_n526), .B2(KEYINPUT95), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(G1gat), .ZN(new_n534));
  AOI21_X1  g333(.A(G8gat), .B1(new_n534), .B2(KEYINPUT97), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n533), .B1(new_n536), .B2(G1gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n535), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n527), .A2(new_n530), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n532), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n531), .A2(new_n539), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n531), .B2(new_n539), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n546), .B(KEYINPUT13), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n549), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT18), .B1(new_n545), .B2(new_n546), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n519), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  INV_X1    g356(.A(new_n519), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n553), .A4(new_n547), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n512), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G176gat), .ZN(new_n564));
  INV_X1    g363(.A(G204gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G71gat), .B(G78gat), .Z(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT99), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT100), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT101), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT102), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n568), .A2(new_n569), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n575), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n573), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n584), .B2(new_n416), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G99gat), .B(G106gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n577), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT102), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(new_n573), .A3(new_n588), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G230gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n203), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT104), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n590), .B2(new_n595), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT104), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n595), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n580), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(KEYINPUT10), .A3(new_n588), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n598), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n567), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT105), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n608), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n599), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n613), .A2(new_n600), .A3(new_n566), .A4(new_n603), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n610), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n611), .B1(new_n610), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n532), .A2(new_n542), .A3(new_n589), .ZN(new_n618));
  AND2_X1   g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n540), .A2(new_n588), .B1(KEYINPUT41), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G134gat), .B(G162gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n619), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n623), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n539), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(G183gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n350), .A3(new_n539), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT103), .B(KEYINPUT21), .Z(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n607), .B2(new_n634), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n607), .A2(new_n633), .A3(new_n634), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n635), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n630), .A3(new_n631), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n230), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n637), .A2(new_n644), .A3(new_n639), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n627), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n617), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n562), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n490), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g451(.A1(new_n562), .A2(new_n429), .A3(new_n649), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT16), .B(G8gat), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT107), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n653), .B(KEYINPUT106), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n654), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(G8gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(G1325gat));
  NAND2_X1  g461(.A1(new_n486), .A2(new_n487), .ZN(new_n663));
  OAI21_X1  g462(.A(G15gat), .B1(new_n650), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n497), .A2(new_n499), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(G15gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n664), .B1(new_n650), .B2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n267), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT108), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n668), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n627), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT44), .B1(new_n512), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n627), .B(KEYINPUT110), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n511), .A2(new_n677), .B1(new_n457), .B2(new_n492), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT109), .B(new_n500), .C1(new_n508), .C2(new_n510), .ZN(new_n679));
  AOI211_X1 g478(.A(KEYINPUT111), .B(new_n676), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT111), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n511), .A2(new_n677), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n493), .A3(new_n679), .ZN(new_n683));
  INV_X1    g482(.A(new_n676), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n673), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n617), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n646), .A2(new_n647), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n561), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n490), .ZN(new_n693));
  INV_X1    g492(.A(G29gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n490), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n690), .A2(new_n672), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n562), .A2(new_n694), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT45), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n693), .A2(new_n698), .ZN(G1328gat));
  OAI21_X1  g498(.A(G36gat), .B1(new_n692), .B2(new_n428), .ZN(new_n700));
  AOI21_X1  g499(.A(G36gat), .B1(KEYINPUT112), .B2(KEYINPUT46), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n562), .A2(new_n429), .A3(new_n696), .A4(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(G1329gat));
  INV_X1    g504(.A(new_n663), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n686), .A2(new_n706), .A3(new_n691), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT113), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT113), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n686), .A2(new_n709), .A3(new_n706), .A4(new_n691), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(G43gat), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n562), .A2(new_n696), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(G43gat), .A3(new_n665), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n707), .A2(G43gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n714), .B1(new_n717), .B2(new_n713), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n692), .B2(new_n267), .ZN(new_n720));
  INV_X1    g519(.A(G50gat), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n562), .A2(new_n721), .A3(new_n268), .A4(new_n696), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n720), .A2(KEYINPUT48), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1331gat));
  AND4_X1   g526(.A1(new_n561), .A2(new_n683), .A3(new_n648), .A4(new_n687), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n695), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n429), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT49), .B(G64gat), .Z(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(G1333gat));
  NAND2_X1  g533(.A1(new_n728), .A2(new_n706), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n665), .A2(G71gat), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n735), .A2(G71gat), .B1(new_n728), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n728), .A2(new_n268), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g539(.A1(new_n688), .A2(new_n560), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n617), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n686), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G85gat), .B1(new_n744), .B2(new_n490), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n627), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT51), .B1(new_n683), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n683), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n617), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n584), .A3(new_n695), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(KEYINPUT114), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1336gat));
  NAND3_X1  g556(.A1(new_n686), .A2(new_n429), .A3(new_n743), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n686), .A2(KEYINPUT116), .A3(new_n429), .A4(new_n743), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(G92gat), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n428), .A2(G92gat), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT52), .B1(new_n751), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n758), .A2(G92gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n749), .A2(KEYINPUT115), .A3(new_n750), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n617), .B1(new_n748), .B2(new_n768), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n767), .A2(new_n763), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT52), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n771), .ZN(G1337gat));
  INV_X1    g571(.A(new_n665), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT117), .B(G99gat), .Z(new_n774));
  NAND3_X1  g573(.A1(new_n751), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n744), .A2(new_n663), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n776), .B2(new_n774), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n686), .A2(new_n268), .A3(new_n743), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT118), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n686), .A2(new_n780), .A3(new_n268), .A4(new_n743), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(G106gat), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n267), .A2(G106gat), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT53), .B1(new_n751), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n778), .A2(G106gat), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n767), .A2(new_n769), .A3(new_n783), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT53), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1339gat));
  AND3_X1   g588(.A1(new_n617), .A2(new_n648), .A3(new_n561), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n627), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n545), .A2(new_n546), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n518), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n559), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n601), .B(KEYINPUT104), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n566), .B1(new_n798), .B2(new_n613), .ZN(new_n799));
  INV_X1    g598(.A(new_n614), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT105), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n610), .A2(new_n611), .A3(new_n614), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n606), .A2(new_n608), .A3(new_n598), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n609), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n612), .A2(new_n806), .A3(new_n599), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n567), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n804), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n566), .B1(new_n609), .B2(new_n806), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n613), .A2(KEYINPUT54), .ZN(new_n812));
  OAI211_X1 g611(.A(KEYINPUT55), .B(new_n811), .C1(new_n812), .C2(new_n805), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n560), .A2(new_n810), .A3(new_n614), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n793), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n797), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n810), .A2(new_n614), .A3(new_n813), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n674), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n791), .B1(new_n819), .B2(new_n688), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n695), .ZN(new_n821));
  INV_X1    g620(.A(new_n506), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n428), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n561), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n429), .A2(new_n490), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n820), .A2(new_n267), .A3(new_n773), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n560), .A2(G113gat), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n824), .A2(G113gat), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT119), .ZN(G1340gat));
  NOR2_X1   g628(.A1(new_n823), .A2(new_n617), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n687), .A2(G120gat), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n830), .A2(G120gat), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT120), .Z(G1341gat));
  INV_X1    g632(.A(new_n688), .ZN(new_n834));
  OAI21_X1  g633(.A(G127gat), .B1(new_n826), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n688), .A2(new_n276), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n823), .B2(new_n836), .ZN(G1342gat));
  NAND2_X1  g636(.A1(new_n428), .A2(new_n627), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(G134gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n822), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n826), .B2(new_n672), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  NAND4_X1  g643(.A1(new_n820), .A2(new_n695), .A3(new_n268), .A4(new_n663), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n429), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n561), .A2(G141gat), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n663), .A2(new_n825), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT57), .B1(new_n820), .B2(new_n268), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n672), .B1(new_n803), .B2(new_n814), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n818), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n790), .B1(new_n852), .B2(new_n834), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n854), .A3(new_n267), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n849), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G141gat), .B1(new_n856), .B2(new_n561), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n848), .A2(KEYINPUT121), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(G148gat), .C1(new_n856), .C2(new_n617), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n816), .B1(new_n615), .B2(new_n616), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n560), .A2(new_n810), .A3(new_n614), .A4(new_n813), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n627), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n672), .A2(new_n797), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n817), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n834), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n267), .B1(new_n869), .B2(new_n791), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT122), .B1(new_n870), .B2(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n867), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n790), .B1(new_n873), .B2(new_n834), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n872), .B(new_n854), .C1(new_n874), .C2(new_n267), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n267), .A2(new_n854), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n820), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n687), .A3(new_n849), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G148gat), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n862), .B1(new_n880), .B2(KEYINPUT59), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT123), .B(new_n860), .C1(new_n879), .C2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n861), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n846), .A2(new_n209), .A3(new_n687), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1345gat));
  OAI21_X1  g684(.A(G155gat), .B1(new_n856), .B2(new_n834), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n846), .A2(new_n221), .A3(new_n688), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n856), .B2(new_n793), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n428), .A2(new_n222), .A3(new_n627), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n845), .B2(new_n890), .ZN(G1347gat));
  AND2_X1   g690(.A1(new_n820), .A2(new_n490), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n892), .A2(new_n429), .A3(new_n822), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n363), .A3(new_n560), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n429), .A2(new_n490), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n665), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n820), .A2(new_n267), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n820), .A2(KEYINPUT124), .A3(new_n267), .A4(new_n896), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n560), .A3(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(G169gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(G169gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n894), .B1(new_n903), .B2(new_n904), .ZN(G1348gat));
  NAND3_X1  g704(.A1(new_n893), .A2(new_n364), .A3(new_n687), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n899), .A2(new_n687), .A3(new_n900), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n364), .ZN(G1349gat));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n893), .A2(new_n381), .A3(new_n383), .A4(new_n688), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n899), .A2(new_n688), .A3(new_n900), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G183gat), .ZN(new_n914));
  AOI211_X1 g713(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  AND4_X1   g714(.A1(new_n909), .A2(new_n912), .A3(KEYINPUT60), .A4(new_n914), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(G1350gat));
  NAND4_X1  g716(.A1(new_n893), .A2(new_n347), .A3(new_n349), .A4(new_n674), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n627), .A3(new_n900), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(G190gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n919), .B2(G190gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(G1351gat));
  NOR3_X1   g722(.A1(new_n706), .A2(new_n267), .A3(new_n428), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n892), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n560), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n706), .A2(new_n895), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n878), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n560), .A2(G197gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  NAND2_X1  g730(.A1(new_n687), .A2(new_n565), .ZN(new_n932));
  OR3_X1    g731(.A1(new_n925), .A2(KEYINPUT62), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT62), .B1(new_n925), .B2(new_n932), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n878), .A2(new_n687), .A3(new_n928), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n933), .B(new_n934), .C1(new_n935), .C2(new_n565), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n878), .A2(new_n688), .A3(new_n928), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G211gat), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n938), .A2(KEYINPUT63), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(KEYINPUT63), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n926), .A2(new_n230), .A3(new_n688), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n939), .B(new_n940), .C1(new_n943), .C2(new_n944), .ZN(G1354gat));
  AOI21_X1  g744(.A(G218gat), .B1(new_n926), .B2(new_n674), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n627), .A2(new_n227), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n929), .B2(new_n947), .ZN(G1355gat));
endmodule


