

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n571), .A2(n528), .ZN(n789) );
  XNOR2_X1 U556 ( .A(n649), .B(KEYINPUT94), .ZN(n637) );
  AND2_X2 U557 ( .A1(n726), .A2(n604), .ZN(n649) );
  INV_X1 U558 ( .A(KEYINPUT28), .ZN(n643) );
  NAND2_X1 U559 ( .A1(n653), .A2(n652), .ZN(n672) );
  XNOR2_X1 U560 ( .A(n648), .B(n647), .ZN(n653) );
  NOR2_X1 U561 ( .A1(n700), .A2(n689), .ZN(n523) );
  XNOR2_X1 U562 ( .A(n636), .B(KEYINPUT27), .ZN(n639) );
  INV_X1 U563 ( .A(KEYINPUT29), .ZN(n647) );
  AND2_X1 U564 ( .A1(n676), .A2(n675), .ZN(n677) );
  INV_X1 U565 ( .A(n748), .ZN(n737) );
  AND2_X1 U566 ( .A1(n539), .A2(G2104), .ZN(n893) );
  AND2_X1 U567 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U568 ( .A1(G651), .A2(n571), .ZN(n793) );
  NOR2_X1 U569 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U570 ( .A(KEYINPUT7), .B(n537), .Z(G168) );
  INV_X1 U571 ( .A(G651), .ZN(n528) );
  NOR2_X1 U572 ( .A1(G543), .A2(n528), .ZN(n524) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n524), .Z(n786) );
  NAND2_X1 U574 ( .A1(G63), .A2(n786), .ZN(n526) );
  XOR2_X1 U575 ( .A(KEYINPUT0), .B(G543), .Z(n571) );
  NAND2_X1 U576 ( .A1(G51), .A2(n793), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U578 ( .A(KEYINPUT6), .B(n527), .ZN(n535) );
  NAND2_X1 U579 ( .A1(n789), .A2(G76), .ZN(n529) );
  XNOR2_X1 U580 ( .A(KEYINPUT74), .B(n529), .ZN(n532) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n785) );
  NAND2_X1 U582 ( .A1(n785), .A2(G89), .ZN(n530) );
  XNOR2_X1 U583 ( .A(KEYINPUT4), .B(n530), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U585 ( .A(n533), .B(KEYINPUT5), .Z(n534) );
  XOR2_X1 U586 ( .A(KEYINPUT75), .B(n536), .Z(n537) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT17), .B(n538), .Z(n894) );
  NAND2_X1 U589 ( .A1(n894), .A2(G138), .ZN(n542) );
  INV_X1 U590 ( .A(G2105), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G102), .A2(n893), .ZN(n540) );
  XOR2_X1 U592 ( .A(KEYINPUT87), .B(n540), .Z(n541) );
  NAND2_X1 U593 ( .A1(n542), .A2(n541), .ZN(n548) );
  INV_X1 U594 ( .A(G2105), .ZN(n543) );
  NOR2_X2 U595 ( .A1(G2104), .A2(n543), .ZN(n897) );
  NAND2_X1 U596 ( .A1(n897), .A2(G126), .ZN(n546) );
  NAND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n544) );
  XOR2_X1 U598 ( .A(KEYINPUT66), .B(n544), .Z(n898) );
  NAND2_X1 U599 ( .A1(G114), .A2(n898), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U601 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U602 ( .A1(G91), .A2(n785), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G78), .A2(n789), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U605 ( .A1(G65), .A2(n786), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G53), .A2(n793), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U609 ( .A(KEYINPUT68), .B(n555), .Z(G299) );
  NAND2_X1 U610 ( .A1(G64), .A2(n786), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G52), .A2(n793), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U613 ( .A(KEYINPUT67), .B(n558), .Z(n563) );
  NAND2_X1 U614 ( .A1(G90), .A2(n785), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G77), .A2(n789), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U618 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U619 ( .A1(G88), .A2(n785), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G75), .A2(n789), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U622 ( .A1(G62), .A2(n786), .ZN(n567) );
  NAND2_X1 U623 ( .A1(G50), .A2(n793), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U625 ( .A1(n569), .A2(n568), .ZN(G166) );
  INV_X1 U626 ( .A(G166), .ZN(G303) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(n570) );
  XNOR2_X1 U628 ( .A(KEYINPUT76), .B(n570), .ZN(G286) );
  NAND2_X1 U629 ( .A1(G87), .A2(n571), .ZN(n572) );
  XNOR2_X1 U630 ( .A(KEYINPUT81), .B(n572), .ZN(n573) );
  NOR2_X1 U631 ( .A1(n786), .A2(n573), .ZN(n575) );
  NAND2_X1 U632 ( .A1(G651), .A2(G74), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n793), .A2(G49), .ZN(n576) );
  XOR2_X1 U635 ( .A(KEYINPUT80), .B(n576), .Z(n577) );
  NOR2_X1 U636 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U637 ( .A(KEYINPUT82), .B(n579), .Z(G288) );
  NAND2_X1 U638 ( .A1(G73), .A2(n789), .ZN(n580) );
  XNOR2_X1 U639 ( .A(n580), .B(KEYINPUT2), .ZN(n587) );
  NAND2_X1 U640 ( .A1(G61), .A2(n786), .ZN(n582) );
  NAND2_X1 U641 ( .A1(G48), .A2(n793), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G86), .A2(n785), .ZN(n583) );
  XNOR2_X1 U644 ( .A(KEYINPUT83), .B(n583), .ZN(n584) );
  NOR2_X1 U645 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U647 ( .A1(G85), .A2(n785), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G72), .A2(n789), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G60), .A2(n786), .ZN(n591) );
  NAND2_X1 U651 ( .A1(G47), .A2(n793), .ZN(n590) );
  NAND2_X1 U652 ( .A1(n591), .A2(n590), .ZN(n592) );
  OR2_X1 U653 ( .A1(n593), .A2(n592), .ZN(G290) );
  NOR2_X1 U654 ( .A1(G164), .A2(G1384), .ZN(n726) );
  NAND2_X1 U655 ( .A1(G137), .A2(n894), .ZN(n595) );
  NAND2_X1 U656 ( .A1(G113), .A2(n898), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(n602) );
  NAND2_X1 U658 ( .A1(n893), .A2(G101), .ZN(n597) );
  INV_X1 U659 ( .A(KEYINPUT23), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n597), .B(n596), .ZN(n599) );
  NAND2_X1 U661 ( .A1(n897), .A2(G125), .ZN(n598) );
  NAND2_X1 U662 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U663 ( .A(KEYINPUT65), .B(n600), .Z(n601) );
  NOR2_X1 U664 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U665 ( .A(n603), .B(KEYINPUT64), .ZN(n758) );
  NAND2_X1 U666 ( .A1(n758), .A2(G40), .ZN(n725) );
  INV_X1 U667 ( .A(n725), .ZN(n604) );
  NAND2_X1 U668 ( .A1(n726), .A2(n604), .ZN(n666) );
  NOR2_X1 U669 ( .A1(G2084), .A2(n666), .ZN(n654) );
  NAND2_X1 U670 ( .A1(G8), .A2(n654), .ZN(n665) );
  NAND2_X1 U671 ( .A1(G8), .A2(n666), .ZN(n700) );
  NOR2_X1 U672 ( .A1(G1966), .A2(n700), .ZN(n663) );
  NAND2_X1 U673 ( .A1(G2067), .A2(n637), .ZN(n605) );
  XNOR2_X1 U674 ( .A(n605), .B(KEYINPUT95), .ZN(n607) );
  INV_X1 U675 ( .A(G1348), .ZN(n976) );
  NOR2_X1 U676 ( .A1(n976), .A2(n649), .ZN(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n633) );
  NAND2_X1 U678 ( .A1(G92), .A2(n785), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G79), .A2(n789), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U681 ( .A1(G66), .A2(n786), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G54), .A2(n793), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT15), .B(n614), .Z(n909) );
  NAND2_X1 U686 ( .A1(n633), .A2(n909), .ZN(n632) );
  NAND2_X1 U687 ( .A1(n786), .A2(G56), .ZN(n615) );
  XOR2_X1 U688 ( .A(KEYINPUT14), .B(n615), .Z(n621) );
  NAND2_X1 U689 ( .A1(n785), .A2(G81), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT12), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G68), .A2(n789), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U693 ( .A(KEYINPUT13), .B(n619), .Z(n620) );
  NOR2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(KEYINPUT70), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n793), .A2(G43), .ZN(n623) );
  XOR2_X1 U697 ( .A(KEYINPUT71), .B(n623), .Z(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n626), .B(KEYINPUT72), .ZN(n961) );
  AND2_X1 U700 ( .A1(n649), .A2(G1996), .ZN(n627) );
  XOR2_X1 U701 ( .A(n627), .B(KEYINPUT26), .Z(n629) );
  NAND2_X1 U702 ( .A1(n666), .A2(G1341), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U704 ( .A1(n961), .A2(n630), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n635) );
  OR2_X1 U706 ( .A1(n909), .A2(n633), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n641) );
  NAND2_X1 U708 ( .A1(G2072), .A2(n637), .ZN(n636) );
  INV_X1 U709 ( .A(G1956), .ZN(n978) );
  NOR2_X1 U710 ( .A1(n637), .A2(n978), .ZN(n638) );
  NOR2_X1 U711 ( .A1(n639), .A2(n638), .ZN(n642) );
  INV_X1 U712 ( .A(G299), .ZN(n799) );
  NAND2_X1 U713 ( .A1(n642), .A2(n799), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n646) );
  NOR2_X1 U715 ( .A1(n642), .A2(n799), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(n645) );
  NAND2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U718 ( .A(G2078), .B(KEYINPUT25), .ZN(n1002) );
  NAND2_X1 U719 ( .A1(n637), .A2(n1002), .ZN(n651) );
  OR2_X1 U720 ( .A1(G1961), .A2(n649), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n658) );
  NAND2_X1 U722 ( .A1(n658), .A2(G171), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n663), .A2(n654), .ZN(n655) );
  NAND2_X1 U724 ( .A1(G8), .A2(n655), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT30), .B(n656), .ZN(n657) );
  NOR2_X1 U726 ( .A1(G168), .A2(n657), .ZN(n660) );
  NOR2_X1 U727 ( .A1(G171), .A2(n658), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U729 ( .A(KEYINPUT31), .B(n661), .Z(n670) );
  AND2_X1 U730 ( .A1(n672), .A2(n670), .ZN(n662) );
  NOR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n684) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n700), .ZN(n668) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n666), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U736 ( .A1(n669), .A2(G303), .ZN(n673) );
  AND2_X1 U737 ( .A1(n670), .A2(n673), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n676) );
  INV_X1 U739 ( .A(n673), .ZN(n674) );
  OR2_X1 U740 ( .A1(n674), .A2(G286), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n677), .B(KEYINPUT96), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n678), .A2(G8), .ZN(n679) );
  XNOR2_X2 U743 ( .A(KEYINPUT32), .B(n679), .ZN(n686) );
  NAND2_X1 U744 ( .A1(n684), .A2(n686), .ZN(n682) );
  NOR2_X1 U745 ( .A1(G2090), .A2(G303), .ZN(n680) );
  NAND2_X1 U746 ( .A1(G8), .A2(n680), .ZN(n681) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n683), .A2(n700), .ZN(n705) );
  NAND2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n967) );
  AND2_X1 U750 ( .A1(n684), .A2(n967), .ZN(n685) );
  NAND2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n691) );
  INV_X1 U752 ( .A(n967), .ZN(n688) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n693) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n693), .A2(n687), .ZN(n968) );
  OR2_X1 U756 ( .A1(n688), .A2(n968), .ZN(n689) );
  NOR2_X1 U757 ( .A1(KEYINPUT33), .A2(n523), .ZN(n690) );
  AND2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT97), .ZN(n697) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n951) );
  NAND2_X1 U761 ( .A1(KEYINPUT33), .A2(n693), .ZN(n694) );
  OR2_X1 U762 ( .A1(n700), .A2(n694), .ZN(n695) );
  AND2_X1 U763 ( .A1(n951), .A2(n695), .ZN(n696) );
  AND2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n703) );
  NOR2_X1 U765 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XOR2_X1 U766 ( .A(n698), .B(KEYINPUT24), .Z(n699) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U768 ( .A(KEYINPUT93), .B(n701), .Z(n702) );
  NOR2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n741) );
  NAND2_X1 U771 ( .A1(n897), .A2(G119), .ZN(n707) );
  NAND2_X1 U772 ( .A1(G107), .A2(n898), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n713) );
  NAND2_X1 U774 ( .A1(n893), .A2(G95), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n708), .B(KEYINPUT88), .ZN(n710) );
  NAND2_X1 U776 ( .A1(G131), .A2(n894), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U778 ( .A(KEYINPUT89), .B(n711), .Z(n712) );
  NOR2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U780 ( .A(KEYINPUT90), .B(n714), .Z(n905) );
  NAND2_X1 U781 ( .A1(G1991), .A2(n905), .ZN(n724) );
  NAND2_X1 U782 ( .A1(G105), .A2(n893), .ZN(n715) );
  XOR2_X1 U783 ( .A(KEYINPUT38), .B(n715), .Z(n720) );
  NAND2_X1 U784 ( .A1(n897), .A2(G129), .ZN(n717) );
  NAND2_X1 U785 ( .A1(G117), .A2(n898), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U787 ( .A(KEYINPUT91), .B(n718), .Z(n719) );
  NOR2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U789 ( .A1(n894), .A2(G141), .ZN(n721) );
  NAND2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n886) );
  NAND2_X1 U791 ( .A1(G1996), .A2(n886), .ZN(n723) );
  NAND2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n940) );
  NOR2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n753) );
  NAND2_X1 U794 ( .A1(n940), .A2(n753), .ZN(n727) );
  XOR2_X1 U795 ( .A(KEYINPUT92), .B(n727), .Z(n745) );
  XOR2_X1 U796 ( .A(KEYINPUT37), .B(G2067), .Z(n750) );
  NAND2_X1 U797 ( .A1(G104), .A2(n893), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G140), .A2(n894), .ZN(n728) );
  NAND2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U800 ( .A(KEYINPUT34), .B(n730), .ZN(n735) );
  NAND2_X1 U801 ( .A1(n897), .A2(G128), .ZN(n732) );
  NAND2_X1 U802 ( .A1(G116), .A2(n898), .ZN(n731) );
  NAND2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U804 ( .A(KEYINPUT35), .B(n733), .Z(n734) );
  NOR2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U806 ( .A(KEYINPUT36), .B(n736), .Z(n883) );
  AND2_X1 U807 ( .A1(n750), .A2(n883), .ZN(n933) );
  NAND2_X1 U808 ( .A1(n753), .A2(n933), .ZN(n748) );
  NOR2_X1 U809 ( .A1(n745), .A2(n737), .ZN(n739) );
  XNOR2_X1 U810 ( .A(G1986), .B(G290), .ZN(n958) );
  NAND2_X1 U811 ( .A1(n958), .A2(n753), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n756) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n886), .ZN(n927) );
  NOR2_X1 U814 ( .A1(G1986), .A2(G290), .ZN(n743) );
  NOR2_X1 U815 ( .A1(n905), .A2(G1991), .ZN(n742) );
  XNOR2_X1 U816 ( .A(n742), .B(KEYINPUT98), .ZN(n935) );
  NOR2_X1 U817 ( .A1(n743), .A2(n935), .ZN(n744) );
  NOR2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U819 ( .A1(n927), .A2(n746), .ZN(n747) );
  XNOR2_X1 U820 ( .A(n747), .B(KEYINPUT39), .ZN(n749) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n752) );
  NOR2_X1 U822 ( .A1(n883), .A2(n750), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n751), .B(KEYINPUT99), .ZN(n943) );
  NAND2_X1 U824 ( .A1(n752), .A2(n943), .ZN(n754) );
  NAND2_X1 U825 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U826 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U827 ( .A(n757), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U828 ( .A(n758), .Z(G160) );
  AND2_X1 U829 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U830 ( .A(G132), .ZN(G219) );
  INV_X1 U831 ( .A(G82), .ZN(G220) );
  INV_X1 U832 ( .A(G57), .ZN(G237) );
  XOR2_X1 U833 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n760) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n759) );
  XNOR2_X1 U835 ( .A(n760), .B(n759), .ZN(G223) );
  INV_X1 U836 ( .A(G223), .ZN(n825) );
  NAND2_X1 U837 ( .A1(n825), .A2(G567), .ZN(n761) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(n761), .Z(G234) );
  INV_X1 U839 ( .A(G860), .ZN(n767) );
  OR2_X1 U840 ( .A1(n767), .A2(n961), .ZN(G153) );
  NAND2_X1 U841 ( .A1(G868), .A2(G171), .ZN(n763) );
  INV_X1 U842 ( .A(G868), .ZN(n807) );
  NAND2_X1 U843 ( .A1(n909), .A2(n807), .ZN(n762) );
  NAND2_X1 U844 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U845 ( .A(n764), .B(KEYINPUT73), .ZN(G284) );
  NAND2_X1 U846 ( .A1(G868), .A2(G286), .ZN(n766) );
  NAND2_X1 U847 ( .A1(G299), .A2(n807), .ZN(n765) );
  NAND2_X1 U848 ( .A1(n766), .A2(n765), .ZN(G297) );
  NAND2_X1 U849 ( .A1(n767), .A2(G559), .ZN(n768) );
  NAND2_X1 U850 ( .A1(n768), .A2(n909), .ZN(n769) );
  XNOR2_X1 U851 ( .A(n769), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U852 ( .A1(n961), .A2(G868), .ZN(n772) );
  NAND2_X1 U853 ( .A1(G868), .A2(n909), .ZN(n770) );
  NOR2_X1 U854 ( .A1(G559), .A2(n770), .ZN(n771) );
  NOR2_X1 U855 ( .A1(n772), .A2(n771), .ZN(G282) );
  NAND2_X1 U856 ( .A1(G123), .A2(n897), .ZN(n773) );
  XOR2_X1 U857 ( .A(KEYINPUT18), .B(n773), .Z(n774) );
  XNOR2_X1 U858 ( .A(n774), .B(KEYINPUT77), .ZN(n776) );
  NAND2_X1 U859 ( .A1(G99), .A2(n893), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U861 ( .A1(G135), .A2(n894), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G111), .A2(n898), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n932) );
  XNOR2_X1 U865 ( .A(G2096), .B(n932), .ZN(n782) );
  INV_X1 U866 ( .A(G2100), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(G156) );
  NAND2_X1 U868 ( .A1(G559), .A2(n909), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT78), .ZN(n805) );
  XNOR2_X1 U870 ( .A(n961), .B(n805), .ZN(n784) );
  NOR2_X1 U871 ( .A1(G860), .A2(n784), .ZN(n796) );
  NAND2_X1 U872 ( .A1(G93), .A2(n785), .ZN(n788) );
  NAND2_X1 U873 ( .A1(G67), .A2(n786), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G80), .A2(n789), .ZN(n790) );
  XNOR2_X1 U876 ( .A(KEYINPUT79), .B(n790), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U878 ( .A1(n793), .A2(G55), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n808) );
  XOR2_X1 U880 ( .A(n796), .B(n808), .Z(G145) );
  XOR2_X1 U881 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n798) );
  XNOR2_X1 U882 ( .A(G288), .B(G166), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n798), .B(n797), .ZN(n800) );
  XNOR2_X1 U884 ( .A(n800), .B(n799), .ZN(n801) );
  XNOR2_X1 U885 ( .A(n801), .B(n808), .ZN(n802) );
  XNOR2_X1 U886 ( .A(n802), .B(G290), .ZN(n803) );
  XNOR2_X1 U887 ( .A(n803), .B(G305), .ZN(n804) );
  XNOR2_X1 U888 ( .A(n961), .B(n804), .ZN(n911) );
  XNOR2_X1 U889 ( .A(n805), .B(n911), .ZN(n806) );
  NOR2_X1 U890 ( .A1(n807), .A2(n806), .ZN(n810) );
  NOR2_X1 U891 ( .A1(G868), .A2(n808), .ZN(n809) );
  NOR2_X1 U892 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U893 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U894 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U895 ( .A1(G2090), .A2(n812), .ZN(n813) );
  XNOR2_X1 U896 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U897 ( .A1(n814), .A2(G2072), .ZN(G158) );
  XOR2_X1 U898 ( .A(KEYINPUT85), .B(G44), .Z(n815) );
  XNOR2_X1 U899 ( .A(KEYINPUT3), .B(n815), .ZN(G218) );
  NAND2_X1 U900 ( .A1(G120), .A2(G69), .ZN(n816) );
  NOR2_X1 U901 ( .A1(G237), .A2(n816), .ZN(n817) );
  XNOR2_X1 U902 ( .A(KEYINPUT86), .B(n817), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n818), .A2(G108), .ZN(n831) );
  NAND2_X1 U904 ( .A1(G567), .A2(n831), .ZN(n823) );
  NOR2_X1 U905 ( .A1(G220), .A2(G219), .ZN(n819) );
  XOR2_X1 U906 ( .A(KEYINPUT22), .B(n819), .Z(n820) );
  NOR2_X1 U907 ( .A1(G218), .A2(n820), .ZN(n821) );
  NAND2_X1 U908 ( .A1(G96), .A2(n821), .ZN(n832) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n832), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n823), .A2(n822), .ZN(n844) );
  NAND2_X1 U911 ( .A1(G661), .A2(G483), .ZN(n824) );
  NOR2_X1 U912 ( .A1(n844), .A2(n824), .ZN(n830) );
  NAND2_X1 U913 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U914 ( .A1(n825), .A2(G2106), .ZN(n826) );
  XNOR2_X1 U915 ( .A(n826), .B(KEYINPUT102), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U917 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT103), .B(n828), .Z(n829) );
  NAND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G108), .ZN(G238) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U928 ( .A(G2430), .B(G2454), .ZN(n841) );
  XNOR2_X1 U929 ( .A(KEYINPUT100), .B(G2435), .ZN(n839) );
  XOR2_X1 U930 ( .A(G2451), .B(G2427), .Z(n834) );
  XNOR2_X1 U931 ( .A(G2438), .B(G2446), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n835), .B(G2443), .Z(n837) );
  XNOR2_X1 U934 ( .A(G1348), .B(G1341), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n842), .A2(G14), .ZN(n843) );
  XNOR2_X1 U939 ( .A(KEYINPUT101), .B(n843), .ZN(G401) );
  XOR2_X1 U940 ( .A(KEYINPUT104), .B(n844), .Z(G319) );
  XNOR2_X1 U941 ( .A(G1981), .B(KEYINPUT41), .ZN(n854) );
  XOR2_X1 U942 ( .A(G1956), .B(G1971), .Z(n846) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1976), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(G1961), .B(G1966), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1991), .B(G1996), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U949 ( .A(KEYINPUT106), .B(G2474), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT105), .B(G2090), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2072), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(n857), .B(G2096), .Z(n859) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2084), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U958 ( .A(KEYINPUT43), .B(G2678), .Z(n861) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(G2100), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U961 ( .A(n863), .B(n862), .Z(G227) );
  NAND2_X1 U962 ( .A1(G100), .A2(n893), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G136), .A2(n894), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n898), .A2(G112), .ZN(n866) );
  XOR2_X1 U966 ( .A(KEYINPUT108), .B(n866), .Z(n867) );
  NOR2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n870) );
  NAND2_X1 U969 ( .A1(G124), .A2(n897), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT109), .ZN(G162) );
  XNOR2_X1 U973 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G106), .A2(n893), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G142), .A2(n894), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n876), .B(KEYINPUT45), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n897), .A2(G130), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G118), .A2(n898), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n883), .B(G164), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n890) );
  XNOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n886), .B(KEYINPUT112), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n892) );
  XNOR2_X1 U989 ( .A(G160), .B(n932), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n904) );
  NAND2_X1 U991 ( .A1(G103), .A2(n893), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G139), .A2(n894), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U994 ( .A1(n897), .A2(G127), .ZN(n900) );
  NAND2_X1 U995 ( .A1(G115), .A2(n898), .ZN(n899) );
  NAND2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n922) );
  XOR2_X1 U999 ( .A(n904), .B(n922), .Z(n907) );
  XNOR2_X1 U1000 ( .A(n905), .B(G162), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n908), .ZN(G395) );
  INV_X1 U1003 ( .A(n909), .ZN(n954) );
  XNOR2_X1 U1004 ( .A(G171), .B(n954), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n910), .B(G286), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n913), .ZN(G397) );
  INV_X1 U1008 ( .A(G401), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(n914), .A2(G319), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n915) );
  XOR2_X1 U1011 ( .A(KEYINPUT49), .B(n915), .Z(n916) );
  XNOR2_X1 U1012 ( .A(n916), .B(KEYINPUT113), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U1018 ( .A(G164), .B(G2078), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n921), .B(KEYINPUT117), .ZN(n924) );
  XOR2_X1 U1020 ( .A(G2072), .B(n922), .Z(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT50), .B(n925), .ZN(n931) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1025 ( .A(KEYINPUT116), .B(n928), .Z(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT51), .B(n929), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n945) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G2084), .B(KEYINPUT114), .Z(n934) );
  XNOR2_X1 U1030 ( .A(G160), .B(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1034 ( .A(KEYINPUT115), .B(n941), .Z(n942) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n946), .ZN(n948) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1040 ( .A1(n949), .A2(G29), .ZN(n1037) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G168), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(n950), .B(KEYINPUT120), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(n953), .B(KEYINPUT57), .ZN(n966) );
  XNOR2_X1 U1045 ( .A(G301), .B(G1961), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(n954), .B(G1348), .ZN(n955) );
  NOR2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n960) );
  XNOR2_X1 U1048 ( .A(G1956), .B(G299), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n964) );
  XNOR2_X1 U1051 ( .A(G1341), .B(n961), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n962), .ZN(n963) );
  NOR2_X1 U1053 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1054 ( .A1(n966), .A2(n965), .ZN(n973) );
  AND2_X1 U1055 ( .A1(G303), .A2(G1971), .ZN(n970) );
  NAND2_X1 U1056 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1057 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1058 ( .A(KEYINPUT121), .B(n971), .ZN(n972) );
  NOR2_X1 U1059 ( .A1(n973), .A2(n972), .ZN(n1026) );
  NOR2_X1 U1060 ( .A1(KEYINPUT56), .A2(n1026), .ZN(n1000) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G21), .ZN(n975) );
  XNOR2_X1 U1062 ( .A(G5), .B(G1961), .ZN(n974) );
  NOR2_X1 U1063 ( .A1(n975), .A2(n974), .ZN(n996) );
  XNOR2_X1 U1064 ( .A(KEYINPUT59), .B(G4), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(n977), .B(n976), .ZN(n985) );
  XOR2_X1 U1066 ( .A(G1341), .B(G19), .Z(n980) );
  XNOR2_X1 U1067 ( .A(n978), .B(G20), .ZN(n979) );
  NAND2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(G6), .B(G1981), .ZN(n981) );
  NOR2_X1 U1070 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1071 ( .A(KEYINPUT124), .B(n983), .Z(n984) );
  NOR2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(n986), .B(KEYINPUT125), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(n987), .B(KEYINPUT60), .ZN(n994) );
  XNOR2_X1 U1075 ( .A(G1976), .B(G23), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G1971), .B(G22), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n991) );
  XOR2_X1 U1078 ( .A(G1986), .B(G24), .Z(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n992), .ZN(n993) );
  NOR2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(n997), .B(KEYINPUT126), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(KEYINPUT61), .B(n998), .ZN(n1024) );
  NOR2_X1 U1085 ( .A1(n1024), .A2(KEYINPUT123), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1087 ( .A1(G16), .A2(n1001), .ZN(n1034) );
  XNOR2_X1 U1088 ( .A(G27), .B(n1002), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(G2067), .B(G26), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(G1996), .B(G32), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G33), .B(G2072), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(KEYINPUT118), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1096 ( .A(G1991), .B(G25), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(G28), .A2(n1012), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1013), .B(KEYINPUT53), .ZN(n1016) );
  XOR2_X1 U1100 ( .A(G2084), .B(G34), .Z(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT54), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(G35), .B(G2090), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT55), .B(n1019), .ZN(n1021) );
  INV_X1 U1106 ( .A(G29), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(G11), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(n1023), .B(KEYINPUT119), .ZN(n1032) );
  INV_X1 U1110 ( .A(n1024), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(KEYINPUT123), .A2(n1025), .ZN(n1029) );
  INV_X1 U1112 ( .A(n1026), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(KEYINPUT56), .A2(n1027), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(G16), .A2(n1030), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1118 ( .A(KEYINPUT127), .B(n1035), .Z(n1036) );
  NAND2_X1 U1119 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1038), .Z(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

