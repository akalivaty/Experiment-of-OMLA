

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U322 ( .A(n570), .B(KEYINPUT41), .Z(n543) );
  XNOR2_X1 U323 ( .A(n326), .B(KEYINPUT46), .ZN(n327) );
  XNOR2_X1 U324 ( .A(n328), .B(n327), .ZN(n346) );
  XNOR2_X1 U325 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n371) );
  XNOR2_X1 U326 ( .A(n372), .B(n371), .ZN(n523) );
  XNOR2_X1 U327 ( .A(n321), .B(n380), .ZN(n322) );
  XNOR2_X1 U328 ( .A(n323), .B(n322), .ZN(n324) );
  NOR2_X1 U329 ( .A1(n555), .A2(n564), .ZN(n448) );
  XOR2_X1 U330 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n291) );
  XNOR2_X1 U331 ( .A(KEYINPUT64), .B(KEYINPUT30), .ZN(n290) );
  XOR2_X1 U332 ( .A(n291), .B(n290), .Z(n295) );
  XOR2_X1 U333 ( .A(G43GAT), .B(G50GAT), .Z(n293) );
  XOR2_X1 U334 ( .A(G1GAT), .B(KEYINPUT68), .Z(n341) );
  XNOR2_X1 U335 ( .A(n341), .B(KEYINPUT69), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n297) );
  NAND2_X1 U338 ( .A1(G229GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U340 ( .A(G197GAT), .B(G22GAT), .Z(n299) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G141GAT), .ZN(n298) );
  XOR2_X1 U342 ( .A(n299), .B(n298), .Z(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n309) );
  XOR2_X1 U344 ( .A(KEYINPUT67), .B(KEYINPUT8), .Z(n303) );
  XNOR2_X1 U345 ( .A(G36GAT), .B(G29GAT), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U347 ( .A(KEYINPUT7), .B(n304), .Z(n352) );
  XOR2_X1 U348 ( .A(KEYINPUT66), .B(G8GAT), .Z(n306) );
  XNOR2_X1 U349 ( .A(G15GAT), .B(G113GAT), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U351 ( .A(n352), .B(n307), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n309), .B(n308), .ZN(n564) );
  XOR2_X1 U353 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n311) );
  XNOR2_X1 U354 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n325) );
  XNOR2_X1 U356 ( .A(G106GAT), .B(G78GAT), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n312), .B(G148GAT), .ZN(n391) );
  XOR2_X1 U358 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n314) );
  XNOR2_X1 U359 ( .A(G71GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n333) );
  XNOR2_X1 U361 ( .A(n391), .B(n333), .ZN(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT72), .B(KEYINPUT74), .Z(n316) );
  NAND2_X1 U363 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n317), .B(KEYINPUT73), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U367 ( .A(G176GAT), .B(G120GAT), .Z(n437) );
  XOR2_X1 U368 ( .A(G99GAT), .B(G85GAT), .Z(n350) );
  XNOR2_X1 U369 ( .A(n437), .B(n350), .ZN(n321) );
  XNOR2_X1 U370 ( .A(G204GAT), .B(G92GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n320), .B(G64GAT), .ZN(n380) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n570) );
  NOR2_X1 U373 ( .A1(n564), .A2(n543), .ZN(n328) );
  INV_X1 U374 ( .A(KEYINPUT112), .ZN(n326) );
  XOR2_X1 U375 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n330) );
  XNOR2_X1 U376 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n345) );
  XOR2_X1 U378 ( .A(G8GAT), .B(G211GAT), .Z(n384) );
  XOR2_X1 U379 ( .A(n384), .B(G78GAT), .Z(n332) );
  XOR2_X1 U380 ( .A(G15GAT), .B(G127GAT), .Z(n432) );
  XNOR2_X1 U381 ( .A(G183GAT), .B(n432), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U383 ( .A(G22GAT), .B(G155GAT), .Z(n395) );
  XOR2_X1 U384 ( .A(n333), .B(n395), .Z(n335) );
  NAND2_X1 U385 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U387 ( .A(n337), .B(n336), .Z(n343) );
  XOR2_X1 U388 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n339) );
  XNOR2_X1 U389 ( .A(KEYINPUT78), .B(KEYINPUT12), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U393 ( .A(n345), .B(n344), .ZN(n575) );
  XOR2_X1 U394 ( .A(n575), .B(KEYINPUT111), .Z(n553) );
  NAND2_X1 U395 ( .A1(n346), .A2(n553), .ZN(n347) );
  XNOR2_X1 U396 ( .A(n347), .B(KEYINPUT113), .ZN(n364) );
  XOR2_X1 U397 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n349) );
  XNOR2_X1 U398 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n351) );
  XOR2_X1 U400 ( .A(n351), .B(n350), .Z(n354) );
  XOR2_X1 U401 ( .A(G43GAT), .B(G134GAT), .Z(n435) );
  XNOR2_X1 U402 ( .A(n352), .B(n435), .ZN(n353) );
  XNOR2_X1 U403 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U404 ( .A(G50GAT), .B(G162GAT), .Z(n396) );
  XOR2_X1 U405 ( .A(G92GAT), .B(n396), .Z(n356) );
  NAND2_X1 U406 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U408 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U409 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n360) );
  XNOR2_X1 U410 ( .A(G190GAT), .B(KEYINPUT10), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U412 ( .A(G106GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U413 ( .A(n363), .B(n362), .ZN(n556) );
  NAND2_X1 U414 ( .A1(n364), .A2(n556), .ZN(n365) );
  XNOR2_X1 U415 ( .A(n365), .B(KEYINPUT47), .ZN(n370) );
  XNOR2_X1 U416 ( .A(KEYINPUT36), .B(n556), .ZN(n578) );
  NOR2_X1 U417 ( .A1(n578), .A2(n575), .ZN(n366) );
  XNOR2_X1 U418 ( .A(KEYINPUT45), .B(n366), .ZN(n367) );
  NAND2_X1 U419 ( .A1(n367), .A2(n564), .ZN(n368) );
  INV_X1 U420 ( .A(n570), .ZN(n451) );
  NOR2_X1 U421 ( .A1(n368), .A2(n451), .ZN(n369) );
  NOR2_X1 U422 ( .A1(n370), .A2(n369), .ZN(n372) );
  XOR2_X1 U423 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n374) );
  XNOR2_X1 U424 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U426 ( .A(n375), .B(KEYINPUT17), .Z(n377) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(G183GAT), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n377), .B(n376), .ZN(n444) );
  XOR2_X1 U429 ( .A(KEYINPUT21), .B(KEYINPUT88), .Z(n379) );
  XNOR2_X1 U430 ( .A(G197GAT), .B(G218GAT), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n392) );
  XNOR2_X1 U432 ( .A(n392), .B(n380), .ZN(n388) );
  XOR2_X1 U433 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n382) );
  XNOR2_X1 U434 ( .A(G36GAT), .B(G176GAT), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U436 ( .A(n384), .B(n383), .Z(n386) );
  NAND2_X1 U437 ( .A1(G226GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U439 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U440 ( .A(n444), .B(n389), .Z(n486) );
  INV_X1 U441 ( .A(n486), .ZN(n511) );
  NOR2_X1 U442 ( .A1(n523), .A2(n511), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n390), .B(KEYINPUT54), .ZN(n561) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n408) );
  XOR2_X1 U445 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n394) );
  XNOR2_X1 U446 ( .A(G211GAT), .B(G204GAT), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n400) );
  XOR2_X1 U448 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n398) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U451 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U452 ( .A1(G228GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U453 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U454 ( .A(n403), .B(KEYINPUT87), .Z(n406) );
  XNOR2_X1 U455 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U456 ( .A(n404), .B(KEYINPUT2), .ZN(n411) );
  XNOR2_X1 U457 ( .A(n411), .B(KEYINPUT89), .ZN(n405) );
  XNOR2_X1 U458 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U459 ( .A(n408), .B(n407), .ZN(n458) );
  XOR2_X1 U460 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n410) );
  XNOR2_X1 U461 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n409) );
  XNOR2_X1 U462 ( .A(n410), .B(n409), .ZN(n415) );
  XOR2_X1 U463 ( .A(G162GAT), .B(n411), .Z(n413) );
  XOR2_X1 U464 ( .A(G113GAT), .B(KEYINPUT0), .Z(n438) );
  XNOR2_X1 U465 ( .A(n438), .B(G134GAT), .ZN(n412) );
  XNOR2_X1 U466 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n428) );
  XOR2_X1 U468 ( .A(G85GAT), .B(G155GAT), .Z(n417) );
  XNOR2_X1 U469 ( .A(G29GAT), .B(G148GAT), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U471 ( .A(G57GAT), .B(G127GAT), .Z(n419) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G120GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U474 ( .A(n421), .B(n420), .Z(n426) );
  XOR2_X1 U475 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n423) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U478 ( .A(KEYINPUT92), .B(n424), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U480 ( .A(n428), .B(n427), .Z(n560) );
  AND2_X1 U481 ( .A1(n458), .A2(n560), .ZN(n429) );
  NAND2_X1 U482 ( .A1(n561), .A2(n429), .ZN(n431) );
  XOR2_X1 U483 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n447) );
  XOR2_X1 U485 ( .A(G71GAT), .B(n432), .Z(n434) );
  NAND2_X1 U486 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U488 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n446) );
  XOR2_X1 U491 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n442) );
  XNOR2_X1 U492 ( .A(G99GAT), .B(KEYINPUT83), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U494 ( .A(n444), .B(n443), .Z(n445) );
  XOR2_X1 U495 ( .A(n446), .B(n445), .Z(n514) );
  INV_X1 U496 ( .A(n514), .ZN(n527) );
  NAND2_X1 U497 ( .A1(n447), .A2(n527), .ZN(n555) );
  XNOR2_X1 U498 ( .A(n448), .B(G169GAT), .ZN(n450) );
  INV_X1 U499 ( .A(KEYINPUT120), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(G1348GAT) );
  NOR2_X1 U501 ( .A1(n564), .A2(n451), .ZN(n480) );
  XNOR2_X1 U502 ( .A(n514), .B(KEYINPUT85), .ZN(n454) );
  XNOR2_X1 U503 ( .A(n458), .B(KEYINPUT28), .ZN(n526) );
  INV_X1 U504 ( .A(n526), .ZN(n491) );
  INV_X1 U505 ( .A(n560), .ZN(n482) );
  XNOR2_X1 U506 ( .A(KEYINPUT27), .B(n486), .ZN(n456) );
  NAND2_X1 U507 ( .A1(n482), .A2(n456), .ZN(n524) );
  NOR2_X1 U508 ( .A1(n491), .A2(n524), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n452), .B(KEYINPUT95), .ZN(n453) );
  NOR2_X1 U510 ( .A1(n454), .A2(n453), .ZN(n465) );
  NOR2_X1 U511 ( .A1(n527), .A2(n458), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n455), .B(KEYINPUT26), .ZN(n562) );
  NAND2_X1 U513 ( .A1(n456), .A2(n562), .ZN(n461) );
  NAND2_X1 U514 ( .A1(n486), .A2(n527), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n458), .A2(n457), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT25), .B(n459), .Z(n460) );
  NAND2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U518 ( .A1(n462), .A2(n560), .ZN(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT96), .B(n463), .Z(n464) );
  NOR2_X1 U520 ( .A1(n465), .A2(n464), .ZN(n477) );
  INV_X1 U521 ( .A(n575), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n556), .A2(n466), .ZN(n467) );
  XNOR2_X1 U523 ( .A(KEYINPUT16), .B(n467), .ZN(n468) );
  NOR2_X1 U524 ( .A1(n477), .A2(n468), .ZN(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT97), .B(n469), .Z(n496) );
  NAND2_X1 U526 ( .A1(n480), .A2(n496), .ZN(n475) );
  NOR2_X1 U527 ( .A1(n560), .A2(n475), .ZN(n470) );
  XOR2_X1 U528 ( .A(G1GAT), .B(n470), .Z(n471) );
  XNOR2_X1 U529 ( .A(KEYINPUT34), .B(n471), .ZN(G1324GAT) );
  NOR2_X1 U530 ( .A1(n511), .A2(n475), .ZN(n472) );
  XOR2_X1 U531 ( .A(G8GAT), .B(n472), .Z(G1325GAT) );
  NOR2_X1 U532 ( .A1(n514), .A2(n475), .ZN(n474) );
  XNOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NOR2_X1 U535 ( .A1(n526), .A2(n475), .ZN(n476) );
  XOR2_X1 U536 ( .A(G22GAT), .B(n476), .Z(G1327GAT) );
  NOR2_X1 U537 ( .A1(n477), .A2(n578), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n575), .A2(n478), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n479), .B(KEYINPUT37), .ZN(n507) );
  NAND2_X1 U540 ( .A1(n480), .A2(n507), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT38), .B(n481), .Z(n492) );
  NAND2_X1 U542 ( .A1(n482), .A2(n492), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT98), .B(KEYINPUT39), .Z(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(n485), .ZN(G1328GAT) );
  XOR2_X1 U546 ( .A(G36GAT), .B(KEYINPUT99), .Z(n488) );
  NAND2_X1 U547 ( .A1(n486), .A2(n492), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1329GAT) );
  NAND2_X1 U549 ( .A1(n492), .A2(n527), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  NAND2_X1 U552 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT100), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  INV_X1 U555 ( .A(n564), .ZN(n495) );
  XOR2_X1 U556 ( .A(KEYINPUT101), .B(n543), .Z(n549) );
  NOR2_X1 U557 ( .A1(n495), .A2(n549), .ZN(n506) );
  NAND2_X1 U558 ( .A1(n496), .A2(n506), .ZN(n502) );
  NOR2_X1 U559 ( .A1(n560), .A2(n502), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U562 ( .A(G57GAT), .B(n499), .Z(G1332GAT) );
  NOR2_X1 U563 ( .A1(n511), .A2(n502), .ZN(n500) );
  XOR2_X1 U564 ( .A(G64GAT), .B(n500), .Z(G1333GAT) );
  NOR2_X1 U565 ( .A1(n514), .A2(n502), .ZN(n501) );
  XOR2_X1 U566 ( .A(G71GAT), .B(n501), .Z(G1334GAT) );
  NOR2_X1 U567 ( .A1(n526), .A2(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT43), .B(KEYINPUT103), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U570 ( .A(G78GAT), .B(n505), .Z(G1335GAT) );
  NAND2_X1 U571 ( .A1(n507), .A2(n506), .ZN(n520) );
  NOR2_X1 U572 ( .A1(n560), .A2(n520), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NOR2_X1 U576 ( .A1(n511), .A2(n520), .ZN(n512) );
  XOR2_X1 U577 ( .A(KEYINPUT106), .B(n512), .Z(n513) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(n513), .ZN(G1337GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n520), .ZN(n516) );
  XNOR2_X1 U580 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n517), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n519) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n522) );
  NOR2_X1 U586 ( .A1(n526), .A2(n520), .ZN(n521) );
  XOR2_X1 U587 ( .A(n522), .B(n521), .Z(G1339GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U589 ( .A(n525), .B(KEYINPUT115), .Z(n538) );
  AND2_X1 U590 ( .A1(n526), .A2(n538), .ZN(n528) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n535) );
  NOR2_X1 U592 ( .A1(n564), .A2(n535), .ZN(n529) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n529), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n549), .A2(n535), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U597 ( .A1(n553), .A2(n535), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  NOR2_X1 U601 ( .A1(n556), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n538), .A2(n562), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n564), .A2(n547), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n542) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n543), .A2(n547), .ZN(n544) );
  XOR2_X1 U612 ( .A(n545), .B(n544), .Z(G1345GAT) );
  NOR2_X1 U613 ( .A1(n575), .A2(n547), .ZN(n546) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n546), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n556), .A2(n547), .ZN(n548) );
  XOR2_X1 U616 ( .A(G162GAT), .B(n548), .Z(G1347GAT) );
  NOR2_X1 U617 ( .A1(n555), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(n552), .ZN(G1349GAT) );
  NOR2_X1 U621 ( .A1(n553), .A2(n555), .ZN(n554) );
  XOR2_X1 U622 ( .A(G183GAT), .B(n554), .Z(G1350GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n558) );
  INV_X1 U624 ( .A(KEYINPUT58), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G190GAT), .ZN(G1351GAT) );
  AND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n577) );
  NOR2_X1 U629 ( .A1(n564), .A2(n577), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n566) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT121), .B(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n577), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n577), .ZN(n576) );
  XOR2_X1 U641 ( .A(G211GAT), .B(n576), .Z(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n583) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(KEYINPUT125), .B(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1355GAT) );
endmodule

