

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738;

  XOR2_X1 U375 ( .A(KEYINPUT4), .B(KEYINPUT71), .Z(n427) );
  XNOR2_X1 U376 ( .A(G146), .B(G125), .ZN(n458) );
  XNOR2_X1 U377 ( .A(n393), .B(n392), .ZN(n690) );
  INV_X1 U378 ( .A(G953), .ZN(n725) );
  NOR2_X1 U379 ( .A1(n690), .A2(n584), .ZN(n391) );
  NOR2_X2 U380 ( .A1(n671), .A2(n670), .ZN(n582) );
  NOR2_X2 U381 ( .A1(n507), .A2(n508), .ZN(n539) );
  NOR2_X1 U382 ( .A1(n616), .A2(n709), .ZN(n617) );
  XNOR2_X1 U383 ( .A(n401), .B(n400), .ZN(n735) );
  XNOR2_X1 U384 ( .A(n377), .B(n376), .ZN(n737) );
  OR2_X1 U385 ( .A1(n555), .A2(n645), .ZN(n377) );
  XNOR2_X1 U386 ( .A(n570), .B(n569), .ZN(n594) );
  XNOR2_X1 U387 ( .A(n387), .B(G134), .ZN(n486) );
  XNOR2_X1 U388 ( .A(n435), .B(n434), .ZN(n436) );
  AND2_X1 U389 ( .A1(n527), .A2(n528), .ZN(n551) );
  NOR2_X1 U390 ( .A1(n737), .A2(n738), .ZN(n543) );
  OR2_X1 U391 ( .A1(n625), .A2(G902), .ZN(n394) );
  OR2_X1 U392 ( .A1(n707), .A2(G902), .ZN(n374) );
  XNOR2_X1 U393 ( .A(n422), .B(n421), .ZN(n441) );
  XNOR2_X1 U394 ( .A(n420), .B(KEYINPUT3), .ZN(n421) );
  XNOR2_X1 U395 ( .A(G113), .B(KEYINPUT75), .ZN(n419) );
  NAND2_X1 U396 ( .A1(n386), .A2(n553), .ZN(n384) );
  INV_X1 U397 ( .A(n653), .ZN(n363) );
  AND2_X1 U398 ( .A1(n551), .A2(n360), .ZN(n379) );
  NAND2_X1 U399 ( .A1(KEYINPUT44), .A2(n603), .ZN(n389) );
  XOR2_X1 U400 ( .A(KEYINPUT107), .B(KEYINPUT7), .Z(n489) );
  XNOR2_X1 U401 ( .A(G122), .B(KEYINPUT106), .ZN(n488) );
  XOR2_X1 U402 ( .A(G131), .B(G140), .Z(n472) );
  XNOR2_X1 U403 ( .A(n531), .B(n530), .ZN(n665) );
  XNOR2_X1 U404 ( .A(n676), .B(n444), .ZN(n556) );
  XNOR2_X1 U405 ( .A(KEYINPUT108), .B(KEYINPUT6), .ZN(n444) );
  XNOR2_X1 U406 ( .A(G137), .B(KEYINPUT24), .ZN(n459) );
  INV_X1 U407 ( .A(G119), .ZN(n407) );
  XNOR2_X1 U408 ( .A(G143), .B(G122), .ZN(n473) );
  XNOR2_X1 U409 ( .A(n423), .B(n366), .ZN(n431) );
  INV_X1 U410 ( .A(G107), .ZN(n366) );
  XNOR2_X1 U411 ( .A(n395), .B(n717), .ZN(n618) );
  XNOR2_X1 U412 ( .A(n397), .B(n396), .ZN(n395) );
  XNOR2_X1 U413 ( .A(n540), .B(n378), .ZN(n555) );
  INV_X1 U414 ( .A(KEYINPUT39), .ZN(n378) );
  AND2_X1 U415 ( .A1(n365), .A2(n404), .ZN(n536) );
  XNOR2_X1 U416 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n569) );
  NAND2_X1 U417 ( .A1(n568), .A2(n567), .ZN(n570) );
  AND2_X1 U418 ( .A1(n659), .A2(n566), .ZN(n567) );
  NOR2_X2 U419 ( .A1(n594), .A2(n583), .ZN(n592) );
  INV_X1 U420 ( .A(KEYINPUT84), .ZN(n511) );
  INV_X1 U421 ( .A(n506), .ZN(n402) );
  XNOR2_X1 U422 ( .A(G116), .B(G119), .ZN(n420) );
  XOR2_X1 U423 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n416) );
  XNOR2_X1 U424 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n529) );
  NOR2_X1 U425 ( .A1(G237), .A2(G902), .ZN(n425) );
  XNOR2_X1 U426 ( .A(n443), .B(n442), .ZN(n625) );
  NOR2_X1 U427 ( .A1(n385), .A2(n363), .ZN(n362) );
  NAND2_X1 U428 ( .A1(n382), .A2(n384), .ZN(n381) );
  NOR2_X1 U429 ( .A1(n602), .A2(n411), .ZN(n606) );
  XNOR2_X1 U430 ( .A(G116), .B(G107), .ZN(n487) );
  XOR2_X1 U431 ( .A(KEYINPUT15), .B(G902), .Z(n608) );
  INV_X1 U432 ( .A(KEYINPUT33), .ZN(n392) );
  BUF_X1 U433 ( .A(n676), .Z(n364) );
  XNOR2_X1 U434 ( .A(n441), .B(n398), .ZN(n717) );
  XNOR2_X1 U435 ( .A(n431), .B(n424), .ZN(n398) );
  XNOR2_X1 U436 ( .A(n375), .B(n405), .ZN(n707) );
  XNOR2_X1 U437 ( .A(n471), .B(n406), .ZN(n405) );
  XNOR2_X1 U438 ( .A(n459), .B(n407), .ZN(n406) );
  XNOR2_X1 U439 ( .A(G113), .B(G104), .ZN(n480) );
  NOR2_X1 U440 ( .A1(G952), .A2(n725), .ZN(n709) );
  INV_X1 U441 ( .A(KEYINPUT40), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n593), .B(KEYINPUT80), .ZN(n400) );
  NAND2_X1 U443 ( .A1(n592), .A2(n591), .ZN(n401) );
  INV_X1 U444 ( .A(KEYINPUT111), .ZN(n408) );
  XOR2_X1 U445 ( .A(KEYINPUT81), .B(n519), .Z(n643) );
  NAND2_X1 U446 ( .A1(n372), .A2(n404), .ZN(n574) );
  NAND2_X1 U447 ( .A1(n402), .A2(KEYINPUT79), .ZN(n352) );
  AND2_X1 U448 ( .A1(n549), .A2(n652), .ZN(n353) );
  XNOR2_X1 U449 ( .A(KEYINPUT109), .B(n502), .ZN(n354) );
  AND2_X1 U450 ( .A1(n539), .A2(n513), .ZN(n355) );
  INV_X1 U451 ( .A(n518), .ZN(n404) );
  AND2_X1 U452 ( .A1(n453), .A2(G210), .ZN(n356) );
  AND2_X1 U453 ( .A1(n383), .A2(n381), .ZN(n357) );
  AND2_X1 U454 ( .A1(n353), .A2(n386), .ZN(n358) );
  AND2_X1 U455 ( .A1(n604), .A2(n389), .ZN(n359) );
  AND2_X1 U456 ( .A1(n353), .A2(n553), .ZN(n360) );
  INV_X1 U457 ( .A(KEYINPUT79), .ZN(n403) );
  XOR2_X1 U458 ( .A(n612), .B(n611), .Z(n361) );
  NOR2_X2 U459 ( .A1(n700), .A2(n709), .ZN(n701) );
  NOR2_X2 U460 ( .A1(n623), .A2(n709), .ZN(n624) );
  NOR2_X2 U461 ( .A1(n628), .A2(n709), .ZN(n630) );
  NOR2_X2 U462 ( .A1(n724), .A2(n714), .ZN(n609) );
  NOR2_X2 U463 ( .A1(n609), .A2(KEYINPUT2), .ZN(n656) );
  XNOR2_X1 U464 ( .A(n417), .B(n414), .ZN(n397) );
  NAND2_X1 U465 ( .A1(n673), .A2(n566), .ZN(n505) );
  XNOR2_X2 U466 ( .A(n374), .B(n470), .ZN(n673) );
  XNOR2_X1 U467 ( .A(n466), .B(n469), .ZN(n375) );
  NAND2_X1 U468 ( .A1(n357), .A2(n362), .ZN(n724) );
  NOR2_X2 U469 ( .A1(G902), .A2(n613), .ZN(n437) );
  XNOR2_X2 U470 ( .A(n518), .B(KEYINPUT1), .ZN(n670) );
  XNOR2_X2 U471 ( .A(n437), .B(n436), .ZN(n518) );
  NAND2_X2 U472 ( .A1(n609), .A2(KEYINPUT2), .ZN(n657) );
  NAND2_X1 U473 ( .A1(n380), .A2(n379), .ZN(n383) );
  XNOR2_X2 U474 ( .A(n722), .B(G146), .ZN(n443) );
  XNOR2_X2 U475 ( .A(n486), .B(n428), .ZN(n722) );
  XNOR2_X1 U476 ( .A(n517), .B(KEYINPUT28), .ZN(n365) );
  NAND2_X1 U477 ( .A1(n582), .A2(n583), .ZN(n393) );
  NOR2_X2 U478 ( .A1(n735), .A2(n639), .ZN(n604) );
  AND2_X1 U479 ( .A1(n368), .A2(n367), .ZN(n370) );
  NAND2_X1 U480 ( .A1(n671), .A2(n403), .ZN(n367) );
  XNOR2_X2 U481 ( .A(n505), .B(n504), .ZN(n671) );
  NAND2_X1 U482 ( .A1(n373), .A2(n403), .ZN(n368) );
  NAND2_X1 U483 ( .A1(n370), .A2(n369), .ZN(n507) );
  NAND2_X1 U484 ( .A1(n371), .A2(n372), .ZN(n369) );
  NOR2_X1 U485 ( .A1(n518), .A2(n352), .ZN(n371) );
  INV_X1 U486 ( .A(n671), .ZN(n372) );
  NAND2_X1 U487 ( .A1(n404), .A2(n402), .ZN(n373) );
  INV_X1 U488 ( .A(n550), .ZN(n380) );
  NAND2_X1 U489 ( .A1(n551), .A2(n358), .ZN(n382) );
  AND2_X1 U490 ( .A1(n550), .A2(n554), .ZN(n385) );
  INV_X1 U491 ( .A(n654), .ZN(n386) );
  XNOR2_X1 U492 ( .A(n387), .B(n418), .ZN(n396) );
  XNOR2_X2 U493 ( .A(n412), .B(G143), .ZN(n387) );
  NAND2_X1 U494 ( .A1(n388), .A2(n603), .ZN(n390) );
  XNOR2_X1 U495 ( .A(n736), .B(KEYINPUT68), .ZN(n388) );
  NAND2_X1 U496 ( .A1(n390), .A2(n359), .ZN(n605) );
  XNOR2_X1 U497 ( .A(n391), .B(n585), .ZN(n586) );
  XNOR2_X2 U498 ( .A(n394), .B(G472), .ZN(n676) );
  AND2_X2 U499 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X2 U500 ( .A(G128), .B(KEYINPUT82), .ZN(n412) );
  NAND2_X1 U501 ( .A1(n562), .A2(n563), .ZN(n564) );
  XNOR2_X2 U502 ( .A(n399), .B(n514), .ZN(n562) );
  NAND2_X1 U503 ( .A1(n513), .A2(n660), .ZN(n399) );
  XNOR2_X2 U504 ( .A(n426), .B(n356), .ZN(n513) );
  XNOR2_X2 U505 ( .A(n409), .B(n408), .ZN(n734) );
  NAND2_X1 U506 ( .A1(n410), .A2(n354), .ZN(n409) );
  XNOR2_X1 U507 ( .A(n355), .B(KEYINPUT110), .ZN(n410) );
  XNOR2_X1 U508 ( .A(n512), .B(n511), .ZN(n528) );
  XNOR2_X1 U509 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X2 U510 ( .A(n607), .B(KEYINPUT45), .ZN(n714) );
  XNOR2_X1 U511 ( .A(n513), .B(n529), .ZN(n661) );
  XNOR2_X2 U512 ( .A(n564), .B(KEYINPUT0), .ZN(n584) );
  AND2_X1 U513 ( .A1(n601), .A2(n600), .ZN(n411) );
  XNOR2_X1 U514 ( .A(KEYINPUT17), .B(KEYINPUT92), .ZN(n413) );
  XNOR2_X1 U515 ( .A(n541), .B(KEYINPUT46), .ZN(n542) );
  INV_X1 U516 ( .A(KEYINPUT88), .ZN(n552) );
  XNOR2_X1 U517 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U518 ( .A(n552), .B(KEYINPUT48), .ZN(n553) );
  INV_X1 U519 ( .A(n565), .ZN(n566) );
  INV_X1 U520 ( .A(n553), .ZN(n554) );
  INV_X1 U521 ( .A(KEYINPUT112), .ZN(n530) );
  INV_X1 U522 ( .A(G469), .ZN(n434) );
  XNOR2_X1 U523 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U524 ( .A(n441), .B(n440), .ZN(n442) );
  INV_X1 U525 ( .A(KEYINPUT32), .ZN(n593) );
  INV_X1 U526 ( .A(KEYINPUT63), .ZN(n629) );
  XNOR2_X1 U527 ( .A(n427), .B(n413), .ZN(n414) );
  INV_X1 U528 ( .A(n458), .ZN(n415) );
  AND2_X1 U529 ( .A1(G224), .A2(n725), .ZN(n418) );
  XOR2_X1 U530 ( .A(G122), .B(KEYINPUT16), .Z(n424) );
  XNOR2_X1 U531 ( .A(n419), .B(G101), .ZN(n422) );
  XNOR2_X1 U532 ( .A(G104), .B(G110), .ZN(n423) );
  INV_X1 U533 ( .A(n608), .ZN(n445) );
  NAND2_X1 U534 ( .A1(n618), .A2(n445), .ZN(n426) );
  XOR2_X1 U535 ( .A(KEYINPUT78), .B(n425), .Z(n453) );
  INV_X1 U536 ( .A(n513), .ZN(n546) );
  XNOR2_X1 U537 ( .A(G137), .B(n427), .ZN(n428) );
  XOR2_X1 U538 ( .A(G101), .B(n472), .Z(n430) );
  NAND2_X1 U539 ( .A1(G227), .A2(n725), .ZN(n429) );
  XNOR2_X1 U540 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X2 U541 ( .A(n443), .B(n433), .ZN(n613) );
  XNOR2_X1 U542 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n435) );
  INV_X1 U543 ( .A(n670), .ZN(n595) );
  XOR2_X1 U544 ( .A(G131), .B(KEYINPUT5), .Z(n439) );
  NOR2_X1 U545 ( .A1(G953), .A2(G237), .ZN(n476) );
  NAND2_X1 U546 ( .A1(n476), .A2(G210), .ZN(n438) );
  XNOR2_X1 U547 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U548 ( .A1(G234), .A2(n445), .ZN(n446) );
  XNOR2_X1 U549 ( .A(KEYINPUT20), .B(n446), .ZN(n455) );
  NAND2_X1 U550 ( .A1(G221), .A2(n455), .ZN(n447) );
  XNOR2_X1 U551 ( .A(n447), .B(KEYINPUT21), .ZN(n565) );
  XOR2_X1 U552 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n449) );
  NAND2_X1 U553 ( .A1(G234), .A2(G237), .ZN(n448) );
  XNOR2_X1 U554 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U555 ( .A1(G952), .A2(n450), .ZN(n688) );
  NOR2_X1 U556 ( .A1(G953), .A2(n688), .ZN(n560) );
  NAND2_X1 U557 ( .A1(G902), .A2(n450), .ZN(n558) );
  OR2_X1 U558 ( .A1(n725), .A2(n558), .ZN(n451) );
  NOR2_X1 U559 ( .A1(G900), .A2(n451), .ZN(n452) );
  NOR2_X1 U560 ( .A1(n560), .A2(n452), .ZN(n506) );
  NOR2_X1 U561 ( .A1(n565), .A2(n506), .ZN(n515) );
  NAND2_X1 U562 ( .A1(n453), .A2(G214), .ZN(n660) );
  NAND2_X1 U563 ( .A1(n515), .A2(n660), .ZN(n454) );
  NOR2_X1 U564 ( .A1(n556), .A2(n454), .ZN(n499) );
  XOR2_X1 U565 ( .A(KEYINPUT25), .B(KEYINPUT100), .Z(n457) );
  NAND2_X1 U566 ( .A1(n455), .A2(G217), .ZN(n456) );
  XNOR2_X1 U567 ( .A(n457), .B(n456), .ZN(n470) );
  XNOR2_X1 U568 ( .A(KEYINPUT10), .B(n458), .ZN(n471) );
  XOR2_X1 U569 ( .A(KEYINPUT86), .B(G140), .Z(n461) );
  XNOR2_X1 U570 ( .A(G128), .B(G110), .ZN(n460) );
  XNOR2_X1 U571 ( .A(n461), .B(n460), .ZN(n465) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(KEYINPUT98), .Z(n463) );
  XNOR2_X1 U573 ( .A(KEYINPUT97), .B(KEYINPUT99), .ZN(n462) );
  XNOR2_X1 U574 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U575 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U576 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n468) );
  NAND2_X1 U577 ( .A1(G234), .A2(n725), .ZN(n467) );
  XNOR2_X1 U578 ( .A(n468), .B(n467), .ZN(n492) );
  AND2_X1 U579 ( .A1(G221), .A2(n492), .ZN(n469) );
  XNOR2_X1 U580 ( .A(KEYINPUT13), .B(G475), .ZN(n485) );
  XOR2_X1 U581 ( .A(n472), .B(n471), .Z(n723) );
  XOR2_X1 U582 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n474) );
  XNOR2_X1 U583 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U584 ( .A(n723), .B(n475), .ZN(n483) );
  XOR2_X1 U585 ( .A(KEYINPUT105), .B(KEYINPUT11), .Z(n478) );
  NAND2_X1 U586 ( .A1(G214), .A2(n476), .ZN(n477) );
  XNOR2_X1 U587 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U588 ( .A(n479), .B(KEYINPUT12), .Z(n481) );
  XNOR2_X1 U589 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n483), .B(n482), .ZN(n697) );
  NOR2_X1 U591 ( .A1(G902), .A2(n697), .ZN(n484) );
  XNOR2_X1 U592 ( .A(n485), .B(n484), .ZN(n533) );
  INV_X1 U593 ( .A(n486), .ZN(n496) );
  XNOR2_X1 U594 ( .A(n487), .B(KEYINPUT9), .ZN(n491) );
  XNOR2_X1 U595 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U596 ( .A(n491), .B(n490), .Z(n494) );
  NAND2_X1 U597 ( .A1(n492), .A2(G217), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U599 ( .A(n496), .B(n495), .ZN(n703) );
  NOR2_X1 U600 ( .A1(G902), .A2(n703), .ZN(n497) );
  XNOR2_X1 U601 ( .A(G478), .B(n497), .ZN(n509) );
  NAND2_X1 U602 ( .A1(n533), .A2(n509), .ZN(n645) );
  NOR2_X1 U603 ( .A1(n673), .A2(n645), .ZN(n498) );
  NAND2_X1 U604 ( .A1(n499), .A2(n498), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n595), .A2(n545), .ZN(n500) );
  XNOR2_X1 U606 ( .A(n500), .B(KEYINPUT43), .ZN(n501) );
  NOR2_X1 U607 ( .A1(n513), .A2(n501), .ZN(n654) );
  INV_X1 U608 ( .A(n509), .ZN(n532) );
  NAND2_X1 U609 ( .A1(n533), .A2(n532), .ZN(n502) );
  NAND2_X1 U610 ( .A1(n676), .A2(n660), .ZN(n503) );
  XNOR2_X1 U611 ( .A(KEYINPUT30), .B(n503), .ZN(n508) );
  INV_X1 U612 ( .A(KEYINPUT69), .ZN(n504) );
  OR2_X1 U613 ( .A1(n533), .A2(n509), .ZN(n647) );
  NAND2_X1 U614 ( .A1(n645), .A2(n647), .ZN(n664) );
  INV_X1 U615 ( .A(n664), .ZN(n521) );
  NAND2_X1 U616 ( .A1(KEYINPUT47), .A2(n521), .ZN(n510) );
  NAND2_X1 U617 ( .A1(n734), .A2(n510), .ZN(n512) );
  XOR2_X1 U618 ( .A(KEYINPUT19), .B(KEYINPUT67), .Z(n514) );
  INV_X1 U619 ( .A(n676), .ZN(n576) );
  INV_X1 U620 ( .A(n673), .ZN(n596) );
  NAND2_X1 U621 ( .A1(n515), .A2(n596), .ZN(n516) );
  NOR2_X1 U622 ( .A1(n576), .A2(n516), .ZN(n517) );
  NAND2_X1 U623 ( .A1(n562), .A2(n536), .ZN(n519) );
  XNOR2_X1 U624 ( .A(KEYINPUT47), .B(KEYINPUT70), .ZN(n520) );
  NOR2_X1 U625 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U626 ( .A1(KEYINPUT85), .A2(n522), .ZN(n523) );
  NOR2_X1 U627 ( .A1(n643), .A2(n523), .ZN(n526) );
  NAND2_X1 U628 ( .A1(KEYINPUT47), .A2(n643), .ZN(n524) );
  NOR2_X1 U629 ( .A1(KEYINPUT85), .A2(n524), .ZN(n525) );
  NOR2_X1 U630 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U631 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n535) );
  NAND2_X1 U632 ( .A1(n661), .A2(n660), .ZN(n531) );
  NOR2_X1 U633 ( .A1(n533), .A2(n532), .ZN(n659) );
  NAND2_X1 U634 ( .A1(n665), .A2(n659), .ZN(n534) );
  XNOR2_X1 U635 ( .A(n535), .B(n534), .ZN(n689) );
  INV_X1 U636 ( .A(n536), .ZN(n537) );
  NOR2_X1 U637 ( .A1(n689), .A2(n537), .ZN(n538) );
  XNOR2_X1 U638 ( .A(KEYINPUT42), .B(n538), .ZN(n738) );
  NAND2_X1 U639 ( .A1(n661), .A2(n539), .ZN(n540) );
  XNOR2_X1 U640 ( .A(KEYINPUT89), .B(KEYINPUT64), .ZN(n541) );
  XNOR2_X1 U641 ( .A(n543), .B(n542), .ZN(n550) );
  INV_X1 U642 ( .A(KEYINPUT47), .ZN(n544) );
  NAND2_X1 U643 ( .A1(KEYINPUT85), .A2(n544), .ZN(n549) );
  NOR2_X1 U644 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U645 ( .A(KEYINPUT36), .B(n547), .ZN(n548) );
  NAND2_X1 U646 ( .A1(n548), .A2(n595), .ZN(n652) );
  OR2_X1 U647 ( .A1(n555), .A2(n647), .ZN(n653) );
  INV_X1 U648 ( .A(n556), .ZN(n583) );
  XOR2_X1 U649 ( .A(G898), .B(KEYINPUT94), .Z(n713) );
  NAND2_X1 U650 ( .A1(n713), .A2(G953), .ZN(n557) );
  XOR2_X1 U651 ( .A(KEYINPUT95), .B(n557), .Z(n718) );
  NOR2_X1 U652 ( .A1(n558), .A2(n718), .ZN(n559) );
  NOR2_X1 U653 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U654 ( .A(KEYINPUT96), .B(n561), .Z(n563) );
  INV_X1 U655 ( .A(n584), .ZN(n568) );
  NAND2_X1 U656 ( .A1(n592), .A2(n670), .ZN(n571) );
  NOR2_X1 U657 ( .A1(n596), .A2(n571), .ZN(n631) );
  NAND2_X1 U658 ( .A1(n364), .A2(n582), .ZN(n679) );
  NOR2_X1 U659 ( .A1(n584), .A2(n679), .ZN(n573) );
  XNOR2_X1 U660 ( .A(KEYINPUT31), .B(KEYINPUT102), .ZN(n572) );
  XNOR2_X1 U661 ( .A(n573), .B(n572), .ZN(n648) );
  OR2_X1 U662 ( .A1(n584), .A2(n574), .ZN(n575) );
  XNOR2_X1 U663 ( .A(n575), .B(KEYINPUT101), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n634) );
  NAND2_X1 U665 ( .A1(n648), .A2(n634), .ZN(n578) );
  NAND2_X1 U666 ( .A1(n578), .A2(n664), .ZN(n580) );
  INV_X1 U667 ( .A(KEYINPUT44), .ZN(n599) );
  NAND2_X1 U668 ( .A1(KEYINPUT65), .A2(n599), .ZN(n579) );
  NAND2_X1 U669 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U670 ( .A1(n631), .A2(n581), .ZN(n590) );
  XNOR2_X1 U671 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n585) );
  NAND2_X1 U672 ( .A1(n586), .A2(n354), .ZN(n588) );
  XOR2_X1 U673 ( .A(KEYINPUT35), .B(KEYINPUT87), .Z(n587) );
  XNOR2_X2 U674 ( .A(n588), .B(n587), .ZN(n736) );
  NAND2_X1 U675 ( .A1(n736), .A2(KEYINPUT44), .ZN(n589) );
  NAND2_X1 U676 ( .A1(n590), .A2(n589), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n670), .A2(n673), .ZN(n591) );
  NOR2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U680 ( .A1(n364), .A2(n598), .ZN(n639) );
  NAND2_X1 U681 ( .A1(KEYINPUT68), .A2(n604), .ZN(n601) );
  NOR2_X1 U682 ( .A1(KEYINPUT65), .A2(n599), .ZN(n600) );
  INV_X1 U683 ( .A(KEYINPUT65), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n657), .A2(n608), .ZN(n610) );
  NOR2_X4 U685 ( .A1(n610), .A2(n656), .ZN(n705) );
  NAND2_X1 U686 ( .A1(n705), .A2(G469), .ZN(n615) );
  XOR2_X1 U687 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n612) );
  XNOR2_X1 U688 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n611) );
  XNOR2_X1 U689 ( .A(n613), .B(n361), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n617), .B(KEYINPUT124), .ZN(G54) );
  XNOR2_X1 U691 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n618), .B(KEYINPUT90), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n705), .A2(G210), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n624), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U697 ( .A(n625), .B(KEYINPUT62), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n705), .A2(G472), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(G57) );
  XOR2_X1 U701 ( .A(G101), .B(n631), .Z(G3) );
  NOR2_X1 U702 ( .A1(n645), .A2(n634), .ZN(n632) );
  XOR2_X1 U703 ( .A(KEYINPUT114), .B(n632), .Z(n633) );
  XNOR2_X1 U704 ( .A(G104), .B(n633), .ZN(G6) );
  NOR2_X1 U705 ( .A1(n634), .A2(n647), .ZN(n638) );
  XOR2_X1 U706 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n636) );
  XNOR2_X1 U707 ( .A(G107), .B(KEYINPUT115), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(G9) );
  XOR2_X1 U710 ( .A(G110), .B(n639), .Z(G12) );
  NOR2_X1 U711 ( .A1(n647), .A2(n643), .ZN(n641) );
  XNOR2_X1 U712 ( .A(KEYINPUT29), .B(KEYINPUT116), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U714 ( .A(G128), .B(n642), .ZN(G30) );
  NOR2_X1 U715 ( .A1(n645), .A2(n643), .ZN(n644) );
  XOR2_X1 U716 ( .A(G146), .B(n644), .Z(G48) );
  NOR2_X1 U717 ( .A1(n648), .A2(n645), .ZN(n646) );
  XOR2_X1 U718 ( .A(G113), .B(n646), .Z(G15) );
  NOR2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U720 ( .A(KEYINPUT118), .B(n649), .Z(n650) );
  XNOR2_X1 U721 ( .A(G116), .B(n650), .ZN(G18) );
  XOR2_X1 U722 ( .A(G125), .B(KEYINPUT37), .Z(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(G27) );
  XNOR2_X1 U724 ( .A(G134), .B(n653), .ZN(G36) );
  XNOR2_X1 U725 ( .A(G140), .B(n654), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n655), .B(KEYINPUT119), .ZN(G42) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT83), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n694) );
  INV_X1 U729 ( .A(n659), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U733 ( .A(KEYINPUT120), .B(n666), .Z(n667) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n669), .A2(n690), .ZN(n684) );
  NAND2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(KEYINPUT50), .ZN(n678) );
  NOR2_X1 U738 ( .A1(n566), .A2(n673), .ZN(n674) );
  XOR2_X1 U739 ( .A(KEYINPUT49), .B(n674), .Z(n675) );
  NOR2_X1 U740 ( .A1(n364), .A2(n675), .ZN(n677) );
  NAND2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n680) );
  NAND2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U743 ( .A(KEYINPUT51), .B(n681), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n682), .A2(n689), .ZN(n683) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U746 ( .A(n685), .B(KEYINPUT52), .Z(n686) );
  XNOR2_X1 U747 ( .A(KEYINPUT121), .B(n686), .ZN(n687) );
  NOR2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n692) );
  NOR2_X1 U749 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U750 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U751 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U752 ( .A1(n695), .A2(G953), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n696), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U754 ( .A(n697), .B(KEYINPUT59), .Z(n699) );
  NAND2_X1 U755 ( .A1(n705), .A2(G475), .ZN(n698) );
  XNOR2_X1 U756 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n701), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U758 ( .A1(G478), .A2(n705), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n709), .A2(n704), .ZN(G63) );
  NAND2_X1 U761 ( .A1(G217), .A2(n705), .ZN(n706) );
  XNOR2_X1 U762 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n709), .A2(n708), .ZN(G66) );
  NAND2_X1 U764 ( .A1(G224), .A2(G953), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n710), .B(KEYINPUT125), .ZN(n711) );
  XNOR2_X1 U766 ( .A(n711), .B(KEYINPUT61), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U768 ( .A1(G953), .A2(n714), .ZN(n715) );
  NOR2_X1 U769 ( .A1(n716), .A2(n715), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U771 ( .A(n719), .B(KEYINPUT126), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(G69) );
  XOR2_X1 U773 ( .A(n722), .B(n723), .Z(n727) );
  XNOR2_X1 U774 ( .A(n727), .B(n724), .ZN(n726) );
  NAND2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n732) );
  XNOR2_X1 U776 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n728), .A2(G900), .ZN(n729) );
  XOR2_X1 U778 ( .A(KEYINPUT127), .B(n729), .Z(n730) );
  NAND2_X1 U779 ( .A1(G953), .A2(n730), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n732), .A2(n731), .ZN(G72) );
  XOR2_X1 U781 ( .A(G143), .B(KEYINPUT117), .Z(n733) );
  XNOR2_X1 U782 ( .A(n734), .B(n733), .ZN(G45) );
  XOR2_X1 U783 ( .A(n735), .B(G119), .Z(G21) );
  XOR2_X1 U784 ( .A(n736), .B(G122), .Z(G24) );
  XOR2_X1 U785 ( .A(G131), .B(n737), .Z(G33) );
  XOR2_X1 U786 ( .A(G137), .B(n738), .Z(G39) );
endmodule

