//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1' ..
//Module:
 module locked_c3540( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  , KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0);
input KEYINPUT0;
input KEYINPUT1;
input KEYINPUT2;
input KEYINPUT3;
input KEYINPUT4;
input KEYINPUT5;
input KEYINPUT6;
input KEYINPUT7;
input KEYINPUT8;
input KEYINPUT9;
input KEYINPUT10;
input KEYINPUT11;
input KEYINPUT12;
input KEYINPUT13;
input KEYINPUT14;
input KEYINPUT15;
input KEYINPUT16;
input KEYINPUT17;
input KEYINPUT18;
input KEYINPUT19;
input KEYINPUT20;
input KEYINPUT21;
input KEYINPUT22;
input KEYINPUT23;
input KEYINPUT24;
input KEYINPUT25;
input KEYINPUT26;
input KEYINPUT27;
input KEYINPUT28;
input KEYINPUT29;
input KEYINPUT30;
input KEYINPUT31;
input KEYINPUT32;
input KEYINPUT33;
input KEYINPUT34;
input KEYINPUT35;
input KEYINPUT36;
input KEYINPUT37;
input KEYINPUT38;
input KEYINPUT39;
input KEYINPUT40;
input KEYINPUT41;
input KEYINPUT42;
input KEYINPUT43;
input KEYINPUT44;
input KEYINPUT45;
input KEYINPUT46;
input KEYINPUT47;
input KEYINPUT48;
input KEYINPUT49;
input KEYINPUT50;
input KEYINPUT51;
input KEYINPUT52;
input KEYINPUT53;
input KEYINPUT54;
input KEYINPUT55;
input KEYINPUT56;
input KEYINPUT57;
input KEYINPUT58;
input KEYINPUT59;
input KEYINPUT60;
input KEYINPUT61;
input KEYINPUT62;
input KEYINPUT63;
//Header:
   input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n73_, new_n74_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_,
    new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_,
    new_n96_, new_n97_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n106_, new_n107_, new_n108_, new_n109_,
    new_n110_, new_n111_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_;
wire RLL_wire_A_0;
wire RLL_wire_A_1;
wire RLL_wire_A_2;
wire RLL_wire_A_3;
wire RLL_wire_A_4;
wire RLL_wire_A_5;
wire RLL_wire_A_6;
wire RLL_wire_A_7;
wire RLL_wire_A_8;
wire RLL_wire_A_9;
wire RLL_wire_A_10;
wire RLL_wire_A_11;
wire RLL_wire_A_12;
wire RLL_wire_A_13;
wire RLL_wire_A_14;
wire RLL_wire_A_15;
wire RLL_wire_A_16;
wire RLL_wire_A_17;
wire RLL_wire_A_18;
wire RLL_wire_A_19;
wire RLL_wire_A_20;
wire RLL_wire_A_21;
wire RLL_wire_A_22;
wire RLL_wire_A_23;
wire RLL_wire_A_24;
wire RLL_wire_A_25;
wire RLL_wire_A_26;
wire RLL_wire_A_27;
wire RLL_wire_A_28;
wire RLL_wire_A_29;
wire RLL_wire_A_30;
wire RLL_wire_A_31;
wire RLL_wire_A_32;
wire RLL_wire_A_33;
wire RLL_wire_A_34;
wire RLL_wire_A_35;
wire RLL_wire_A_36;
wire RLL_wire_A_37;
wire RLL_wire_A_38;
wire RLL_wire_A_39;
wire RLL_wire_A_40;
wire RLL_wire_A_41;
wire RLL_wire_A_42;
wire RLL_wire_A_43;
wire RLL_wire_A_44;
wire RLL_wire_A_45;
wire RLL_wire_A_46;
wire RLL_wire_A_47;
wire RLL_wire_A_48;
wire RLL_wire_A_49;
wire RLL_wire_A_50;
wire RLL_wire_A_51;
wire RLL_wire_A_52;
wire RLL_wire_A_53;
wire RLL_wire_A_54;
wire RLL_wire_A_55;
wire RLL_wire_A_56;
wire RLL_wire_A_57;
wire RLL_wire_A_58;
wire RLL_wire_A_59;
wire RLL_wire_A_60;
wire RLL_wire_A_61;
wire RLL_wire_A_62;
wire RLL_wire_A_63;

//Body:
  NOR3_X1   g000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n73_));
  INV_X1    g001(.A(G77), .ZN(new_n74_));
  AND2_X1   g002(.A1(new_n73_), .A2(new_n74_), .ZN(G353));
  OAI21_X1  g003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g004(.A(G1), .ZN(new_n77_));
  INV_X1    g005(.A(G20), .ZN(new_n78_));
  NOR3_X1   g006(.A1(new_n77_), .A2(new_n78_), .A3(G13), .ZN(new_n79_));
  INV_X1    g007(.A(new_n79_), .ZN(new_n80_));
  OAI21_X1  g008(.A(G250), .B1(G257), .B2(G264), .ZN(new_n81_));
  NOR2_X1   g009(.A1(new_n80_), .A2(new_n81_), .ZN(RLL_wire_A_0));
  XNOR2_X1 RLL_XNOR_0 (.A(RLL_wire_A_0), .B(KEYINPUT0), .ZN(new_n82_) );
  AOI22_X1  g010(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n83_));
  INV_X1    g011(.A(G50), .ZN(new_n84_));
  INV_X1    g012(.A(G226), .ZN(new_n85_));
  OAI21_X1  g013(.A(new_n83_), .B1(new_n84_), .B2(new_n85_), .ZN(new_n86_));
  AOI22_X1  g014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n87_));
  NAND2_X1  g015(.A1(G87), .A2(G250), .ZN(new_n88_));
  INV_X1    g016(.A(G97), .ZN(new_n89_));
  INV_X1    g017(.A(G257), .ZN(new_n90_));
  OAI211_X1 g018(.A(new_n87_), .B(new_n88_), .C1(new_n89_), .C2(new_n90_), .ZN(new_n91_));
  AOI211_X1 g019(.A(new_n86_), .B(new_n91_), .C1(G58), .C2(G232), .ZN(new_n92_));
  INV_X1    g020(.A(G13), .ZN(new_n93_));
  NOR3_X1   g021(.A1(new_n77_), .A2(new_n93_), .A3(new_n78_), .ZN(new_n94_));
  NOR3_X1   g022(.A1(new_n92_), .A2(new_n79_), .A3(new_n94_), .ZN(RLL_wire_A_1));
  XOR2_X1 RLL_XOR_1 (.A(RLL_wire_A_1), .B(KEYINPUT1), .Z(new_n95_) );
  OAI21_X1  g023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n96_));
  INV_X1    g024(.A(new_n96_), .ZN(new_n97_));
  AOI211_X1 g025(.A(new_n82_), .B(new_n95_), .C1(new_n94_), .C2(new_n97_), .ZN(G361));
  XOR2_X1   g026(.A(G264), .B(G270), .Z(new_n99_));
  XNOR2_X1  g027(.A(G250), .B(G257), .ZN(new_n100_));
  XNOR2_X1  g028(.A(new_n99_), .B(new_n100_), .ZN(new_n101_));
  XOR2_X1   g029(.A(G238), .B(G244), .Z(RLL_wire_A_2));
  XOR2_X1 RLL_XOR_2 (.A(RLL_wire_A_2), .B(KEYINPUT2), .Z(new_n102_) );
  XNOR2_X1  g030(.A(G226), .B(G232), .ZN(new_n103_));
  XNOR2_X1  g031(.A(new_n102_), .B(new_n103_), .ZN(new_n104_));
  XNOR2_X1  g032(.A(new_n101_), .B(new_n104_), .ZN(G358));
  XOR2_X1   g033(.A(G68), .B(G77), .Z(new_n106_));
  XNOR2_X1  g034(.A(G50), .B(G58), .ZN(new_n107_));
  XNOR2_X1  g035(.A(new_n106_), .B(new_n107_), .ZN(new_n108_));
  XOR2_X1   g036(.A(G107), .B(G116), .Z(new_n109_));
  XNOR2_X1  g037(.A(G87), .B(G97), .ZN(new_n110_));
  XNOR2_X1  g038(.A(new_n109_), .B(new_n110_), .ZN(new_n111_));
  XNOR2_X1  g039(.A(new_n108_), .B(new_n111_), .ZN(G351));
  INV_X1    g040(.A(G33), .ZN(RLL_wire_A_3));
  XOR2_X1 RLL_XOR_3 (.A(RLL_wire_A_3), .B(KEYINPUT3), .Z(new_n113_) );
  INV_X1    g041(.A(G1698), .ZN(new_n114_));
  NAND3_X1  g042(.A1(new_n113_), .A2(new_n114_), .A3(G244), .ZN(RLL_wire_A_4));
  XNOR2_X1 RLL_XNOR_4 (.A(RLL_wire_A_4), .B(KEYINPUT4), .ZN(new_n115_) );
  NAND3_X1  g043(.A1(new_n113_), .A2(G250), .A3(G1698), .ZN(new_n116_));
  NAND2_X1  g044(.A1(G33), .A2(G283), .ZN(new_n117_));
  NAND3_X1  g045(.A1(new_n115_), .A2(new_n116_), .A3(new_n117_), .ZN(new_n118_));
  NAND2_X1  g046(.A1(G33), .A2(G41), .ZN(new_n119_));
  AND3_X1   g047(.A1(new_n119_), .A2(G1), .A3(G13), .ZN(new_n120_));
  NAND2_X1  g048(.A1(new_n118_), .A2(new_n120_), .ZN(new_n121_));
  INV_X1    g049(.A(G41), .ZN(RLL_wire_A_5));
  XOR2_X1 RLL_XOR_5 (.A(RLL_wire_A_5), .B(KEYINPUT5), .Z(new_n122_) );
  NAND3_X1  g050(.A1(new_n77_), .A2(new_n122_), .A3(G45), .ZN(new_n123_));
  INV_X1    g051(.A(new_n123_), .ZN(new_n124_));
  NAND3_X1  g052(.A1(new_n119_), .A2(G1), .A3(G13), .ZN(new_n125_));
  NAND3_X1  g053(.A1(new_n124_), .A2(new_n125_), .A3(G274), .ZN(new_n126_));
  NAND3_X1  g054(.A1(new_n125_), .A2(new_n123_), .A3(G257), .ZN(new_n127_));
  NAND3_X1  g055(.A1(new_n121_), .A2(new_n126_), .A3(new_n127_), .ZN(new_n128_));
  NAND2_X1  g056(.A1(new_n128_), .A2(G200), .ZN(new_n129_));
  NAND3_X1  g057(.A1(new_n77_), .A2(G13), .A3(G20), .ZN(new_n130_));
  INV_X1    g058(.A(new_n130_), .ZN(new_n131_));
  NAND2_X1  g059(.A1(new_n131_), .A2(new_n89_), .ZN(new_n132_));
  NAND3_X1  g060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n133_));
  NAND2_X1  g061(.A1(G1), .A2(G13), .ZN(new_n134_));
  NAND2_X1  g062(.A1(new_n133_), .A2(new_n134_), .ZN(new_n135_));
  NAND2_X1  g063(.A1(new_n89_), .A2(G107), .ZN(new_n136_));
  INV_X1    g064(.A(G107), .ZN(new_n137_));
  NAND2_X1  g065(.A1(new_n137_), .A2(G97), .ZN(RLL_wire_A_6));
  XOR2_X1 RLL_XOR_6 (.A(RLL_wire_A_6), .B(KEYINPUT6), .Z(new_n138_) );
  NAND3_X1  g066(.A1(new_n136_), .A2(new_n138_), .A3(G20), .ZN(new_n139_));
  NOR2_X1   g067(.A1(new_n113_), .A2(G20), .ZN(RLL_wire_A_7));
  XNOR2_X1 RLL_XNOR_7 (.A(RLL_wire_A_7), .B(KEYINPUT7), .ZN(new_n140_) );
  NAND2_X1  g068(.A1(new_n140_), .A2(G107), .ZN(new_n141_));
  NOR2_X1   g069(.A1(G20), .A2(G33), .ZN(new_n142_));
  NAND2_X1  g070(.A1(new_n142_), .A2(G77), .ZN(new_n143_));
  NAND3_X1  g071(.A1(new_n139_), .A2(new_n141_), .A3(new_n143_), .ZN(new_n144_));
  AND4_X1   g072(.A1(G97), .A2(new_n130_), .A3(new_n134_), .A4(new_n133_), .ZN(new_n145_));
  NAND2_X1  g073(.A1(new_n77_), .A2(G33), .ZN(new_n146_));
  AOI22_X1  g074(.A1(new_n135_), .A2(new_n144_), .B1(new_n145_), .B2(new_n146_), .ZN(new_n147_));
  NAND4_X1  g075(.A1(new_n121_), .A2(new_n126_), .A3(G190), .A4(new_n127_), .ZN(new_n148_));
  NAND4_X1  g076(.A1(new_n129_), .A2(new_n132_), .A3(new_n147_), .A4(new_n148_), .ZN(new_n149_));
  NAND2_X1  g077(.A1(new_n144_), .A2(new_n135_), .ZN(new_n150_));
  NAND2_X1  g078(.A1(new_n145_), .A2(new_n146_), .ZN(new_n151_));
  NAND3_X1  g079(.A1(new_n150_), .A2(new_n151_), .A3(new_n132_), .ZN(new_n152_));
  NAND3_X1  g080(.A1(new_n152_), .A2(G169), .A3(new_n128_), .ZN(new_n153_));
  INV_X1    g081(.A(new_n128_), .ZN(new_n154_));
  NAND3_X1  g082(.A1(new_n152_), .A2(G179), .A3(new_n154_), .ZN(new_n155_));
  AND3_X1   g083(.A1(new_n149_), .A2(new_n153_), .A3(new_n155_), .ZN(new_n156_));
  NAND2_X1  g084(.A1(new_n142_), .A2(G150), .ZN(new_n157_));
  NAND2_X1  g085(.A1(new_n78_), .A2(G33), .ZN(new_n158_));
  INV_X1    g086(.A(G58), .ZN(RLL_wire_A_8));
  XOR2_X1 RLL_XOR_8 (.A(RLL_wire_A_8), .B(KEYINPUT8), .Z(new_n159_) );
  OAI221_X1 g087(.A(new_n157_), .B1(new_n158_), .B2(new_n159_), .C1(new_n73_), .C2(new_n78_), .ZN(new_n160_));
  NOR3_X1   g088(.A1(new_n131_), .A2(new_n135_), .A3(new_n84_), .ZN(new_n161_));
  NAND2_X1  g089(.A1(new_n77_), .A2(G20), .ZN(new_n162_));
  AOI22_X1  g090(.A1(new_n135_), .A2(new_n160_), .B1(new_n161_), .B2(new_n162_), .ZN(new_n163_));
  NAND2_X1  g091(.A1(new_n131_), .A2(new_n84_), .ZN(new_n164_));
  NAND2_X1  g092(.A1(new_n163_), .A2(new_n164_), .ZN(new_n165_));
  INV_X1    g093(.A(new_n165_), .ZN(RLL_wire_A_9));
  XOR2_X1 RLL_XOR_9 (.A(RLL_wire_A_9), .B(KEYINPUT9), .Z(new_n166_) );
  NAND3_X1  g094(.A1(new_n113_), .A2(new_n114_), .A3(G222), .ZN(new_n167_));
  INV_X1    g095(.A(G223), .ZN(new_n168_));
  NAND2_X1  g096(.A1(new_n113_), .A2(G1698), .ZN(new_n169_));
  OAI221_X1 g097(.A(new_n167_), .B1(new_n113_), .B2(new_n74_), .C1(new_n168_), .C2(new_n169_), .ZN(new_n170_));
  NAND2_X1  g098(.A1(new_n170_), .A2(new_n120_), .ZN(new_n171_));
  OAI21_X1  g099(.A(new_n77_), .B1(G41), .B2(G45), .ZN(new_n172_));
  NOR2_X1   g100(.A1(new_n120_), .A2(new_n172_), .ZN(new_n173_));
  NAND2_X1  g101(.A1(new_n173_), .A2(G274), .ZN(new_n174_));
  AND2_X1   g102(.A1(new_n125_), .A2(new_n172_), .ZN(new_n175_));
  NAND2_X1  g103(.A1(new_n175_), .A2(G226), .ZN(new_n176_));
  NAND3_X1  g104(.A1(new_n171_), .A2(new_n174_), .A3(new_n176_), .ZN(new_n177_));
  NAND2_X1  g105(.A1(new_n177_), .A2(G200), .ZN(new_n178_));
  INV_X1    g106(.A(G190), .ZN(new_n179_));
  OAI211_X1 g107(.A(new_n166_), .B(new_n178_), .C1(new_n179_), .C2(new_n177_), .ZN(RLL_wire_A_10));
  XNOR2_X1 RLL_XNOR_10 (.A(RLL_wire_A_10), .B(KEYINPUT10), .ZN(new_n180_) );
  AND2_X1   g108(.A1(new_n177_), .A2(G169), .ZN(new_n181_));
  INV_X1    g109(.A(G179), .ZN(new_n182_));
  NOR2_X1   g110(.A1(new_n177_), .A2(new_n182_), .ZN(new_n183_));
  OAI21_X1  g111(.A(new_n165_), .B1(new_n181_), .B2(new_n183_), .ZN(new_n184_));
  NAND2_X1  g112(.A1(new_n180_), .A2(new_n184_), .ZN(new_n185_));
  INV_X1    g113(.A(new_n142_), .ZN(new_n186_));
  OAI22_X1  g114(.A1(new_n186_), .A2(new_n84_), .B1(new_n78_), .B2(G68), .ZN(new_n187_));
  NOR2_X1   g115(.A1(new_n158_), .A2(new_n74_), .ZN(new_n188_));
  OAI21_X1  g116(.A(new_n135_), .B1(new_n187_), .B2(new_n188_), .ZN(RLL_wire_A_11));
  XNOR2_X1 RLL_XNOR_11 (.A(RLL_wire_A_11), .B(KEYINPUT11), .ZN(new_n189_) );
  NOR2_X1   g117(.A1(new_n131_), .A2(new_n135_), .ZN(new_n190_));
  NAND3_X1  g118(.A1(new_n190_), .A2(G68), .A3(new_n162_), .ZN(new_n191_));
  INV_X1    g119(.A(G68), .ZN(new_n192_));
  NAND2_X1  g120(.A1(new_n131_), .A2(new_n192_), .ZN(RLL_wire_A_12));
  XNOR2_X1 RLL_XNOR_12 (.A(RLL_wire_A_12), .B(KEYINPUT12), .ZN(new_n193_) );
  NAND3_X1  g121(.A1(new_n189_), .A2(new_n191_), .A3(new_n193_), .ZN(new_n194_));
  NAND2_X1  g122(.A1(G33), .A2(G97), .ZN(new_n195_));
  INV_X1    g123(.A(G232), .ZN(new_n196_));
  NAND2_X1  g124(.A1(new_n113_), .A2(new_n114_), .ZN(new_n197_));
  OAI221_X1 g125(.A(new_n195_), .B1(new_n169_), .B2(new_n196_), .C1(new_n85_), .C2(new_n197_), .ZN(new_n198_));
  NAND2_X1  g126(.A1(new_n198_), .A2(new_n120_), .ZN(new_n199_));
  NAND2_X1  g127(.A1(new_n175_), .A2(G238), .ZN(new_n200_));
  NAND3_X1  g128(.A1(new_n199_), .A2(new_n174_), .A3(new_n200_), .ZN(RLL_wire_A_13));
  XNOR2_X1 RLL_XNOR_13 (.A(RLL_wire_A_13), .B(KEYINPUT13), .ZN(new_n201_) );
  AND2_X1   g129(.A1(new_n201_), .A2(G169), .ZN(RLL_wire_A_14));
  XOR2_X1 RLL_XOR_14 (.A(RLL_wire_A_14), .B(KEYINPUT14), .Z(new_n202_) );
  NOR2_X1   g130(.A1(new_n201_), .A2(new_n182_), .ZN(new_n203_));
  OAI21_X1  g131(.A(new_n194_), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g132(.A1(new_n201_), .A2(G200), .ZN(new_n205_));
  INV_X1    g133(.A(new_n194_), .ZN(new_n206_));
  OAI211_X1 g134(.A(new_n205_), .B(new_n206_), .C1(new_n179_), .C2(new_n201_), .ZN(new_n207_));
  NAND2_X1  g135(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  OAI22_X1  g136(.A1(new_n186_), .A2(new_n159_), .B1(new_n78_), .B2(new_n74_), .ZN(new_n209_));
  INV_X1    g137(.A(G87), .ZN(RLL_wire_A_15));
  XOR2_X1 RLL_XOR_15 (.A(RLL_wire_A_15), .B(KEYINPUT15), .Z(new_n210_) );
  NOR2_X1   g138(.A1(new_n158_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g139(.A(new_n135_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g140(.A1(new_n190_), .A2(G77), .A3(new_n162_), .ZN(new_n213_));
  NAND2_X1  g141(.A1(new_n131_), .A2(new_n74_), .ZN(new_n214_));
  AND3_X1   g142(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND3_X1  g143(.A1(new_n113_), .A2(G238), .A3(G1698), .ZN(new_n216_));
  OAI221_X1 g144(.A(new_n216_), .B1(new_n113_), .B2(new_n137_), .C1(new_n197_), .C2(new_n196_), .ZN(new_n217_));
  NAND2_X1  g145(.A1(new_n217_), .A2(new_n120_), .ZN(new_n218_));
  NAND2_X1  g146(.A1(new_n175_), .A2(G244), .ZN(new_n219_));
  NAND3_X1  g147(.A1(new_n218_), .A2(new_n174_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g148(.A1(new_n220_), .A2(G169), .ZN(new_n221_));
  NAND4_X1  g149(.A1(new_n218_), .A2(new_n174_), .A3(G179), .A4(new_n219_), .ZN(new_n222_));
  AOI21_X1  g150(.A(new_n215_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g151(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g152(.A1(new_n220_), .A2(G200), .ZN(new_n225_));
  NAND4_X1  g153(.A1(new_n218_), .A2(new_n174_), .A3(G190), .A4(new_n219_), .ZN(new_n226_));
  NAND3_X1  g154(.A1(new_n225_), .A2(new_n215_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g155(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NOR3_X1   g156(.A1(new_n185_), .A2(new_n208_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g157(.A1(new_n131_), .A2(new_n159_), .ZN(new_n230_));
  NAND2_X1  g158(.A1(G33), .A2(G87), .ZN(new_n231_));
  OAI221_X1 g159(.A(new_n231_), .B1(new_n169_), .B2(new_n85_), .C1(new_n168_), .C2(new_n197_), .ZN(new_n232_));
  NAND2_X1  g160(.A1(new_n232_), .A2(new_n120_), .ZN(new_n233_));
  NAND2_X1  g161(.A1(new_n175_), .A2(G232), .ZN(new_n234_));
  NAND3_X1  g162(.A1(new_n233_), .A2(new_n174_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g163(.A1(new_n235_), .A2(G200), .ZN(new_n236_));
  NAND2_X1  g164(.A1(new_n140_), .A2(G68), .ZN(new_n237_));
  INV_X1    g165(.A(G159), .ZN(new_n238_));
  XOR2_X1   g166(.A(G58), .B(G68), .Z(new_n239_));
  OAI221_X1 g167(.A(new_n237_), .B1(new_n238_), .B2(new_n186_), .C1(new_n239_), .C2(new_n78_), .ZN(RLL_wire_A_16));
  XNOR2_X1 RLL_XNOR_16 (.A(RLL_wire_A_16), .B(KEYINPUT16), .ZN(new_n240_) );
  NOR3_X1   g168(.A1(new_n131_), .A2(new_n135_), .A3(new_n159_), .ZN(new_n241_));
  AOI22_X1  g169(.A1(new_n240_), .A2(new_n135_), .B1(new_n241_), .B2(new_n162_), .ZN(new_n242_));
  NAND4_X1  g170(.A1(new_n233_), .A2(new_n234_), .A3(G190), .A4(new_n174_), .ZN(new_n243_));
  AND4_X1   g171(.A1(new_n230_), .A2(new_n236_), .A3(new_n242_), .A4(new_n243_), .ZN(RLL_wire_A_17));
  XNOR2_X1 RLL_XNOR_17 (.A(RLL_wire_A_17), .B(KEYINPUT17), .ZN(new_n244_) );
  NAND2_X1  g172(.A1(new_n235_), .A2(G169), .ZN(new_n245_));
  NAND4_X1  g173(.A1(new_n233_), .A2(new_n234_), .A3(G179), .A4(new_n174_), .ZN(new_n246_));
  AOI22_X1  g174(.A1(new_n245_), .A2(new_n246_), .B1(new_n242_), .B2(new_n230_), .ZN(RLL_wire_A_18));
  XOR2_X1 RLL_XOR_18 (.A(RLL_wire_A_18), .B(KEYINPUT18), .Z(new_n247_) );
  NOR2_X1   g175(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  AND2_X1   g176(.A1(new_n229_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g177(.A1(new_n78_), .A2(G33), .A3(G97), .ZN(RLL_wire_A_19));
  XNOR2_X1 RLL_XNOR_19 (.A(RLL_wire_A_19), .B(KEYINPUT19), .ZN(new_n250_) );
  NAND3_X1  g178(.A1(new_n78_), .A2(new_n113_), .A3(G68), .ZN(new_n251_));
  NOR3_X1   g179(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n252_));
  OAI211_X1 g180(.A(new_n250_), .B(new_n251_), .C1(new_n252_), .C2(new_n78_), .ZN(new_n253_));
  NAND2_X1  g181(.A1(new_n253_), .A2(new_n135_), .ZN(new_n254_));
  NAND2_X1  g182(.A1(new_n131_), .A2(new_n210_), .ZN(new_n255_));
  INV_X1    g183(.A(new_n135_), .ZN(new_n256_));
  NAND4_X1  g184(.A1(new_n256_), .A2(G87), .A3(new_n130_), .A4(new_n146_), .ZN(new_n257_));
  AND3_X1   g185(.A1(new_n254_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g186(.A1(new_n113_), .A2(new_n114_), .A3(G238), .ZN(new_n259_));
  NAND3_X1  g187(.A1(new_n113_), .A2(G244), .A3(G1698), .ZN(new_n260_));
  NAND2_X1  g188(.A1(G33), .A2(G116), .ZN(new_n261_));
  NAND3_X1  g189(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g190(.A1(new_n262_), .A2(new_n120_), .ZN(new_n263_));
  NAND4_X1  g191(.A1(new_n125_), .A2(new_n77_), .A3(G45), .A4(G274), .ZN(new_n264_));
  INV_X1    g192(.A(G45), .ZN(new_n265_));
  OAI211_X1 g193(.A(new_n125_), .B(G250), .C1(G1), .C2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g194(.A1(new_n263_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g195(.A1(new_n267_), .A2(G200), .ZN(new_n268_));
  NAND4_X1  g196(.A1(new_n263_), .A2(new_n264_), .A3(G190), .A4(new_n266_), .ZN(new_n269_));
  AND3_X1   g197(.A1(new_n258_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g198(.A1(new_n267_), .A2(G169), .ZN(new_n271_));
  NAND4_X1  g199(.A1(new_n263_), .A2(new_n264_), .A3(G179), .A4(new_n266_), .ZN(new_n272_));
  NOR3_X1   g200(.A1(new_n131_), .A2(new_n135_), .A3(new_n210_), .ZN(new_n273_));
  AOI22_X1  g201(.A1(new_n273_), .A2(new_n146_), .B1(new_n253_), .B2(new_n135_), .ZN(new_n274_));
  AOI22_X1  g202(.A1(new_n271_), .A2(new_n272_), .B1(new_n274_), .B2(new_n255_), .ZN(new_n275_));
  NOR2_X1   g203(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g204(.A1(new_n113_), .A2(G264), .A3(G1698), .ZN(new_n277_));
  INV_X1    g205(.A(G303), .ZN(new_n278_));
  OAI221_X1 g206(.A(new_n277_), .B1(new_n113_), .B2(new_n278_), .C1(new_n197_), .C2(new_n90_), .ZN(new_n279_));
  NAND2_X1  g207(.A1(new_n279_), .A2(new_n120_), .ZN(new_n280_));
  NAND3_X1  g208(.A1(new_n125_), .A2(new_n123_), .A3(G270), .ZN(new_n281_));
  NAND4_X1  g209(.A1(new_n280_), .A2(G179), .A3(new_n126_), .A4(new_n281_), .ZN(new_n282_));
  INV_X1    g210(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g211(.A(G116), .ZN(new_n284_));
  OAI22_X1  g212(.A1(new_n186_), .A2(new_n89_), .B1(new_n78_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g213(.A(G283), .ZN(new_n286_));
  NOR2_X1   g214(.A1(new_n158_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g215(.A(new_n135_), .B1(new_n285_), .B2(new_n287_), .ZN(RLL_wire_A_20));
  XOR2_X1 RLL_XOR_20 (.A(RLL_wire_A_20), .B(KEYINPUT20), .Z(new_n288_) );
  NAND3_X1  g216(.A1(new_n190_), .A2(G116), .A3(new_n146_), .ZN(new_n289_));
  NAND2_X1  g217(.A1(new_n131_), .A2(new_n284_), .ZN(new_n290_));
  NAND3_X1  g218(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g219(.A1(new_n283_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g220(.A1(new_n280_), .A2(new_n126_), .A3(new_n281_), .ZN(new_n293_));
  NAND3_X1  g221(.A1(new_n291_), .A2(new_n293_), .A3(G169), .ZN(RLL_wire_A_21));
  XNOR2_X1 RLL_XNOR_21 (.A(RLL_wire_A_21), .B(KEYINPUT21), .ZN(new_n294_) );
  NAND2_X1  g222(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g223(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g224(.A1(new_n293_), .A2(G200), .ZN(new_n297_));
  INV_X1    g225(.A(new_n291_), .ZN(new_n298_));
  OAI211_X1 g226(.A(new_n297_), .B(new_n298_), .C1(new_n179_), .C2(new_n293_), .ZN(new_n299_));
  NAND3_X1  g227(.A1(new_n113_), .A2(new_n114_), .A3(G250), .ZN(new_n300_));
  NAND3_X1  g228(.A1(new_n113_), .A2(G257), .A3(G1698), .ZN(new_n301_));
  NAND2_X1  g229(.A1(G33), .A2(G294), .ZN(new_n302_));
  NAND3_X1  g230(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g231(.A1(new_n303_), .A2(new_n120_), .ZN(new_n304_));
  NAND3_X1  g232(.A1(new_n125_), .A2(new_n123_), .A3(G264), .ZN(new_n305_));
  NAND3_X1  g233(.A1(new_n304_), .A2(new_n126_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g234(.A1(new_n306_), .A2(G200), .ZN(new_n307_));
  NAND4_X1  g235(.A1(new_n256_), .A2(G107), .A3(new_n130_), .A4(new_n146_), .ZN(new_n308_));
  NAND3_X1  g236(.A1(new_n78_), .A2(new_n113_), .A3(G87), .ZN(RLL_wire_A_22));
  XNOR2_X1 RLL_XNOR_22 (.A(RLL_wire_A_22), .B(KEYINPUT22), .ZN(new_n309_) );
  NAND3_X1  g237(.A1(new_n78_), .A2(G33), .A3(G116), .ZN(new_n310_));
  NAND2_X1  g238(.A1(new_n137_), .A2(G20), .ZN(RLL_wire_A_23));
  XOR2_X1 RLL_XOR_23 (.A(RLL_wire_A_23), .B(KEYINPUT23), .Z(new_n311_) );
  NAND3_X1  g239(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(RLL_wire_A_24));
  XNOR2_X1 RLL_XNOR_24 (.A(RLL_wire_A_24), .B(KEYINPUT24), .ZN(new_n312_) );
  NAND2_X1  g240(.A1(new_n312_), .A2(new_n135_), .ZN(new_n313_));
  NAND2_X1  g241(.A1(new_n131_), .A2(new_n137_), .ZN(RLL_wire_A_25));
  XOR2_X1 RLL_XOR_25 (.A(RLL_wire_A_25), .B(KEYINPUT25), .Z(new_n314_) );
  AND3_X1   g242(.A1(new_n308_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  NAND4_X1  g243(.A1(new_n304_), .A2(new_n126_), .A3(G190), .A4(new_n305_), .ZN(new_n316_));
  AND3_X1   g244(.A1(new_n307_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g245(.A1(new_n306_), .A2(G169), .ZN(new_n318_));
  NAND4_X1  g246(.A1(new_n304_), .A2(new_n126_), .A3(G179), .A4(new_n305_), .ZN(new_n319_));
  AOI21_X1  g247(.A(new_n315_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g248(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  AND3_X1   g249(.A1(new_n296_), .A2(new_n299_), .A3(new_n321_), .ZN(new_n322_));
  AND4_X1   g250(.A1(new_n156_), .A2(new_n249_), .A3(new_n276_), .A4(new_n322_), .ZN(G372));
  NOR2_X1   g251(.A1(new_n185_), .A2(new_n208_), .ZN(new_n324_));
  NAND3_X1  g252(.A1(new_n324_), .A2(new_n248_), .A3(new_n223_), .ZN(new_n325_));
  INV_X1    g253(.A(new_n185_), .ZN(new_n326_));
  NAND2_X1  g254(.A1(new_n326_), .A2(new_n247_), .ZN(new_n327_));
  INV_X1    g255(.A(new_n204_), .ZN(new_n328_));
  NAND3_X1  g256(.A1(new_n326_), .A2(new_n248_), .A3(new_n328_), .ZN(new_n329_));
  AND4_X1   g257(.A1(new_n184_), .A2(new_n325_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n330_));
  NAND4_X1  g258(.A1(new_n156_), .A2(new_n276_), .A3(new_n321_), .A4(new_n295_), .ZN(new_n331_));
  NAND3_X1  g259(.A1(new_n156_), .A2(new_n276_), .A3(new_n320_), .ZN(new_n332_));
  INV_X1    g260(.A(new_n275_), .ZN(new_n333_));
  NAND2_X1  g261(.A1(new_n153_), .A2(new_n155_), .ZN(new_n334_));
  NAND2_X1  g262(.A1(new_n276_), .A2(new_n334_), .ZN(RLL_wire_A_26));
  XOR2_X1 RLL_XOR_26 (.A(RLL_wire_A_26), .B(KEYINPUT26), .Z(new_n335_) );
  NAND4_X1  g263(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .A4(new_n335_), .ZN(new_n336_));
  NAND2_X1  g264(.A1(new_n249_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g265(.A1(new_n330_), .A2(new_n337_), .ZN(G369));
  NOR3_X1   g266(.A1(new_n93_), .A2(G1), .A3(G20), .ZN(RLL_wire_A_27));
  XNOR2_X1 RLL_XNOR_27 (.A(RLL_wire_A_27), .B(KEYINPUT27), .ZN(new_n339_) );
  NAND3_X1  g267(.A1(new_n339_), .A2(G213), .A3(G343), .ZN(new_n340_));
  AND2_X1   g268(.A1(new_n320_), .A2(new_n340_), .ZN(new_n341_));
  OR2_X1    g269(.A1(new_n315_), .A2(new_n340_), .ZN(new_n342_));
  XNOR2_X1  g270(.A(new_n321_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g271(.A(new_n340_), .ZN(new_n344_));
  NOR2_X1   g272(.A1(new_n296_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g273(.A(new_n341_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g274(.A1(new_n296_), .A2(new_n299_), .ZN(new_n347_));
  NOR2_X1   g275(.A1(new_n298_), .A2(new_n340_), .ZN(new_n348_));
  XNOR2_X1  g276(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g277(.A1(new_n349_), .A2(new_n343_), .ZN(new_n350_));
  INV_X1    g278(.A(G330), .ZN(new_n351_));
  OAI21_X1  g279(.A(new_n346_), .B1(new_n350_), .B2(new_n351_), .ZN(G399));
  NOR4_X1   g280(.A1(new_n77_), .A2(new_n78_), .A3(G13), .A4(G41), .ZN(new_n353_));
  NOR2_X1   g281(.A1(new_n353_), .A2(new_n77_), .ZN(new_n354_));
  AND2_X1   g282(.A1(new_n252_), .A2(new_n284_), .ZN(new_n355_));
  AOI22_X1  g283(.A1(new_n354_), .A2(new_n355_), .B1(new_n97_), .B2(new_n353_), .ZN(RLL_wire_A_28));
  XOR2_X1 RLL_XOR_28 (.A(RLL_wire_A_28), .B(KEYINPUT28), .Z(new_n356_) );
  NAND2_X1  g284(.A1(new_n336_), .A2(new_n340_), .ZN(new_n357_));
  INV_X1    g285(.A(new_n357_), .ZN(RLL_wire_A_29));
  XOR2_X1 RLL_XOR_29 (.A(RLL_wire_A_29), .B(KEYINPUT29), .Z(new_n358_) );
  NAND4_X1  g286(.A1(new_n322_), .A2(new_n156_), .A3(new_n276_), .A4(new_n340_), .ZN(new_n359_));
  NAND4_X1  g287(.A1(new_n293_), .A2(new_n182_), .A3(new_n267_), .A4(new_n306_), .ZN(new_n360_));
  NOR2_X1   g288(.A1(new_n360_), .A2(new_n154_), .ZN(new_n361_));
  NOR4_X1   g289(.A1(new_n282_), .A2(new_n128_), .A3(new_n267_), .A4(new_n306_), .ZN(RLL_wire_A_30));
  XNOR2_X1 RLL_XNOR_30 (.A(RLL_wire_A_30), .B(KEYINPUT30), .ZN(new_n362_) );
  OAI21_X1  g290(.A(new_n344_), .B1(new_n361_), .B2(new_n362_), .ZN(RLL_wire_A_31));
  XNOR2_X1 RLL_XNOR_31 (.A(RLL_wire_A_31), .B(KEYINPUT31), .ZN(new_n363_) );
  NAND2_X1  g291(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g292(.A(new_n358_), .B1(new_n364_), .B2(G330), .ZN(new_n365_));
  OAI21_X1  g293(.A(new_n356_), .B1(new_n365_), .B2(G1), .ZN(G364));
  XNOR2_X1  g294(.A(new_n349_), .B(G330), .ZN(new_n367_));
  INV_X1    g295(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g296(.A1(new_n368_), .A2(new_n353_), .ZN(new_n369_));
  NOR2_X1   g297(.A1(new_n93_), .A2(new_n265_), .ZN(new_n370_));
  AOI21_X1  g298(.A(new_n77_), .B1(new_n370_), .B2(new_n78_), .ZN(new_n371_));
  INV_X1    g299(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g300(.A1(new_n368_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g301(.A1(new_n179_), .A2(G20), .ZN(new_n374_));
  OAI21_X1  g302(.A(G20), .B1(G179), .B2(G200), .ZN(new_n375_));
  NAND2_X1  g303(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g304(.A1(new_n376_), .A2(new_n89_), .ZN(new_n377_));
  INV_X1    g305(.A(new_n374_), .ZN(new_n378_));
  NAND2_X1  g306(.A1(G20), .A2(G179), .ZN(new_n379_));
  NOR3_X1   g307(.A1(new_n378_), .A2(G200), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g308(.A(G200), .ZN(new_n381_));
  NOR2_X1   g309(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  AND2_X1   g310(.A1(new_n382_), .A2(new_n374_), .ZN(new_n383_));
  AOI22_X1  g311(.A1(new_n380_), .A2(G58), .B1(new_n383_), .B2(G50), .ZN(new_n384_));
  NAND2_X1  g312(.A1(new_n378_), .A2(new_n382_), .ZN(new_n385_));
  NAND4_X1  g313(.A1(new_n179_), .A2(new_n381_), .A3(G20), .A4(G179), .ZN(new_n386_));
  OAI221_X1 g314(.A(new_n384_), .B1(new_n192_), .B2(new_n385_), .C1(new_n74_), .C2(new_n386_), .ZN(new_n387_));
  NOR4_X1   g315(.A1(new_n78_), .A2(new_n179_), .A3(new_n381_), .A4(G179), .ZN(new_n388_));
  AOI211_X1 g316(.A(new_n377_), .B(new_n387_), .C1(G87), .C2(new_n388_), .ZN(new_n389_));
  NOR4_X1   g317(.A1(new_n78_), .A2(new_n381_), .A3(G179), .A4(G190), .ZN(new_n390_));
  NAND2_X1  g318(.A1(new_n390_), .A2(G107), .ZN(new_n391_));
  AND2_X1   g319(.A1(new_n378_), .A2(new_n375_), .ZN(new_n392_));
  NAND2_X1  g320(.A1(new_n392_), .A2(G159), .ZN(RLL_wire_A_32));
  XOR2_X1 RLL_XOR_32 (.A(RLL_wire_A_32), .B(KEYINPUT32), .Z(new_n393_) );
  NAND4_X1  g321(.A1(new_n389_), .A2(new_n113_), .A3(new_n391_), .A4(new_n393_), .ZN(new_n394_));
  INV_X1    g322(.A(new_n388_), .ZN(new_n395_));
  NOR2_X1   g323(.A1(new_n395_), .A2(new_n278_), .ZN(new_n396_));
  AOI22_X1  g324(.A1(new_n380_), .A2(G322), .B1(new_n383_), .B2(G326), .ZN(new_n397_));
  INV_X1    g325(.A(G311), .ZN(new_n398_));
  INV_X1    g326(.A(G317), .ZN(RLL_wire_A_33));
  XNOR2_X1 RLL_XNOR_33 (.A(RLL_wire_A_33), .B(KEYINPUT33), .ZN(new_n399_) );
  OAI221_X1 g327(.A(new_n397_), .B1(new_n398_), .B2(new_n386_), .C1(new_n399_), .C2(new_n385_), .ZN(new_n400_));
  INV_X1    g328(.A(new_n376_), .ZN(new_n401_));
  AOI211_X1 g329(.A(new_n396_), .B(new_n400_), .C1(G294), .C2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g330(.A1(new_n390_), .A2(G283), .ZN(new_n403_));
  NAND2_X1  g331(.A1(new_n392_), .A2(G329), .ZN(new_n404_));
  NAND3_X1  g332(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g333(.A(new_n394_), .B1(new_n405_), .B2(new_n113_), .ZN(new_n406_));
  OAI211_X1 g334(.A(G1), .B(G13), .C1(new_n78_), .C2(G169), .ZN(new_n407_));
  INV_X1    g335(.A(new_n407_), .ZN(new_n408_));
  NOR2_X1   g336(.A1(new_n80_), .A2(new_n113_), .ZN(new_n409_));
  NAND2_X1  g337(.A1(new_n97_), .A2(new_n265_), .ZN(new_n410_));
  OAI211_X1 g338(.A(new_n409_), .B(new_n410_), .C1(new_n108_), .C2(new_n265_), .ZN(new_n411_));
  NAND3_X1  g339(.A1(new_n93_), .A2(G1), .A3(G20), .ZN(new_n412_));
  INV_X1    g340(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g341(.A(G355), .ZN(new_n414_));
  NAND2_X1  g342(.A1(new_n79_), .A2(new_n113_), .ZN(new_n415_));
  OAI221_X1 g343(.A(new_n411_), .B1(G116), .B2(new_n413_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g344(.A1(G13), .A2(G33), .ZN(new_n417_));
  INV_X1    g345(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g346(.A1(new_n418_), .A2(G20), .ZN(new_n419_));
  NOR2_X1   g347(.A1(new_n419_), .A2(new_n408_), .ZN(new_n420_));
  AOI22_X1  g348(.A1(new_n406_), .A2(new_n408_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g349(.A1(new_n372_), .A2(new_n353_), .ZN(new_n422_));
  INV_X1    g350(.A(new_n419_), .ZN(new_n423_));
  OAI211_X1 g351(.A(new_n421_), .B(new_n422_), .C1(new_n349_), .C2(new_n423_), .ZN(new_n424_));
  AND3_X1   g352(.A1(new_n369_), .A2(new_n373_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g353(.A(new_n425_), .ZN(G396));
  OAI211_X1 g354(.A(new_n224_), .B(new_n227_), .C1(new_n215_), .C2(new_n340_), .ZN(new_n427_));
  NOR2_X1   g355(.A1(new_n215_), .A2(new_n340_), .ZN(new_n428_));
  INV_X1    g356(.A(new_n227_), .ZN(new_n429_));
  OAI21_X1  g357(.A(new_n428_), .B1(new_n429_), .B2(new_n223_), .ZN(new_n430_));
  NAND2_X1  g358(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g359(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g360(.A(new_n357_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g361(.A(new_n364_), .ZN(new_n434_));
  NOR2_X1   g362(.A1(new_n434_), .A2(new_n351_), .ZN(new_n435_));
  AND2_X1   g363(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g364(.A1(new_n433_), .A2(new_n435_), .ZN(new_n437_));
  OAI21_X1  g365(.A(new_n353_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g366(.A(new_n372_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n439_));
  NOR2_X1   g367(.A1(new_n395_), .A2(new_n84_), .ZN(new_n440_));
  AOI22_X1  g368(.A1(new_n380_), .A2(G143), .B1(new_n383_), .B2(G137), .ZN(new_n441_));
  INV_X1    g369(.A(G150), .ZN(new_n442_));
  OAI221_X1 g370(.A(new_n441_), .B1(new_n442_), .B2(new_n385_), .C1(new_n238_), .C2(new_n386_), .ZN(RLL_wire_A_34));
  XOR2_X1 RLL_XOR_34 (.A(RLL_wire_A_34), .B(KEYINPUT34), .Z(new_n443_) );
  AOI211_X1 g371(.A(new_n440_), .B(new_n443_), .C1(G58), .C2(new_n401_), .ZN(new_n444_));
  NAND2_X1  g372(.A1(new_n390_), .A2(G68), .ZN(new_n445_));
  NAND2_X1  g373(.A1(new_n392_), .A2(G132), .ZN(new_n446_));
  NAND4_X1  g374(.A1(new_n444_), .A2(new_n113_), .A3(new_n445_), .A4(new_n446_), .ZN(new_n447_));
  AOI22_X1  g375(.A1(new_n380_), .A2(G294), .B1(new_n383_), .B2(G303), .ZN(new_n448_));
  OAI221_X1 g376(.A(new_n448_), .B1(new_n284_), .B2(new_n386_), .C1(new_n286_), .C2(new_n385_), .ZN(new_n449_));
  AOI211_X1 g377(.A(new_n377_), .B(new_n449_), .C1(G107), .C2(new_n388_), .ZN(new_n450_));
  NAND2_X1  g378(.A1(new_n390_), .A2(G87), .ZN(new_n451_));
  NAND2_X1  g379(.A1(new_n392_), .A2(G311), .ZN(new_n452_));
  NAND3_X1  g380(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  OAI21_X1  g381(.A(new_n447_), .B1(new_n453_), .B2(new_n113_), .ZN(new_n454_));
  NOR2_X1   g382(.A1(new_n408_), .A2(new_n417_), .ZN(new_n455_));
  AOI22_X1  g383(.A1(new_n454_), .A2(new_n408_), .B1(new_n74_), .B2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g384(.A(new_n456_), .B(new_n422_), .C1(new_n418_), .C2(new_n431_), .ZN(new_n457_));
  NAND3_X1  g385(.A1(new_n438_), .A2(new_n439_), .A3(new_n457_), .ZN(G384));
  NAND2_X1  g386(.A1(new_n136_), .A2(new_n138_), .ZN(RLL_wire_A_35));
  XNOR2_X1 RLL_XNOR_35 (.A(RLL_wire_A_35), .B(KEYINPUT35), .ZN(new_n459_) );
  NAND3_X1  g387(.A1(new_n94_), .A2(new_n459_), .A3(G116), .ZN(RLL_wire_A_36));
  XNOR2_X1 RLL_XNOR_36 (.A(RLL_wire_A_36), .B(KEYINPUT36), .ZN(new_n460_) );
  AND3_X1   g388(.A1(new_n239_), .A2(G50), .A3(G77), .ZN(new_n461_));
  NOR2_X1   g389(.A1(new_n192_), .A2(G50), .ZN(new_n462_));
  OAI211_X1 g390(.A(G1), .B(new_n93_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g391(.A1(new_n339_), .A2(G213), .ZN(new_n464_));
  NAND2_X1  g392(.A1(new_n247_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g393(.A1(new_n194_), .A2(new_n344_), .ZN(new_n466_));
  INV_X1    g394(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g395(.A1(new_n208_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g396(.A1(new_n204_), .A2(new_n207_), .A3(new_n466_), .ZN(new_n469_));
  NAND2_X1  g397(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g398(.A1(new_n242_), .A2(new_n230_), .ZN(new_n471_));
  INV_X1    g399(.A(new_n464_), .ZN(new_n472_));
  NAND2_X1  g400(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g401(.A(new_n473_), .ZN(new_n474_));
  OAI21_X1  g402(.A(new_n474_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n475_));
  INV_X1    g403(.A(new_n471_), .ZN(new_n476_));
  NAND3_X1  g404(.A1(new_n476_), .A2(new_n236_), .A3(new_n243_), .ZN(new_n477_));
  AND2_X1   g405(.A1(new_n235_), .A2(G169), .ZN(new_n478_));
  INV_X1    g406(.A(new_n246_), .ZN(new_n479_));
  OAI21_X1  g407(.A(new_n471_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g408(.A1(new_n477_), .A2(new_n480_), .A3(new_n473_), .ZN(RLL_wire_A_37));
  XNOR2_X1 RLL_XNOR_37 (.A(RLL_wire_A_37), .B(KEYINPUT37), .ZN(new_n481_) );
  NAND2_X1  g409(.A1(new_n475_), .A2(new_n481_), .ZN(RLL_wire_A_38));
  XOR2_X1 RLL_XOR_38 (.A(RLL_wire_A_38), .B(KEYINPUT38), .Z(new_n482_) );
  NOR2_X1   g410(.A1(new_n224_), .A2(new_n344_), .ZN(new_n483_));
  NAND3_X1  g411(.A1(new_n470_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND4_X1  g412(.A1(new_n336_), .A2(new_n340_), .A3(new_n431_), .A4(new_n482_), .ZN(new_n485_));
  INV_X1    g413(.A(new_n470_), .ZN(new_n486_));
  OAI211_X1 g414(.A(new_n465_), .B(new_n484_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  INV_X1    g415(.A(new_n482_), .ZN(RLL_wire_A_39));
  XNOR2_X1 RLL_XNOR_39 (.A(RLL_wire_A_39), .B(KEYINPUT39), .ZN(new_n488_) );
  NOR2_X1   g416(.A1(new_n204_), .A2(new_n344_), .ZN(new_n489_));
  INV_X1    g417(.A(new_n489_), .ZN(new_n490_));
  NOR2_X1   g418(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g419(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g420(.A1(new_n358_), .A2(new_n249_), .ZN(new_n493_));
  NAND2_X1  g421(.A1(new_n330_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g422(.A(new_n492_), .B(new_n494_), .ZN(new_n495_));
  NAND4_X1  g423(.A1(new_n364_), .A2(new_n431_), .A3(new_n482_), .A4(new_n470_), .ZN(RLL_wire_A_40));
  XOR2_X1 RLL_XOR_40 (.A(RLL_wire_A_40), .B(KEYINPUT40), .Z(new_n496_) );
  NAND2_X1  g424(.A1(new_n249_), .A2(new_n364_), .ZN(new_n497_));
  XNOR2_X1  g425(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NOR2_X1   g426(.A1(new_n498_), .A2(new_n351_), .ZN(new_n499_));
  XNOR2_X1  g427(.A(new_n495_), .B(new_n499_), .ZN(new_n500_));
  AOI21_X1  g428(.A(new_n77_), .B1(G13), .B2(new_n78_), .ZN(new_n501_));
  OAI211_X1 g429(.A(new_n460_), .B(new_n463_), .C1(new_n500_), .C2(new_n501_), .ZN(G367));
  INV_X1    g430(.A(new_n353_), .ZN(RLL_wire_A_41));
  XNOR2_X1 RLL_XNOR_41 (.A(RLL_wire_A_41), .B(KEYINPUT41), .ZN(new_n503_) );
  NAND3_X1  g431(.A1(new_n149_), .A2(new_n153_), .A3(new_n155_), .ZN(new_n504_));
  NAND2_X1  g432(.A1(new_n152_), .A2(new_n344_), .ZN(new_n505_));
  INV_X1    g433(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g434(.A(new_n504_), .B(new_n506_), .ZN(new_n507_));
  NAND3_X1  g435(.A1(new_n343_), .A2(new_n345_), .A3(new_n507_), .ZN(RLL_wire_A_42));
  XOR2_X1 RLL_XOR_42 (.A(RLL_wire_A_42), .B(KEYINPUT42), .Z(new_n508_) );
  NAND2_X1  g436(.A1(new_n507_), .A2(new_n341_), .ZN(new_n509_));
  NAND2_X1  g437(.A1(new_n334_), .A2(new_n340_), .ZN(new_n510_));
  NAND3_X1  g438(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NOR2_X1   g439(.A1(new_n258_), .A2(new_n340_), .ZN(new_n512_));
  XOR2_X1   g440(.A(new_n276_), .B(new_n512_), .Z(new_n513_));
  INV_X1    g441(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g442(.A1(new_n511_), .A2(new_n514_), .ZN(RLL_wire_A_43));
  XOR2_X1 RLL_XOR_43 (.A(RLL_wire_A_43), .B(KEYINPUT43), .Z(new_n515_) );
  INV_X1    g443(.A(new_n515_), .ZN(new_n516_));
  NAND4_X1  g444(.A1(new_n349_), .A2(G330), .A3(new_n343_), .A4(new_n507_), .ZN(new_n517_));
  NOR2_X1   g445(.A1(new_n511_), .A2(new_n514_), .ZN(new_n518_));
  OR3_X1    g446(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g447(.A(new_n517_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n520_));
  NAND2_X1  g448(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g449(.A1(new_n350_), .A2(new_n351_), .ZN(new_n522_));
  OR2_X1    g450(.A1(new_n346_), .A2(new_n507_), .ZN(RLL_wire_A_44));
  XOR2_X1 RLL_XOR_44 (.A(RLL_wire_A_44), .B(KEYINPUT44), .Z(new_n523_) );
  NAND2_X1  g451(.A1(new_n346_), .A2(new_n507_), .ZN(RLL_wire_A_45));
  XOR2_X1 RLL_XOR_45 (.A(RLL_wire_A_45), .B(KEYINPUT45), .Z(new_n524_) );
  NAND3_X1  g452(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g453(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g454(.A(new_n522_), .B1(new_n524_), .B2(new_n523_), .ZN(new_n527_));
  OR2_X1    g455(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g456(.A(new_n343_), .B(new_n345_), .ZN(new_n529_));
  NAND2_X1  g457(.A1(new_n349_), .A2(G330), .ZN(new_n530_));
  XNOR2_X1  g458(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g459(.A(new_n531_), .ZN(new_n532_));
  NAND4_X1  g460(.A1(new_n521_), .A2(new_n528_), .A3(new_n365_), .A4(new_n532_), .ZN(new_n533_));
  INV_X1    g461(.A(new_n365_), .ZN(new_n534_));
  NAND2_X1  g462(.A1(new_n521_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g463(.A(new_n503_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g464(.A1(new_n521_), .A2(new_n372_), .ZN(new_n537_));
  INV_X1    g465(.A(new_n420_), .ZN(new_n538_));
  AOI22_X1  g466(.A1(new_n101_), .A2(new_n409_), .B1(new_n210_), .B2(new_n412_), .ZN(new_n539_));
  AOI21_X1  g467(.A(new_n538_), .B1(new_n539_), .B2(new_n415_), .ZN(new_n540_));
  NOR2_X1   g468(.A1(new_n376_), .A2(new_n192_), .ZN(new_n541_));
  AOI22_X1  g469(.A1(new_n380_), .A2(G150), .B1(new_n383_), .B2(G143), .ZN(new_n542_));
  OAI221_X1 g470(.A(new_n542_), .B1(new_n84_), .B2(new_n386_), .C1(new_n238_), .C2(new_n385_), .ZN(new_n543_));
  AOI211_X1 g471(.A(new_n541_), .B(new_n543_), .C1(G58), .C2(new_n388_), .ZN(new_n544_));
  NAND2_X1  g472(.A1(new_n390_), .A2(G77), .ZN(new_n545_));
  NAND2_X1  g473(.A1(new_n392_), .A2(G137), .ZN(new_n546_));
  NAND4_X1  g474(.A1(new_n544_), .A2(new_n113_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  NOR2_X1   g475(.A1(new_n395_), .A2(new_n284_), .ZN(RLL_wire_A_46));
  XNOR2_X1 RLL_XNOR_46 (.A(RLL_wire_A_46), .B(KEYINPUT46), .ZN(new_n548_) );
  AOI22_X1  g476(.A1(new_n380_), .A2(G303), .B1(new_n383_), .B2(G311), .ZN(new_n549_));
  INV_X1    g477(.A(G294), .ZN(new_n550_));
  OAI221_X1 g478(.A(new_n549_), .B1(new_n286_), .B2(new_n386_), .C1(new_n550_), .C2(new_n385_), .ZN(new_n551_));
  AOI211_X1 g479(.A(new_n548_), .B(new_n551_), .C1(G107), .C2(new_n401_), .ZN(new_n552_));
  NAND2_X1  g480(.A1(new_n390_), .A2(G97), .ZN(new_n553_));
  NAND2_X1  g481(.A1(new_n392_), .A2(G317), .ZN(new_n554_));
  NAND3_X1  g482(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OAI21_X1  g483(.A(new_n547_), .B1(new_n555_), .B2(new_n113_), .ZN(RLL_wire_A_47));
  XNOR2_X1 RLL_XNOR_47 (.A(RLL_wire_A_47), .B(KEYINPUT47), .ZN(new_n556_) );
  AOI21_X1  g484(.A(new_n540_), .B1(new_n556_), .B2(new_n408_), .ZN(new_n557_));
  OAI211_X1 g485(.A(new_n557_), .B(new_n422_), .C1(new_n423_), .C2(new_n513_), .ZN(new_n558_));
  NAND2_X1  g486(.A1(new_n537_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g487(.A1(new_n536_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g488(.A(new_n560_), .ZN(G387));
  NAND2_X1  g489(.A1(new_n532_), .A2(new_n365_), .ZN(new_n562_));
  NAND2_X1  g490(.A1(new_n531_), .A2(new_n534_), .ZN(new_n563_));
  NAND3_X1  g491(.A1(new_n562_), .A2(new_n353_), .A3(new_n563_), .ZN(new_n564_));
  NOR2_X1   g492(.A1(new_n376_), .A2(new_n210_), .ZN(new_n565_));
  AOI22_X1  g493(.A1(new_n380_), .A2(G50), .B1(new_n383_), .B2(G159), .ZN(new_n566_));
  OAI221_X1 g494(.A(new_n566_), .B1(new_n159_), .B2(new_n385_), .C1(new_n192_), .C2(new_n386_), .ZN(new_n567_));
  AOI211_X1 g495(.A(new_n565_), .B(new_n567_), .C1(G77), .C2(new_n388_), .ZN(new_n568_));
  NAND2_X1  g496(.A1(new_n392_), .A2(G150), .ZN(new_n569_));
  NAND4_X1  g497(.A1(new_n568_), .A2(new_n113_), .A3(new_n553_), .A4(new_n569_), .ZN(new_n570_));
  NOR2_X1   g498(.A1(new_n395_), .A2(new_n550_), .ZN(new_n571_));
  AOI22_X1  g499(.A1(new_n380_), .A2(G317), .B1(new_n383_), .B2(G322), .ZN(new_n572_));
  OAI221_X1 g500(.A(new_n572_), .B1(new_n278_), .B2(new_n386_), .C1(new_n398_), .C2(new_n385_), .ZN(RLL_wire_A_48));
  XOR2_X1 RLL_XOR_48 (.A(RLL_wire_A_48), .B(KEYINPUT48), .Z(new_n573_) );
  AOI211_X1 g501(.A(new_n571_), .B(new_n573_), .C1(G283), .C2(new_n401_), .ZN(RLL_wire_A_49));
  XOR2_X1 RLL_XOR_49 (.A(RLL_wire_A_49), .B(KEYINPUT49), .Z(new_n574_) );
  NAND2_X1  g502(.A1(new_n390_), .A2(G116), .ZN(new_n575_));
  NAND2_X1  g503(.A1(new_n392_), .A2(G326), .ZN(new_n576_));
  NAND3_X1  g504(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  OAI21_X1  g505(.A(new_n570_), .B1(new_n577_), .B2(new_n113_), .ZN(new_n578_));
  NAND2_X1  g506(.A1(G68), .A2(G77), .ZN(new_n579_));
  NOR2_X1   g507(.A1(new_n159_), .A2(G50), .ZN(RLL_wire_A_50));
  XNOR2_X1 RLL_XNOR_50 (.A(RLL_wire_A_50), .B(KEYINPUT50), .ZN(new_n580_) );
  NAND4_X1  g508(.A1(new_n355_), .A2(new_n265_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n581_));
  OAI211_X1 g509(.A(new_n409_), .B(new_n581_), .C1(new_n104_), .C2(new_n265_), .ZN(new_n582_));
  OAI221_X1 g510(.A(new_n582_), .B1(G107), .B2(new_n413_), .C1(new_n355_), .C2(new_n415_), .ZN(new_n583_));
  AOI22_X1  g511(.A1(new_n578_), .A2(new_n408_), .B1(new_n420_), .B2(new_n583_), .ZN(new_n584_));
  OR2_X1    g512(.A1(new_n343_), .A2(new_n423_), .ZN(new_n585_));
  NAND3_X1  g513(.A1(new_n584_), .A2(new_n422_), .A3(new_n585_), .ZN(new_n586_));
  OAI211_X1 g514(.A(new_n564_), .B(new_n586_), .C1(new_n371_), .C2(new_n531_), .ZN(G393));
  NOR2_X1   g515(.A1(new_n528_), .A2(new_n562_), .ZN(new_n588_));
  INV_X1    g516(.A(new_n527_), .ZN(new_n589_));
  AOI22_X1  g517(.A1(new_n532_), .A2(new_n365_), .B1(new_n525_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g518(.A(new_n353_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  AOI22_X1  g519(.A1(new_n111_), .A2(new_n409_), .B1(new_n89_), .B2(new_n412_), .ZN(new_n592_));
  AOI21_X1  g520(.A(new_n538_), .B1(new_n592_), .B2(new_n415_), .ZN(new_n593_));
  NOR2_X1   g521(.A1(new_n376_), .A2(new_n74_), .ZN(new_n594_));
  AOI22_X1  g522(.A1(new_n380_), .A2(G159), .B1(new_n383_), .B2(G150), .ZN(RLL_wire_A_51));
  XOR2_X1 RLL_XOR_51 (.A(RLL_wire_A_51), .B(KEYINPUT51), .Z(new_n595_) );
  OAI221_X1 g523(.A(new_n595_), .B1(new_n84_), .B2(new_n385_), .C1(new_n159_), .C2(new_n386_), .ZN(new_n596_));
  AOI211_X1 g524(.A(new_n594_), .B(new_n596_), .C1(G68), .C2(new_n388_), .ZN(new_n597_));
  NAND2_X1  g525(.A1(new_n392_), .A2(G143), .ZN(new_n598_));
  NAND4_X1  g526(.A1(new_n597_), .A2(new_n113_), .A3(new_n451_), .A4(new_n598_), .ZN(new_n599_));
  NOR2_X1   g527(.A1(new_n395_), .A2(new_n286_), .ZN(new_n600_));
  AOI22_X1  g528(.A1(new_n380_), .A2(G311), .B1(new_n383_), .B2(G317), .ZN(RLL_wire_A_52));
  XOR2_X1 RLL_XOR_52 (.A(RLL_wire_A_52), .B(KEYINPUT52), .Z(new_n601_) );
  OAI221_X1 g529(.A(new_n601_), .B1(new_n550_), .B2(new_n386_), .C1(new_n278_), .C2(new_n385_), .ZN(new_n602_));
  AOI211_X1 g530(.A(new_n600_), .B(new_n602_), .C1(G116), .C2(new_n401_), .ZN(new_n603_));
  NAND2_X1  g531(.A1(new_n392_), .A2(G322), .ZN(new_n604_));
  NAND3_X1  g532(.A1(new_n603_), .A2(new_n391_), .A3(new_n604_), .ZN(new_n605_));
  OAI21_X1  g533(.A(new_n599_), .B1(new_n605_), .B2(new_n113_), .ZN(new_n606_));
  AOI21_X1  g534(.A(new_n593_), .B1(new_n606_), .B2(new_n408_), .ZN(new_n607_));
  OAI211_X1 g535(.A(new_n607_), .B(new_n422_), .C1(new_n423_), .C2(new_n507_), .ZN(new_n608_));
  INV_X1    g536(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g537(.A(new_n609_), .B1(new_n528_), .B2(new_n372_), .ZN(new_n610_));
  NAND2_X1  g538(.A1(new_n591_), .A2(new_n610_), .ZN(G390));
  NAND4_X1  g539(.A1(new_n336_), .A2(new_n470_), .A3(new_n340_), .A4(new_n431_), .ZN(new_n612_));
  NAND2_X1  g540(.A1(new_n470_), .A2(new_n483_), .ZN(new_n613_));
  NAND3_X1  g541(.A1(new_n612_), .A2(new_n490_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g542(.A1(new_n614_), .A2(new_n488_), .ZN(new_n615_));
  NAND4_X1  g543(.A1(new_n612_), .A2(new_n482_), .A3(new_n490_), .A4(new_n613_), .ZN(new_n616_));
  NAND2_X1  g544(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g545(.A1(new_n364_), .A2(G330), .A3(new_n431_), .A4(new_n470_), .ZN(new_n618_));
  NAND2_X1  g546(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g547(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g548(.A1(new_n615_), .A2(new_n620_), .A3(new_n616_), .ZN(new_n621_));
  NAND2_X1  g549(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g550(.A1(new_n336_), .A2(new_n340_), .A3(new_n431_), .ZN(new_n623_));
  INV_X1    g551(.A(new_n483_), .ZN(new_n624_));
  NAND2_X1  g552(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g553(.A1(new_n625_), .A2(new_n486_), .ZN(new_n626_));
  AOI211_X1 g554(.A(new_n351_), .B(new_n432_), .C1(new_n359_), .C2(new_n363_), .ZN(new_n627_));
  NAND3_X1  g555(.A1(new_n623_), .A2(new_n470_), .A3(new_n624_), .ZN(new_n628_));
  NAND3_X1  g556(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g557(.A1(new_n364_), .A2(G330), .A3(new_n431_), .ZN(new_n630_));
  AND3_X1   g558(.A1(new_n623_), .A2(new_n470_), .A3(new_n624_), .ZN(new_n631_));
  AOI21_X1  g559(.A(new_n470_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n632_));
  OAI21_X1  g560(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g561(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g562(.A(new_n330_), .B(new_n493_), .C1(new_n497_), .C2(new_n351_), .ZN(new_n635_));
  INV_X1    g563(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g564(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g565(.A1(new_n622_), .A2(new_n637_), .ZN(new_n638_));
  AOI22_X1  g566(.A1(new_n621_), .A2(new_n619_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n639_));
  OAI21_X1  g567(.A(new_n353_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g568(.A1(new_n395_), .A2(new_n442_), .ZN(RLL_wire_A_53));
  XOR2_X1 RLL_XOR_53 (.A(RLL_wire_A_53), .B(KEYINPUT53), .Z(new_n641_) );
  AOI22_X1  g569(.A1(new_n380_), .A2(G132), .B1(new_n383_), .B2(G128), .ZN(new_n642_));
  INV_X1    g570(.A(G137), .ZN(new_n643_));
  INV_X1    g571(.A(G143), .ZN(RLL_wire_A_54));
  XOR2_X1 RLL_XOR_54 (.A(RLL_wire_A_54), .B(KEYINPUT54), .Z(new_n644_) );
  OAI221_X1 g572(.A(new_n642_), .B1(new_n643_), .B2(new_n385_), .C1(new_n644_), .C2(new_n386_), .ZN(new_n645_));
  AOI211_X1 g573(.A(new_n641_), .B(new_n645_), .C1(G159), .C2(new_n401_), .ZN(new_n646_));
  NAND2_X1  g574(.A1(new_n390_), .A2(G50), .ZN(new_n647_));
  NAND2_X1  g575(.A1(new_n392_), .A2(G125), .ZN(new_n648_));
  NAND4_X1  g576(.A1(new_n646_), .A2(new_n113_), .A3(new_n647_), .A4(new_n648_), .ZN(new_n649_));
  AOI22_X1  g577(.A1(new_n380_), .A2(G116), .B1(new_n383_), .B2(G283), .ZN(new_n650_));
  OAI221_X1 g578(.A(new_n650_), .B1(new_n89_), .B2(new_n386_), .C1(new_n137_), .C2(new_n385_), .ZN(new_n651_));
  AOI211_X1 g579(.A(new_n594_), .B(new_n651_), .C1(G87), .C2(new_n388_), .ZN(new_n652_));
  NAND2_X1  g580(.A1(new_n392_), .A2(G294), .ZN(new_n653_));
  NAND3_X1  g581(.A1(new_n652_), .A2(new_n445_), .A3(new_n653_), .ZN(new_n654_));
  OAI21_X1  g582(.A(new_n649_), .B1(new_n654_), .B2(new_n113_), .ZN(new_n655_));
  AOI22_X1  g583(.A1(new_n655_), .A2(new_n408_), .B1(new_n159_), .B2(new_n455_), .ZN(new_n656_));
  NAND2_X1  g584(.A1(new_n488_), .A2(new_n417_), .ZN(new_n657_));
  NAND3_X1  g585(.A1(new_n656_), .A2(new_n422_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g586(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g587(.A(new_n659_), .B1(new_n622_), .B2(new_n372_), .ZN(new_n660_));
  NAND2_X1  g588(.A1(new_n640_), .A2(new_n660_), .ZN(G378));
  AND3_X1   g589(.A1(new_n470_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n662_));
  AND4_X1   g590(.A1(new_n336_), .A2(new_n340_), .A3(new_n431_), .A4(new_n482_), .ZN(new_n663_));
  AOI21_X1  g591(.A(new_n662_), .B1(new_n663_), .B2(new_n470_), .ZN(new_n664_));
  INV_X1    g592(.A(new_n491_), .ZN(new_n665_));
  NAND2_X1  g593(.A1(new_n165_), .A2(new_n472_), .ZN(RLL_wire_A_55));
  XOR2_X1 RLL_XOR_55 (.A(RLL_wire_A_55), .B(KEYINPUT55), .Z(new_n666_) );
  XNOR2_X1  g594(.A(new_n185_), .B(new_n666_), .ZN(RLL_wire_A_56));
  XNOR2_X1 RLL_XNOR_56 (.A(RLL_wire_A_56), .B(KEYINPUT56), .ZN(new_n667_) );
  INV_X1    g595(.A(new_n667_), .ZN(new_n668_));
  NAND4_X1  g596(.A1(new_n664_), .A2(new_n665_), .A3(new_n465_), .A4(new_n668_), .ZN(new_n669_));
  NOR2_X1   g597(.A1(new_n496_), .A2(new_n351_), .ZN(new_n670_));
  OAI21_X1  g598(.A(new_n667_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n671_));
  AND3_X1   g599(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g600(.A(new_n670_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g601(.A(new_n635_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g602(.A(new_n634_), .B(new_n636_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n675_));
  INV_X1    g603(.A(new_n622_), .ZN(new_n676_));
  OAI21_X1  g604(.A(new_n674_), .B1(new_n675_), .B2(new_n676_), .ZN(RLL_wire_A_57));
  XOR2_X1 RLL_XOR_57 (.A(RLL_wire_A_57), .B(KEYINPUT57), .Z(new_n677_) );
  NAND2_X1  g605(.A1(new_n677_), .A2(new_n353_), .ZN(new_n678_));
  INV_X1    g606(.A(new_n670_), .ZN(new_n679_));
  INV_X1    g607(.A(new_n487_), .ZN(new_n680_));
  AOI21_X1  g608(.A(new_n668_), .B1(new_n680_), .B2(new_n665_), .ZN(new_n681_));
  NOR3_X1   g609(.A1(new_n487_), .A2(new_n491_), .A3(new_n667_), .ZN(new_n682_));
  OAI21_X1  g610(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g611(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n684_));
  NAND2_X1  g612(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g613(.A1(new_n685_), .A2(new_n372_), .ZN(new_n686_));
  AOI22_X1  g614(.A1(new_n380_), .A2(G107), .B1(new_n383_), .B2(G116), .ZN(new_n687_));
  OAI221_X1 g615(.A(new_n687_), .B1(new_n210_), .B2(new_n386_), .C1(new_n89_), .C2(new_n385_), .ZN(new_n688_));
  AOI211_X1 g616(.A(new_n541_), .B(new_n688_), .C1(G77), .C2(new_n388_), .ZN(new_n689_));
  NOR2_X1   g617(.A1(new_n113_), .A2(G41), .ZN(new_n690_));
  NAND2_X1  g618(.A1(new_n390_), .A2(G58), .ZN(new_n691_));
  NAND2_X1  g619(.A1(new_n392_), .A2(G283), .ZN(new_n692_));
  NAND4_X1  g620(.A1(new_n689_), .A2(new_n690_), .A3(new_n691_), .A4(new_n692_), .ZN(RLL_wire_A_58));
  XNOR2_X1 RLL_XNOR_58 (.A(RLL_wire_A_58), .B(KEYINPUT58), .ZN(new_n693_) );
  NOR2_X1   g621(.A1(new_n395_), .A2(new_n644_), .ZN(new_n694_));
  AOI22_X1  g622(.A1(new_n380_), .A2(G128), .B1(new_n383_), .B2(G125), .ZN(new_n695_));
  INV_X1    g623(.A(G132), .ZN(new_n696_));
  OAI221_X1 g624(.A(new_n695_), .B1(new_n696_), .B2(new_n385_), .C1(new_n643_), .C2(new_n386_), .ZN(new_n697_));
  AOI211_X1 g625(.A(new_n694_), .B(new_n697_), .C1(G150), .C2(new_n401_), .ZN(RLL_wire_A_59));
  XNOR2_X1 RLL_XNOR_59 (.A(RLL_wire_A_59), .B(KEYINPUT59), .ZN(new_n698_) );
  NOR2_X1   g626(.A1(G33), .A2(G41), .ZN(new_n699_));
  NAND2_X1  g627(.A1(new_n390_), .A2(G159), .ZN(new_n700_));
  NAND2_X1  g628(.A1(new_n392_), .A2(G124), .ZN(new_n701_));
  NAND4_X1  g629(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .A4(new_n701_), .ZN(new_n702_));
  OR3_X1    g630(.A1(new_n690_), .A2(G50), .A3(new_n699_), .ZN(new_n703_));
  NAND3_X1  g631(.A1(new_n693_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  AOI22_X1  g632(.A1(new_n704_), .A2(new_n408_), .B1(new_n84_), .B2(new_n455_), .ZN(new_n705_));
  OAI211_X1 g633(.A(new_n705_), .B(new_n422_), .C1(new_n668_), .C2(new_n418_), .ZN(new_n706_));
  NAND2_X1  g634(.A1(new_n686_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g635(.A(new_n707_), .ZN(new_n708_));
  NAND2_X1  g636(.A1(new_n678_), .A2(new_n708_), .ZN(G375));
  INV_X1    g637(.A(new_n637_), .ZN(new_n710_));
  NOR2_X1   g638(.A1(new_n634_), .A2(new_n636_), .ZN(new_n711_));
  NOR3_X1   g639(.A1(new_n710_), .A2(new_n711_), .A3(new_n503_), .ZN(new_n712_));
  NAND2_X1  g640(.A1(new_n634_), .A2(new_n372_), .ZN(new_n713_));
  NOR2_X1   g641(.A1(new_n395_), .A2(new_n238_), .ZN(new_n714_));
  AOI22_X1  g642(.A1(new_n380_), .A2(G137), .B1(new_n383_), .B2(G132), .ZN(new_n715_));
  OAI221_X1 g643(.A(new_n715_), .B1(new_n644_), .B2(new_n385_), .C1(new_n442_), .C2(new_n386_), .ZN(new_n716_));
  AOI211_X1 g644(.A(new_n714_), .B(new_n716_), .C1(G50), .C2(new_n401_), .ZN(new_n717_));
  NAND2_X1  g645(.A1(new_n392_), .A2(G128), .ZN(new_n718_));
  NAND4_X1  g646(.A1(new_n717_), .A2(new_n113_), .A3(new_n691_), .A4(new_n718_), .ZN(new_n719_));
  AOI22_X1  g647(.A1(new_n380_), .A2(G283), .B1(new_n383_), .B2(G294), .ZN(new_n720_));
  OAI221_X1 g648(.A(new_n720_), .B1(new_n137_), .B2(new_n386_), .C1(new_n284_), .C2(new_n385_), .ZN(new_n721_));
  AOI211_X1 g649(.A(new_n565_), .B(new_n721_), .C1(G97), .C2(new_n388_), .ZN(new_n722_));
  NAND2_X1  g650(.A1(new_n392_), .A2(G303), .ZN(new_n723_));
  NAND3_X1  g651(.A1(new_n722_), .A2(new_n545_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g652(.A(new_n719_), .B1(new_n724_), .B2(new_n113_), .ZN(new_n725_));
  AOI22_X1  g653(.A1(new_n725_), .A2(new_n408_), .B1(new_n192_), .B2(new_n455_), .ZN(new_n726_));
  NAND2_X1  g654(.A1(new_n486_), .A2(new_n417_), .ZN(new_n727_));
  NAND3_X1  g655(.A1(new_n726_), .A2(new_n422_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g656(.A1(new_n713_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g657(.A1(new_n712_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g658(.A(new_n730_), .ZN(G381));
  NOR4_X1   g659(.A1(G375), .A2(G384), .A3(G381), .A4(G378), .ZN(new_n732_));
  NOR4_X1   g660(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n733_));
  NAND2_X1  g661(.A1(new_n732_), .A2(new_n733_), .ZN(G407));
  INV_X1    g662(.A(G343), .ZN(new_n735_));
  NAND2_X1  g663(.A1(new_n735_), .A2(G213), .ZN(new_n736_));
  OR3_X1    g664(.A1(G375), .A2(G378), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g665(.A1(G407), .A2(G213), .A3(new_n737_), .ZN(G409));
  INV_X1    g666(.A(new_n660_), .ZN(new_n739_));
  XNOR2_X1  g667(.A(new_n622_), .B(new_n637_), .ZN(new_n740_));
  AOI21_X1  g668(.A(new_n739_), .B1(new_n740_), .B2(new_n353_), .ZN(new_n741_));
  NAND4_X1  g669(.A1(new_n685_), .A2(new_n622_), .A3(new_n634_), .A4(new_n636_), .ZN(new_n742_));
  AOI21_X1  g670(.A(new_n503_), .B1(new_n742_), .B2(new_n674_), .ZN(new_n743_));
  OAI211_X1 g671(.A(new_n741_), .B(new_n736_), .C1(new_n743_), .C2(new_n707_), .ZN(new_n744_));
  NAND4_X1  g672(.A1(new_n678_), .A2(G378), .A3(new_n708_), .A4(new_n736_), .ZN(new_n745_));
  NAND2_X1  g673(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g674(.A(new_n711_), .ZN(RLL_wire_A_60));
  XNOR2_X1 RLL_XNOR_60 (.A(RLL_wire_A_60), .B(KEYINPUT60), .ZN(new_n747_) );
  NAND3_X1  g675(.A1(new_n747_), .A2(new_n353_), .A3(new_n637_), .ZN(new_n748_));
  INV_X1    g676(.A(new_n729_), .ZN(new_n749_));
  AND3_X1   g677(.A1(new_n748_), .A2(G384), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g678(.A(G384), .B1(new_n748_), .B2(new_n749_), .ZN(new_n751_));
  NOR2_X1   g679(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g680(.A1(new_n735_), .A2(G213), .A3(G2897), .ZN(new_n753_));
  NOR2_X1   g681(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g682(.A1(new_n746_), .A2(new_n754_), .ZN(RLL_wire_A_61));
  XOR2_X1 RLL_XOR_61 (.A(RLL_wire_A_61), .B(KEYINPUT61), .Z(new_n755_) );
  INV_X1    g683(.A(new_n751_), .ZN(new_n756_));
  NAND3_X1  g684(.A1(new_n748_), .A2(G384), .A3(new_n749_), .ZN(new_n757_));
  NAND3_X1  g685(.A1(new_n756_), .A2(new_n753_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g686(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g687(.A1(new_n746_), .A2(new_n759_), .ZN(RLL_wire_A_62));
  XOR2_X1 RLL_XOR_62 (.A(RLL_wire_A_62), .B(KEYINPUT62), .Z(new_n760_) );
  INV_X1    g688(.A(new_n752_), .ZN(new_n761_));
  NAND4_X1  g689(.A1(new_n761_), .A2(new_n744_), .A3(new_n745_), .A4(new_n753_), .ZN(new_n762_));
  NOR3_X1   g690(.A1(new_n750_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n763_));
  NAND3_X1  g691(.A1(new_n744_), .A2(new_n745_), .A3(new_n763_), .ZN(new_n764_));
  NAND4_X1  g692(.A1(new_n755_), .A2(new_n760_), .A3(new_n762_), .A4(new_n764_), .ZN(new_n765_));
  NAND2_X1  g693(.A1(new_n560_), .A2(G390), .ZN(new_n766_));
  OAI211_X1 g694(.A(new_n591_), .B(new_n610_), .C1(new_n536_), .C2(new_n559_), .ZN(new_n767_));
  NAND2_X1  g695(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g696(.A(G393), .B(new_n425_), .ZN(new_n769_));
  INV_X1    g697(.A(new_n769_), .ZN(new_n770_));
  NAND2_X1  g698(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g699(.A1(new_n766_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n772_));
  NAND2_X1  g700(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g701(.A1(new_n765_), .A2(new_n773_), .ZN(new_n774_));
  AND3_X1   g702(.A1(new_n744_), .A2(new_n745_), .A3(new_n763_), .ZN(new_n775_));
  AOI21_X1  g703(.A(new_n758_), .B1(new_n744_), .B2(new_n745_), .ZN(RLL_wire_A_63));
  XNOR2_X1 RLL_XNOR_63 (.A(RLL_wire_A_63), .B(KEYINPUT63), .ZN(new_n776_) );
  NOR2_X1   g704(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g705(.A(new_n772_), .ZN(new_n778_));
  AOI21_X1  g706(.A(new_n769_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n779_));
  NOR2_X1   g707(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND4_X1  g708(.A1(new_n777_), .A2(new_n780_), .A3(new_n762_), .A4(new_n755_), .ZN(new_n781_));
  NAND2_X1  g709(.A1(new_n774_), .A2(new_n781_), .ZN(G405));
  NAND3_X1  g710(.A1(new_n678_), .A2(G378), .A3(new_n708_), .ZN(new_n783_));
  INV_X1    g711(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g712(.A(G378), .B1(new_n678_), .B2(new_n708_), .ZN(new_n785_));
  OAI21_X1  g713(.A(new_n752_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g714(.A(new_n785_), .ZN(new_n787_));
  NAND3_X1  g715(.A1(new_n787_), .A2(new_n761_), .A3(new_n783_), .ZN(new_n788_));
  NAND2_X1  g716(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g717(.A(new_n789_), .B(new_n773_), .ZN(G402));

endmodule
