

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U324 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U325 ( .A(KEYINPUT41), .B(n579), .Z(n551) );
  XNOR2_X1 U326 ( .A(KEYINPUT106), .B(KEYINPUT37), .ZN(n482) );
  XNOR2_X1 U327 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n442) );
  NOR2_X1 U328 ( .A1(n567), .A2(n566), .ZN(n292) );
  XOR2_X1 U329 ( .A(n423), .B(n304), .Z(n293) );
  XOR2_X1 U330 ( .A(n333), .B(KEYINPUT74), .Z(n294) );
  XNOR2_X1 U331 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n373) );
  XNOR2_X1 U332 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U333 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U334 ( .A(n422), .B(n313), .ZN(n317) );
  XNOR2_X1 U335 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n371) );
  INV_X1 U336 ( .A(KEYINPUT88), .ZN(n433) );
  XNOR2_X1 U337 ( .A(n372), .B(n371), .ZN(n379) );
  XNOR2_X1 U338 ( .A(n436), .B(n435), .ZN(n437) );
  NOR2_X1 U339 ( .A1(n421), .A2(n520), .ZN(n573) );
  XNOR2_X1 U340 ( .A(n305), .B(n293), .ZN(n306) );
  XNOR2_X1 U341 ( .A(n443), .B(n442), .ZN(n568) );
  XNOR2_X1 U342 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U343 ( .A(n483), .B(n482), .ZN(n518) );
  XNOR2_X1 U344 ( .A(n329), .B(n328), .ZN(n579) );
  XOR2_X1 U345 ( .A(KEYINPUT28), .B(n476), .Z(n527) );
  XNOR2_X1 U346 ( .A(n488), .B(G183GAT), .ZN(n489) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n486) );
  XNOR2_X1 U348 ( .A(n490), .B(n489), .ZN(G1350GAT) );
  XNOR2_X1 U349 ( .A(n487), .B(n486), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n296) );
  XNOR2_X1 U351 ( .A(G92GAT), .B(KEYINPUT73), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n309) );
  XOR2_X1 U353 ( .A(G29GAT), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U354 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n333) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n294), .B(n299), .ZN(n307) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(G85GAT), .ZN(n328) );
  XOR2_X1 U359 ( .A(G36GAT), .B(G190GAT), .Z(n388) );
  XNOR2_X1 U360 ( .A(n328), .B(n388), .ZN(n301) );
  XNOR2_X1 U361 ( .A(G218GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U362 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XOR2_X1 U364 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n303) );
  XNOR2_X1 U365 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n302) );
  XNOR2_X1 U366 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U367 ( .A(n309), .B(n308), .Z(n559) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n310), .B(G148GAT), .ZN(n422) );
  NAND2_X1 U370 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  INV_X1 U371 ( .A(KEYINPUT32), .ZN(n311) );
  XOR2_X1 U372 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n315) );
  XNOR2_X1 U373 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n322) );
  XOR2_X1 U376 ( .A(G64GAT), .B(G92GAT), .Z(n319) );
  XNOR2_X1 U377 ( .A(G176GAT), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n387) );
  XNOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n320), .B(KEYINPUT13), .ZN(n361) );
  XOR2_X1 U381 ( .A(n387), .B(n361), .Z(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U383 ( .A(G120GAT), .B(G71GAT), .Z(n450) );
  NAND2_X1 U384 ( .A1(n323), .A2(n450), .ZN(n327) );
  INV_X1 U385 ( .A(n450), .ZN(n325) );
  INV_X1 U386 ( .A(n323), .ZN(n324) );
  NAND2_X1 U387 ( .A1(n325), .A2(n324), .ZN(n326) );
  AND2_X1 U388 ( .A1(n327), .A2(n326), .ZN(n329) );
  XOR2_X1 U389 ( .A(G197GAT), .B(G113GAT), .Z(n331) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(G36GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U392 ( .A(G15GAT), .B(G1GAT), .Z(n363) );
  XOR2_X1 U393 ( .A(n332), .B(n363), .Z(n338) );
  XOR2_X1 U394 ( .A(n333), .B(KEYINPUT67), .Z(n335) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U397 ( .A(G169GAT), .B(G8GAT), .Z(n392) );
  XNOR2_X1 U398 ( .A(n336), .B(n392), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n346) );
  XOR2_X1 U400 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n340) );
  XNOR2_X1 U401 ( .A(G141GAT), .B(G22GAT), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n342) );
  XNOR2_X1 U404 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U406 ( .A(n344), .B(n343), .Z(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n576) );
  NOR2_X1 U408 ( .A1(n551), .A2(n576), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(KEYINPUT46), .ZN(n368) );
  XOR2_X1 U410 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n349) );
  XNOR2_X1 U411 ( .A(KEYINPUT81), .B(KEYINPUT14), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n367) );
  XOR2_X1 U413 ( .A(G211GAT), .B(G71GAT), .Z(n351) );
  XNOR2_X1 U414 ( .A(G183GAT), .B(G127GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U416 ( .A(KEYINPUT80), .B(G64GAT), .Z(n353) );
  XNOR2_X1 U417 ( .A(G8GAT), .B(G78GAT), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U419 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U420 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n357) );
  NAND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U423 ( .A(KEYINPUT79), .B(n358), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U425 ( .A(n362), .B(n361), .Z(n365) );
  XOR2_X1 U426 ( .A(G22GAT), .B(G155GAT), .Z(n429) );
  XNOR2_X1 U427 ( .A(n363), .B(n429), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n556) );
  NOR2_X1 U430 ( .A1(n368), .A2(n556), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n369), .B(KEYINPUT111), .ZN(n370) );
  NOR2_X1 U432 ( .A1(n559), .A2(n370), .ZN(n372) );
  INV_X1 U433 ( .A(n556), .ZN(n582) );
  INV_X1 U434 ( .A(n559), .ZN(n567) );
  XNOR2_X1 U435 ( .A(KEYINPUT36), .B(n567), .ZN(n585) );
  NOR2_X1 U436 ( .A1(n582), .A2(n585), .ZN(n374) );
  NAND2_X1 U437 ( .A1(n375), .A2(n579), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n376), .B(KEYINPUT113), .ZN(n377) );
  NAND2_X1 U439 ( .A1(n377), .A2(n576), .ZN(n378) );
  NAND2_X1 U440 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n380), .B(KEYINPUT48), .ZN(n543) );
  XOR2_X1 U442 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n382) );
  XNOR2_X1 U443 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U445 ( .A(KEYINPUT86), .B(n383), .Z(n457) );
  XOR2_X1 U446 ( .A(KEYINPUT21), .B(G218GAT), .Z(n385) );
  XNOR2_X1 U447 ( .A(KEYINPUT90), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U449 ( .A(G197GAT), .B(n386), .Z(n439) );
  XNOR2_X1 U450 ( .A(n457), .B(n439), .ZN(n396) );
  XOR2_X1 U451 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U454 ( .A(n391), .B(KEYINPUT97), .Z(n394) );
  XNOR2_X1 U455 ( .A(n392), .B(KEYINPUT98), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n522) );
  NAND2_X1 U458 ( .A1(n543), .A2(n522), .ZN(n398) );
  XOR2_X1 U459 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n421) );
  XOR2_X1 U461 ( .A(G57GAT), .B(G155GAT), .Z(n400) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(G148GAT), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U464 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n402) );
  XNOR2_X1 U465 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U467 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U468 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n406) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U471 ( .A(KEYINPUT5), .B(n407), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n415) );
  XOR2_X1 U473 ( .A(G85GAT), .B(G162GAT), .Z(n413) );
  XOR2_X1 U474 ( .A(KEYINPUT91), .B(KEYINPUT3), .Z(n411) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n432) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(n432), .ZN(n412) );
  XNOR2_X1 U478 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U479 ( .A(n415), .B(n414), .Z(n420) );
  XOR2_X1 U480 ( .A(KEYINPUT0), .B(G134GAT), .Z(n417) );
  XNOR2_X1 U481 ( .A(KEYINPUT83), .B(G127GAT), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U483 ( .A(G113GAT), .B(n418), .Z(n458) );
  XNOR2_X1 U484 ( .A(n458), .B(G120GAT), .ZN(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n520) );
  XOR2_X1 U486 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n438) );
  XOR2_X1 U489 ( .A(G204GAT), .B(KEYINPUT89), .Z(n427) );
  XNOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U492 ( .A(n428), .B(KEYINPUT92), .Z(n431) );
  XNOR2_X1 U493 ( .A(n429), .B(KEYINPUT22), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n432), .B(KEYINPUT93), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n441) );
  INV_X1 U497 ( .A(n439), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n476) );
  NAND2_X1 U499 ( .A1(n573), .A2(n476), .ZN(n443) );
  XOR2_X1 U500 ( .A(KEYINPUT87), .B(G99GAT), .Z(n445) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(G190GAT), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U503 ( .A(KEYINPUT84), .B(G176GAT), .Z(n447) );
  XNOR2_X1 U504 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U506 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U507 ( .A(n450), .B(KEYINPUT85), .Z(n452) );
  NAND2_X1 U508 ( .A1(G227GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U510 ( .A(G169GAT), .B(n453), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(n460) );
  INV_X1 U513 ( .A(n458), .ZN(n459) );
  XNOR2_X2 U514 ( .A(n460), .B(n459), .ZN(n565) );
  NAND2_X1 U515 ( .A1(n568), .A2(n565), .ZN(n562) );
  XNOR2_X1 U516 ( .A(n551), .B(KEYINPUT108), .ZN(n535) );
  NOR2_X1 U517 ( .A1(n562), .A2(n535), .ZN(n464) );
  XNOR2_X1 U518 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n462) );
  XNOR2_X1 U519 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  NOR2_X1 U522 ( .A1(n565), .A2(n476), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT26), .B(n465), .Z(n466) );
  XNOR2_X1 U524 ( .A(KEYINPUT101), .B(n466), .ZN(n574) );
  XNOR2_X1 U525 ( .A(n522), .B(KEYINPUT27), .ZN(n475) );
  NAND2_X1 U526 ( .A1(n574), .A2(n475), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n522), .A2(n565), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n467), .A2(n476), .ZN(n468) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT102), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(KEYINPUT103), .B(n472), .ZN(n473) );
  NOR2_X1 U533 ( .A1(n520), .A2(n473), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT104), .ZN(n480) );
  NAND2_X1 U535 ( .A1(n520), .A2(n475), .ZN(n545) );
  NOR2_X1 U536 ( .A1(n545), .A2(n527), .ZN(n530) );
  XNOR2_X1 U537 ( .A(KEYINPUT99), .B(n530), .ZN(n477) );
  NOR2_X1 U538 ( .A1(n565), .A2(n477), .ZN(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT100), .B(n478), .ZN(n479) );
  NOR2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n494) );
  NOR2_X1 U541 ( .A1(n585), .A2(n494), .ZN(n481) );
  NAND2_X1 U542 ( .A1(n582), .A2(n481), .ZN(n483) );
  INV_X1 U543 ( .A(n576), .ZN(n546) );
  AND2_X1 U544 ( .A1(n546), .A2(n579), .ZN(n495) );
  NAND2_X1 U545 ( .A1(n518), .A2(n495), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(KEYINPUT38), .ZN(n485) );
  XNOR2_X1 U547 ( .A(KEYINPUT107), .B(n485), .ZN(n507) );
  NAND2_X1 U548 ( .A1(n507), .A2(n565), .ZN(n487) );
  NOR2_X1 U549 ( .A1(n582), .A2(n562), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n488) );
  NAND2_X1 U551 ( .A1(n556), .A2(n567), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(KEYINPUT82), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT16), .ZN(n493) );
  NOR2_X1 U554 ( .A1(n494), .A2(n493), .ZN(n509) );
  AND2_X1 U555 ( .A1(n495), .A2(n509), .ZN(n501) );
  NAND2_X1 U556 ( .A1(n501), .A2(n520), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(KEYINPUT34), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(n497), .ZN(G1324GAT) );
  NAND2_X1 U559 ( .A1(n501), .A2(n522), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U562 ( .A1(n501), .A2(n565), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  XOR2_X1 U564 ( .A(G22GAT), .B(KEYINPUT105), .Z(n503) );
  NAND2_X1 U565 ( .A1(n501), .A2(n527), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1327GAT) );
  NAND2_X1 U567 ( .A1(n520), .A2(n507), .ZN(n505) );
  XOR2_X1 U568 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NAND2_X1 U570 ( .A1(n507), .A2(n522), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n507), .A2(n527), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U574 ( .A1(n546), .A2(n535), .ZN(n519) );
  AND2_X1 U575 ( .A1(n519), .A2(n509), .ZN(n515) );
  NAND2_X1 U576 ( .A1(n520), .A2(n515), .ZN(n510) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n510), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n522), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT109), .Z(n514) );
  NAND2_X1 U582 ( .A1(n515), .A2(n565), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U585 ( .A1(n515), .A2(n527), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  AND2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n526) );
  NAND2_X1 U588 ( .A1(n526), .A2(n520), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n521), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n522), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n565), .A2(n526), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n524), .B(KEYINPUT110), .ZN(n525) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n533) );
  AND2_X1 U599 ( .A1(n543), .A2(n530), .ZN(n531) );
  NAND2_X1 U600 ( .A1(n565), .A2(n531), .ZN(n534) );
  INV_X1 U601 ( .A(n534), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n546), .A2(n540), .ZN(n532) );
  XNOR2_X1 U603 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  NOR2_X1 U604 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n556), .A2(n540), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U611 ( .A1(n540), .A2(n559), .ZN(n541) );
  XNOR2_X1 U612 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n543), .A2(n574), .ZN(n544) );
  NOR2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n560), .A2(n546), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n549) );
  XNOR2_X1 U618 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n548) );
  XNOR2_X1 U619 ( .A(n549), .B(n548), .ZN(n555) );
  INV_X1 U620 ( .A(n560), .ZN(n550) );
  NOR2_X1 U621 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n552) );
  XNOR2_X1 U623 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U624 ( .A(n555), .B(n554), .Z(G1345GAT) );
  NAND2_X1 U625 ( .A1(n556), .A2(n560), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n557), .B(KEYINPUT118), .ZN(n558) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n558), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n576), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  INV_X1 U633 ( .A(n565), .ZN(n566) );
  AND2_X1 U634 ( .A1(n568), .A2(n292), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT58), .B(n569), .Z(n570) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(n575), .Z(n584) );
  NOR2_X1 U642 ( .A1(n576), .A2(n584), .ZN(n577) );
  XOR2_X1 U643 ( .A(n578), .B(n577), .Z(G1352GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n584), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

