//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n207), .A3(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n215), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n207), .A2(G1), .ZN(new_n254));
  INV_X1    g0054(.A(G50), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n253), .A2(new_n256), .B1(new_n255), .B2(new_n250), .ZN(new_n257));
  NOR3_X1   g0057(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n258), .A2(new_n207), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n264));
  OAI21_X1  g0064(.A(G58), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT8), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G58), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n270), .B(G58), .C1(new_n263), .C2(new_n264), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n266), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n262), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n252), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n257), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n273), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n288), .A2(KEYINPUT69), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT69), .B1(new_n288), .B2(new_n289), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n279), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n288), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G222), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n299), .A2(new_n300), .B1(new_n221), .B2(new_n293), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n278), .B1(new_n292), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G41), .ZN(new_n303));
  INV_X1    g0103(.A(G45), .ZN(new_n304));
  AOI21_X1  g0104(.A(G1), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n278), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G274), .ZN(new_n307));
  INV_X1    g0107(.A(new_n215), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G41), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n306), .A2(G226), .B1(new_n310), .B2(new_n305), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n277), .B1(new_n313), .B2(G169), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(new_n277), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(KEYINPUT9), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(KEYINPUT9), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(G200), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n302), .A2(G190), .A3(new_n311), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT10), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT10), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n320), .A2(new_n325), .A3(new_n321), .A4(new_n322), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n316), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n249), .A2(G1), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G20), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n272), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n254), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n271), .A2(new_n269), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT70), .B(KEYINPUT8), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n270), .B1(new_n334), .B2(G58), .ZN(new_n335));
  OAI211_X1 g0135(.A(KEYINPUT76), .B(new_n332), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n253), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT76), .B1(new_n272), .B2(new_n332), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G58), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n219), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G58), .A2(G68), .ZN(new_n342));
  OAI21_X1  g0142(.A(G20), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n259), .A2(G159), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n286), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n281), .A2(new_n282), .A3(new_n280), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT67), .B1(new_n285), .B2(new_n286), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n207), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n346), .B1(new_n353), .B2(new_n219), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n285), .A2(new_n207), .A3(new_n286), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n352), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n347), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n345), .B1(new_n359), .B2(G68), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n276), .B1(new_n360), .B2(KEYINPUT16), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n339), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n281), .A2(new_n282), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n294), .A2(new_n296), .A3(G223), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G226), .A2(G1698), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G87), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n273), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n278), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n306), .A2(G232), .B1(new_n310), .B2(new_n305), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n369), .A2(G190), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n369), .B2(new_n370), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT17), .B1(new_n362), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(G20), .B1(new_n283), .B2(new_n287), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n347), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n345), .B1(new_n377), .B2(G68), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n361), .B1(new_n378), .B2(KEYINPUT16), .ZN(new_n379));
  INV_X1    g0179(.A(new_n253), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT70), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n267), .ZN(new_n382));
  NAND2_X1  g0182(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n340), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n268), .B1(new_n384), .B2(new_n270), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n254), .B1(new_n385), .B2(new_n266), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n380), .B1(new_n386), .B2(KEYINPUT76), .ZN(new_n387));
  INV_X1    g0187(.A(new_n338), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n330), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n379), .A2(new_n389), .A3(new_n374), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT77), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT77), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n379), .A2(new_n389), .A3(new_n374), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n375), .B1(new_n394), .B2(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n379), .A2(new_n389), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n369), .B2(new_n370), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n369), .A2(new_n370), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(G179), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n402), .B(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n306), .A2(G244), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n310), .A2(new_n305), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g0208(.A(new_n408), .B(KEYINPUT72), .Z(new_n409));
  AOI21_X1  g0209(.A(new_n220), .B1(new_n290), .B2(new_n291), .ZN(new_n410));
  INV_X1    g0210(.A(G232), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n299), .A2(new_n411), .B1(new_n203), .B2(new_n293), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n308), .A2(new_n309), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n415), .A2(G200), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  INV_X1    g0217(.A(new_n274), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(new_n207), .B2(new_n221), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT8), .B(G58), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(new_n260), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n252), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT73), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n329), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n250), .A2(KEYINPUT74), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n252), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(G77), .A3(new_n332), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(G77), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G190), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n415), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n416), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n415), .A2(G179), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n431), .B1(new_n415), .B2(new_n397), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n327), .A2(new_n405), .A3(new_n434), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n219), .A2(G20), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n439), .B1(new_n260), .B2(new_n255), .C1(new_n418), .C2(new_n221), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n252), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT11), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n427), .A2(G68), .A3(new_n332), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n328), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n445), .A2(KEYINPUT12), .A3(new_n439), .ZN(new_n446));
  INV_X1    g0246(.A(new_n429), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n219), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n448), .B2(KEYINPUT12), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT14), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n306), .A2(G238), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n407), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n283), .A2(new_n287), .A3(G232), .A4(G1698), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(KEYINPUT75), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(KEYINPUT75), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n298), .A2(new_n283), .A3(new_n287), .A4(G226), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n273), .B2(new_n202), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n454), .B1(new_n462), .B2(new_n278), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT13), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n460), .B1(new_n456), .B2(new_n457), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n453), .B(new_n407), .C1(new_n466), .C2(new_n414), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(KEYINPUT13), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n452), .B(G169), .C1(new_n465), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n463), .A2(new_n464), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(KEYINPUT13), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(G179), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n471), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n452), .B1(new_n474), .B2(G169), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n451), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n450), .B1(new_n474), .B2(new_n432), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n372), .B1(new_n470), .B2(new_n471), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n438), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  AND2_X1   g0283(.A1(G264), .A2(G1698), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n281), .B2(new_n282), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n285), .A2(new_n286), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(KEYINPUT81), .A3(new_n484), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(G303), .B1(new_n349), .B2(new_n350), .ZN(new_n491));
  INV_X1    g0291(.A(G257), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n285), .B2(new_n286), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n298), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n288), .A2(G303), .B1(new_n298), .B2(new_n493), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT82), .A3(new_n490), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n414), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT79), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(G41), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n304), .A2(G1), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n303), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n506), .A2(new_n307), .A3(new_n278), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n506), .A2(new_n414), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(G270), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n483), .B1(new_n500), .B2(new_n510), .ZN(new_n511));
  AND4_X1   g0311(.A1(KEYINPUT82), .A2(new_n490), .A3(new_n494), .A4(new_n491), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT82), .B1(new_n498), .B2(new_n490), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n278), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(KEYINPUT83), .A3(new_n509), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G283), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n517), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n252), .C1(new_n207), .C2(G116), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT20), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n521), .A2(new_n522), .B1(new_n447), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n206), .B2(G33), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n427), .A2(KEYINPUT84), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT84), .B1(new_n427), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G169), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n516), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT85), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n516), .A2(G200), .ZN(new_n535));
  INV_X1    g0335(.A(new_n528), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n511), .A2(new_n515), .A3(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n529), .B1(new_n511), .B2(new_n515), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT21), .B1(new_n539), .B2(KEYINPUT85), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n509), .A2(G179), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n497), .A2(new_n499), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n278), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n528), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n534), .A2(new_n538), .A3(new_n540), .A4(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT78), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n329), .B2(G97), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n250), .A2(KEYINPUT78), .A3(new_n202), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n253), .B1(G1), .B2(new_n273), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n202), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n552), .A2(new_n202), .A3(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(G97), .B(G107), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n555), .A2(new_n207), .B1(new_n221), .B2(new_n260), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n377), .B2(G107), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n551), .B1(new_n557), .B2(new_n276), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n222), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n298), .A2(new_n283), .A3(new_n287), .A4(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n283), .A2(new_n287), .A3(G250), .A4(G1698), .ZN(new_n563));
  OAI21_X1  g0363(.A(G244), .B1(new_n281), .B2(new_n282), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n560), .B1(new_n564), .B2(new_n297), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n562), .A2(new_n563), .A3(new_n565), .A4(new_n517), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n278), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n507), .B1(G257), .B2(new_n508), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G200), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n559), .B(new_n570), .C1(new_n432), .C2(new_n569), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n397), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n558), .C1(G179), .C2(new_n569), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G116), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n294), .B(new_n296), .C1(new_n281), .C2(new_n282), .ZN(new_n576));
  OAI221_X1 g0376(.A(new_n575), .B1(new_n564), .B2(new_n289), .C1(new_n220), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n278), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n504), .A2(new_n307), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n414), .C1(G250), .C2(new_n504), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n488), .A2(new_n207), .A3(G68), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n584), .A2(new_n273), .A3(new_n202), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n585), .A2(G20), .B1(G87), .B2(new_n204), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n274), .A2(G97), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n584), .ZN(new_n589));
  AOI211_X1 g0389(.A(KEYINPUT80), .B(KEYINPUT19), .C1(new_n274), .C2(G97), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n583), .B(new_n586), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n252), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n447), .A2(new_n417), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n578), .A2(G190), .A3(new_n580), .ZN(new_n595));
  INV_X1    g0395(.A(new_n549), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G87), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n582), .A2(new_n594), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n581), .A2(new_n397), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n592), .B(new_n593), .C1(new_n417), .C2(new_n549), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n578), .A2(new_n315), .A3(new_n580), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n574), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n545), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n549), .A2(new_n203), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n250), .A2(new_n203), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT25), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n575), .A2(G20), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT86), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT23), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n207), .B2(G107), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT87), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n615), .A2(new_n616), .B1(new_n617), .B2(KEYINPUT24), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n488), .A2(new_n207), .A3(G87), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT22), .ZN(new_n621));
  OR3_X1    g0421(.A1(new_n367), .A2(KEYINPUT22), .A3(G20), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n288), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n617), .A2(KEYINPUT24), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n276), .B1(new_n624), .B2(new_n625), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n611), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n506), .A2(G264), .A3(new_n414), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT88), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n506), .A2(new_n631), .A3(new_n414), .A4(G264), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n634));
  INV_X1    g0434(.A(G294), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n273), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G250), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n576), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n278), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n633), .A2(KEYINPUT89), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT89), .B1(new_n633), .B2(new_n639), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n640), .A2(new_n641), .A3(new_n507), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G179), .ZN(new_n643));
  INV_X1    g0443(.A(new_n507), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n633), .A2(new_n644), .A3(new_n639), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G169), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n628), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n642), .A2(G200), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n645), .A2(G190), .ZN(new_n649));
  OAI211_X1 g0449(.A(KEYINPUT90), .B(new_n628), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n633), .A2(new_n639), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n633), .A2(KEYINPUT89), .A3(new_n639), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n644), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n649), .B1(new_n656), .B2(new_n372), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n626), .A2(new_n627), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n610), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n651), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n647), .B1(new_n650), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n482), .A2(new_n606), .A3(new_n661), .ZN(G372));
  INV_X1    g0462(.A(new_n475), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n472), .A3(new_n469), .ZN(new_n664));
  INV_X1    g0464(.A(new_n437), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n451), .A2(new_n664), .B1(new_n480), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n395), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n404), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n324), .A2(new_n326), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n316), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n482), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n571), .A2(new_n573), .A3(new_n598), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n650), .B2(new_n660), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n534), .A2(new_n540), .A3(new_n544), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n646), .B1(new_n656), .B2(new_n315), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n675), .A2(KEYINPUT91), .A3(new_n659), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT91), .B1(new_n675), .B2(new_n659), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n673), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n602), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n603), .A2(new_n573), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n603), .B2(new_n573), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n670), .B1(new_n671), .B2(new_n687), .ZN(G369));
  OR3_X1    g0488(.A1(new_n445), .A2(KEYINPUT27), .A3(G20), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT27), .B1(new_n445), .B2(G20), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n536), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n545), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n674), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n661), .B1(new_n628), .B2(new_n694), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n647), .A2(new_n693), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(G330), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n674), .A2(new_n694), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT92), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT92), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n674), .B2(new_n694), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n701), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n678), .A2(new_n694), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n702), .A2(new_n707), .A3(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n210), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n213), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g0515(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n716));
  XNOR2_X1  g0516(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT94), .B1(new_n500), .B2(new_n541), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT94), .ZN(new_n720));
  INV_X1    g0520(.A(new_n541), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n514), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n640), .A2(new_n641), .A3(new_n581), .ZN(new_n723));
  INV_X1    g0523(.A(new_n569), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n719), .A2(new_n722), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n569), .A2(new_n315), .A3(new_n581), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n642), .A2(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n725), .A2(new_n726), .B1(new_n728), .B2(new_n516), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n569), .A2(new_n726), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n719), .A2(new_n722), .A3(new_n723), .A4(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT95), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n729), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n578), .A2(new_n580), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n654), .A2(new_n737), .A3(new_n655), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n720), .B2(new_n543), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(KEYINPUT95), .A3(new_n719), .A4(new_n730), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n731), .A2(new_n732), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT96), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(new_n743), .A3(new_n729), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n736), .A2(new_n693), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n694), .A2(new_n746), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n742), .B2(new_n729), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n693), .B(new_n647), .C1(new_n650), .C2(new_n660), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n750), .B1(new_n606), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n718), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT29), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n673), .B1(new_n674), .B2(new_n647), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n684), .B1(new_n682), .B2(KEYINPUT97), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT97), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n758), .B(new_n681), .C1(new_n603), .C2(new_n573), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n680), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n755), .B1(new_n761), .B2(new_n694), .ZN(new_n762));
  AOI211_X1 g0562(.A(KEYINPUT29), .B(new_n693), .C1(new_n679), .C2(new_n685), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n754), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n717), .B1(new_n766), .B2(G1), .ZN(G364));
  NAND2_X1  g0567(.A1(new_n698), .A2(G330), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n696), .A2(new_n718), .A3(new_n697), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n249), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n206), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n711), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n768), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n215), .B1(G20), .B2(new_n397), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(new_n315), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n782), .A2(new_n432), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n432), .A2(new_n372), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n784), .A2(new_n340), .B1(new_n786), .B2(new_n255), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n432), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n207), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n288), .B(new_n787), .C1(G97), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n207), .A2(G179), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n372), .A2(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT99), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G107), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n781), .A2(new_n798), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n785), .A2(new_n792), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n219), .A2(new_n802), .B1(new_n803), .B2(new_n367), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n781), .A2(new_n793), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(G77), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n791), .A2(new_n797), .A3(new_n801), .A4(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n786), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G326), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n784), .B2(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n293), .B(new_n812), .C1(G294), .C2(new_n790), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n803), .B(KEYINPUT100), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G303), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n800), .A2(G283), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n805), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G317), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n819), .A2(KEYINPUT33), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(KEYINPUT33), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n802), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n794), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n818), .B(new_n822), .C1(G329), .C2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n813), .A2(new_n815), .A3(new_n816), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n780), .B1(new_n808), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(G13), .A2(G33), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(G20), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n779), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n213), .A2(G45), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n210), .A2(new_n363), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(new_n247), .C2(G45), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n293), .A2(new_n210), .ZN(new_n834));
  INV_X1    g0634(.A(G355), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n834), .A2(new_n835), .B1(G116), .B2(new_n210), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n774), .B(new_n826), .C1(new_n830), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n829), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n698), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n775), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n780), .A2(new_n828), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n773), .B1(new_n843), .B2(G77), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n783), .A2(G143), .B1(new_n809), .B2(G137), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n261), .B2(new_n802), .C1(new_n795), .C2(new_n805), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT34), .Z(new_n847));
  NAND2_X1  g0647(.A1(new_n814), .A2(G50), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n800), .A2(G68), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n790), .A2(G58), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n363), .B1(new_n823), .B2(G132), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n802), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT101), .B(G283), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n783), .A2(G294), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(new_n288), .C1(new_n202), .C2(new_n789), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n800), .A2(G87), .ZN(new_n858));
  INV_X1    g0658(.A(G303), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n786), .A2(new_n859), .B1(new_n805), .B2(new_n523), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G311), .B2(new_n823), .ZN(new_n861));
  INV_X1    g0661(.A(new_n814), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n858), .B(new_n861), .C1(new_n862), .C2(new_n203), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n847), .A2(new_n852), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n844), .B1(new_n864), .B2(new_n779), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n416), .A2(new_n433), .B1(new_n431), .B2(new_n694), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n437), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n435), .A2(new_n436), .A3(new_n694), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n865), .B1(new_n870), .B2(new_n828), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(new_n687), .B2(new_n693), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n686), .A2(new_n694), .A3(new_n870), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n773), .B1(new_n874), .B2(new_n754), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n754), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(G384));
  NOR2_X1   g0678(.A1(new_n770), .A2(new_n206), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n482), .B1(new_n762), .B2(new_n763), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n670), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT103), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n390), .B1(new_n362), .B2(new_n400), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n362), .A2(new_n691), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT37), .B1(new_n396), .B2(new_n401), .ZN(new_n887));
  INV_X1    g0687(.A(new_n691), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n396), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n887), .A2(new_n391), .A3(new_n393), .A4(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT102), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT102), .B1(new_n886), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n395), .B2(new_n404), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n219), .B1(new_n358), .B2(new_n347), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n355), .B1(new_n897), .B2(new_n345), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n361), .A2(new_n898), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n401), .A2(new_n888), .B1(new_n899), .B2(new_n339), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n391), .A3(new_n393), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n902), .A2(new_n890), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n888), .B1(new_n899), .B2(new_n339), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n395), .B2(new_n404), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n883), .B1(new_n896), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n664), .A2(new_n451), .A3(new_n694), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n902), .A2(new_n890), .ZN(new_n911));
  OAI211_X1 g0711(.A(KEYINPUT38), .B(new_n911), .C1(new_n405), .C2(new_n904), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n906), .B1(new_n903), .B2(new_n905), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT39), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n908), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n451), .B(new_n693), .C1(new_n664), .C2(new_n479), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n450), .A2(new_n694), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n476), .A2(new_n480), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n912), .A2(new_n913), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n693), .B(new_n869), .C1(new_n679), .C2(new_n685), .ZN(new_n922));
  INV_X1    g0722(.A(new_n868), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n920), .B(new_n921), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n404), .A2(new_n888), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n915), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n882), .B(new_n926), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n894), .A2(new_n891), .A3(new_n892), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n912), .B1(new_n928), .B2(KEYINPUT38), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n869), .B1(new_n916), .B2(new_n919), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n742), .A2(new_n743), .A3(new_n729), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n743), .B1(new_n742), .B2(new_n729), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT31), .B1(new_n933), .B2(new_n693), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n736), .A2(new_n744), .A3(new_n748), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n534), .A2(new_n540), .A3(new_n544), .ZN(new_n936));
  INV_X1    g0736(.A(new_n605), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n751), .A2(new_n936), .A3(new_n538), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n929), .B(new_n930), .C1(new_n934), .C2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT40), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT40), .B1(new_n912), .B2(new_n913), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n942), .B(new_n930), .C1(new_n934), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n935), .A2(new_n938), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n671), .B1(new_n747), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n718), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n944), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n879), .B1(new_n927), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n927), .B2(new_n948), .ZN(new_n950));
  INV_X1    g0750(.A(new_n555), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT35), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(G116), .A3(new_n216), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n341), .A2(new_n213), .A3(new_n221), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n219), .A2(G50), .ZN(new_n957));
  OAI211_X1 g0757(.A(G1), .B(new_n249), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n950), .A2(new_n955), .A3(new_n958), .ZN(G367));
  INV_X1    g0759(.A(KEYINPUT104), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n594), .A2(new_n597), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n693), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n604), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n602), .B2(new_n962), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT43), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n703), .B(KEYINPUT92), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n574), .B1(new_n559), .B2(new_n694), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n573), .A2(new_n694), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n966), .A2(KEYINPUT42), .A3(new_n701), .A4(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n701), .B(new_n969), .C1(new_n704), .C2(new_n706), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT42), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n675), .A2(new_n659), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n573), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n694), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n960), .B(new_n965), .C1(new_n974), .C2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n977), .B1(new_n970), .B2(new_n973), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n965), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT104), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n978), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(KEYINPUT105), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n969), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n702), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n984), .A2(KEYINPUT105), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n984), .A2(KEYINPUT105), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n991), .A2(new_n985), .B1(new_n702), .B2(new_n987), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n711), .B(KEYINPUT41), .Z(new_n993));
  AOI21_X1  g0793(.A(new_n969), .B1(new_n707), .B2(new_n708), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n707), .A2(new_n708), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(new_n987), .A3(new_n995), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n707), .A2(new_n708), .A3(new_n969), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1000), .B(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n999), .A2(new_n1004), .A3(new_n702), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n966), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n702), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n701), .B1(new_n698), .B2(G330), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1008), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(new_n702), .A3(new_n966), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n765), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n996), .A2(new_n998), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1007), .B1(new_n1014), .B2(new_n1003), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1005), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n993), .B1(new_n1016), .B2(new_n766), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n990), .B(new_n992), .C1(new_n772), .C2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n830), .B1(new_n210), .B2(new_n417), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n239), .A2(new_n832), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n773), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n786), .A2(new_n817), .B1(new_n802), .B2(new_n635), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n488), .B(new_n1022), .C1(G317), .C2(new_n823), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n803), .A2(new_n523), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1023), .B1(KEYINPUT46), .B2(new_n1024), .C1(new_n203), .C2(new_n789), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n814), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n799), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n783), .A2(G303), .B1(G97), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(new_n805), .C2(new_n854), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n784), .A2(new_n261), .B1(new_n221), .B2(new_n799), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n803), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1030), .B1(G58), .B2(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n255), .A2(new_n805), .B1(new_n802), .B2(new_n795), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT108), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT108), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n809), .A2(G143), .B1(new_n823), .B2(G137), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n293), .C1(new_n219), .C2(new_n789), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1025), .A2(new_n1029), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT47), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n780), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1021), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n964), .B2(new_n839), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1018), .A2(new_n1044), .ZN(G387));
  NAND2_X1  g0845(.A1(new_n1012), .A2(new_n765), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT109), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1013), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(KEYINPUT109), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1047), .A2(new_n711), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1012), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n699), .A2(new_n700), .A3(new_n829), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n789), .A2(new_n854), .B1(new_n803), .B2(new_n635), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G303), .A2(new_n806), .B1(new_n853), .B2(G311), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n811), .B2(new_n786), .C1(new_n819), .C2(new_n784), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT49), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n488), .B1(new_n823), .B2(G326), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n523), .C2(new_n799), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n803), .A2(new_n221), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n786), .A2(new_n795), .B1(new_n805), .B2(new_n219), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G50), .C2(new_n783), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n789), .A2(new_n417), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n363), .B(new_n1065), .C1(G150), .C2(new_n823), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n272), .A2(new_n853), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n800), .A2(G97), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n780), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n236), .A2(new_n304), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1071), .A2(new_n832), .B1(new_n713), .B2(new_n834), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n420), .A2(G50), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT50), .ZN(new_n1074));
  AOI21_X1  g0874(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n713), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(G107), .B2(new_n210), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n774), .B(new_n1070), .C1(new_n830), .C2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1051), .A2(new_n772), .B1(new_n1052), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1050), .A2(new_n1080), .ZN(G393));
  NAND3_X1  g0881(.A1(new_n1005), .A2(new_n772), .A3(new_n1015), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n244), .A2(new_n210), .A3(new_n363), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n830), .B1(new_n202), .B2(new_n210), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n773), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n783), .A2(G159), .B1(new_n809), .B2(G150), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT51), .Z(new_n1087));
  NAND2_X1  g0887(.A1(new_n853), .A2(G50), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n803), .B2(new_n219), .C1(new_n420), .C2(new_n805), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n789), .A2(new_n221), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n363), .B(new_n1091), .C1(G143), .C2(new_n823), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1087), .A2(new_n858), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n784), .A2(new_n817), .B1(new_n786), .B2(new_n819), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1031), .A2(new_n855), .B1(new_n823), .B2(G322), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1096), .B1(KEYINPUT111), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n635), .A2(new_n805), .B1(new_n802), .B2(new_n859), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n293), .B(new_n1102), .C1(G116), .C2(new_n790), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n801), .C1(KEYINPUT111), .C2(new_n1098), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1093), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1085), .B1(new_n1105), .B2(new_n779), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n969), .B2(new_n839), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1082), .A2(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1016), .A2(new_n711), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1005), .A2(new_n1015), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n765), .B2(new_n1012), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G390));
  AOI21_X1  g0913(.A(new_n693), .B1(new_n756), .B2(new_n760), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n923), .B1(new_n1114), .B2(new_n867), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n476), .A2(new_n480), .A3(new_n918), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n918), .B1(new_n476), .B2(new_n480), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n909), .B(new_n929), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n747), .A2(new_n752), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1120), .A2(G330), .A3(new_n920), .A4(new_n870), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n873), .A2(new_n868), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n910), .B1(new_n1122), .B2(new_n920), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n908), .A2(new_n914), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1119), .B(new_n1121), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT112), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n908), .A2(new_n914), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1118), .B1(new_n873), .B2(new_n868), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n910), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT112), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1129), .A2(new_n1130), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1119), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n718), .B1(new_n945), .B2(new_n747), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n930), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1126), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n772), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n773), .B1(new_n843), .B2(new_n272), .ZN(new_n1139));
  INV_X1    g0939(.A(G283), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n786), .A2(new_n1140), .B1(new_n805), .B2(new_n202), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G294), .B2(new_n823), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n849), .B(new_n1142), .C1(new_n862), .C2(new_n367), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n783), .A2(G116), .B1(G107), .B2(new_n853), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(new_n288), .C1(new_n221), .C2(new_n789), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n803), .A2(new_n261), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT53), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT54), .B(G143), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G128), .A2(new_n809), .B1(new_n806), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1027), .A2(G50), .B1(new_n823), .B2(G125), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n783), .A2(G132), .B1(G137), .B2(new_n853), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n293), .C1(new_n795), .C2(new_n789), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1143), .A2(new_n1145), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1139), .B1(new_n1155), .B2(new_n779), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1124), .B2(new_n828), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n920), .B1(new_n1133), .B2(new_n870), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1121), .A2(new_n1115), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n920), .B1(new_n753), .B2(new_n870), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT114), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n718), .B(new_n869), .C1(new_n747), .C2(new_n752), .ZN(new_n1164));
  OAI21_X1  g0964(.A(KEYINPUT114), .B1(new_n1164), .B2(new_n920), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1165), .A3(new_n1134), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1160), .B1(new_n1166), .B2(new_n1122), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n482), .B(G330), .C1(new_n934), .C2(new_n939), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n880), .A2(new_n1168), .A3(new_n670), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT113), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n880), .A2(new_n1168), .A3(new_n670), .A4(KEYINPUT113), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n711), .B1(new_n1174), .B2(new_n1137), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1134), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1164), .A2(KEYINPUT114), .A3(new_n920), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1122), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1173), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1126), .A2(new_n1136), .A3(new_n1131), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1138), .B(new_n1157), .C1(new_n1175), .C2(new_n1184), .ZN(G378));
  OAI21_X1  g0985(.A(new_n1181), .B1(new_n1183), .B2(new_n1167), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n277), .A2(new_n888), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT55), .Z(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n327), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n327), .A2(new_n1189), .ZN(new_n1194));
  OR3_X1    g0994(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n944), .A2(G330), .A3(new_n926), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n926), .B1(new_n944), .B2(G330), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n915), .A2(new_n924), .A3(new_n925), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n870), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n945), .B2(new_n747), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1203), .A2(new_n942), .B1(new_n940), .B2(KEYINPUT40), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1204), .B2(new_n718), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n944), .A2(G330), .A3(new_n926), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1197), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1200), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1186), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1200), .B2(new_n1208), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n712), .B1(new_n1213), .B2(new_n1186), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT119), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n771), .B1(new_n1200), .B2(new_n1208), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n773), .B1(new_n843), .B2(G50), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n794), .A2(new_n1140), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n805), .A2(new_n417), .B1(new_n799), .B2(new_n340), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(G107), .C2(new_n783), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n303), .B(new_n363), .C1(new_n802), .C2(new_n202), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1062), .B(new_n1222), .C1(G116), .C2(new_n809), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(new_n219), .C2(new_n789), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n363), .A2(new_n303), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G50), .B1(new_n273), .B2(new_n303), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1224), .A2(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT115), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G125), .A2(new_n809), .B1(new_n1031), .B2(new_n1149), .ZN(new_n1230));
  INV_X1    g1030(.A(G128), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n784), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G132), .A2(new_n853), .B1(new_n806), .B2(G137), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT116), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(G150), .C2(new_n790), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1027), .A2(G159), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n823), .C2(G124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1229), .B1(new_n1225), .B2(new_n1224), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1218), .B1(new_n1242), .B2(new_n779), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1197), .B2(new_n828), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT118), .Z(new_n1245));
  OAI21_X1  g1045(.A(new_n1216), .B1(new_n1217), .B2(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1207), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n772), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1245), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(KEYINPUT119), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1246), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1215), .A2(new_n1252), .ZN(G375));
  INV_X1    g1053(.A(new_n993), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1178), .A2(new_n1173), .A3(new_n1179), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1182), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT120), .Z(new_n1257));
  NAND2_X1  g1057(.A1(new_n1118), .A2(new_n827), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n773), .B1(new_n843), .B2(G68), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n784), .A2(new_n1140), .B1(new_n786), .B2(new_n635), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G107), .B2(new_n806), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n800), .A2(G77), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n202), .C2(new_n862), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G116), .A2(new_n853), .B1(new_n823), .B2(G303), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(new_n288), .C1(new_n417), .C2(new_n789), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n805), .A2(new_n261), .B1(new_n794), .B2(new_n1231), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n363), .B(new_n1266), .C1(G58), .C2(new_n1027), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1267), .B1(new_n255), .B2(new_n789), .C1(new_n862), .C2(new_n795), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G132), .A2(new_n809), .B1(new_n853), .B2(new_n1149), .ZN(new_n1269));
  INV_X1    g1069(.A(G137), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n784), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT121), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1263), .A2(new_n1265), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1259), .B1(new_n1273), .B2(new_n779), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1180), .A2(new_n772), .B1(new_n1258), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1257), .A2(new_n1275), .ZN(G381));
  AND3_X1   g1076(.A1(new_n1018), .A2(new_n1044), .A3(new_n1112), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1050), .A2(new_n841), .A3(new_n1080), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(G378), .A2(new_n1278), .A3(G384), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1277), .A2(new_n1279), .A3(new_n1275), .A4(new_n1257), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1280), .A2(G375), .ZN(G407));
  NAND2_X1  g1081(.A1(new_n1138), .A2(new_n1157), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1174), .A2(new_n1137), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n712), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n692), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G407), .B(G213), .C1(G375), .C2(new_n1286), .ZN(G409));
  NAND2_X1  g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1278), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1112), .B1(new_n1018), .B2(new_n1044), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1277), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G387), .A2(G390), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1018), .A2(new_n1044), .A3(new_n1112), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1289), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n712), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1178), .A2(KEYINPUT60), .A3(new_n1173), .A4(new_n1179), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT122), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT122), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1167), .A2(new_n1301), .A3(KEYINPUT60), .A4(new_n1173), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1255), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1298), .A2(new_n1300), .A3(new_n1302), .A4(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(G384), .A3(new_n1275), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT123), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT123), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1305), .A2(new_n1308), .A3(G384), .A4(new_n1275), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1275), .ZN(new_n1310));
  INV_X1    g1110(.A(G384), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1307), .A2(new_n1309), .A3(new_n1312), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n692), .A2(G213), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1215), .A2(new_n1252), .A3(G378), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1210), .A2(new_n993), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1285), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1314), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1314), .A2(G2897), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1313), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1307), .A2(new_n1309), .A3(new_n1312), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1320), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1325), .A2(new_n1326), .A3(new_n1330), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1319), .A2(KEYINPUT62), .A3(new_n1323), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT62), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1328), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1297), .B1(new_n1331), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT124), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1325), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1292), .A2(new_n1295), .A3(new_n1326), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT63), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1338), .B1(new_n1339), .B2(new_n1327), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1322), .A2(KEYINPUT124), .A3(new_n1324), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1319), .A2(new_n1323), .A3(KEYINPUT63), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1337), .A2(new_n1340), .A3(new_n1341), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1335), .A2(new_n1343), .ZN(G405));
  INV_X1    g1144(.A(new_n1315), .ZN(new_n1345));
  AOI21_X1  g1145(.A(G378), .B1(new_n1215), .B2(new_n1252), .ZN(new_n1346));
  OR3_X1    g1146(.A1(new_n1345), .A2(new_n1313), .A3(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1313), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1347), .A2(new_n1296), .A3(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1296), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT126), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  AOI211_X1 g1152(.A(KEYINPUT126), .B(new_n1296), .C1(new_n1347), .C2(new_n1348), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(G402));
endmodule


