//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n585, new_n586,
    new_n587, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n608, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n647, new_n648, new_n649, new_n652, new_n654,
    new_n655, new_n656, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AND2_X1   g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  OR2_X1    g038(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(KEYINPUT3), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT69), .B(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G101), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(KEYINPUT70), .A3(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  INV_X1    g056(.A(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n468), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G125), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n471), .A2(new_n480), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NOR2_X1   g064(.A1(new_n469), .A2(new_n474), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT72), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(KEYINPUT72), .A2(G100), .A3(G2105), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G112), .B2(new_n474), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n470), .A2(G136), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n492), .A2(new_n496), .A3(new_n497), .ZN(G162));
  NAND4_X1  g073(.A1(new_n466), .A2(G138), .A3(new_n474), .A4(new_n468), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n474), .A2(G138), .ZN(new_n501));
  OR2_X1    g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n484), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G114), .C2(new_n474), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n503), .A2(KEYINPUT73), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n484), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n511), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n512), .B2(new_n507), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(KEYINPUT76), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n518), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT77), .B1(new_n525), .B2(new_n518), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(G62), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT74), .B(G651), .Z(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT75), .A2(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(KEYINPUT6), .ZN(new_n534));
  OAI21_X1  g109(.A(KEYINPUT6), .B1(KEYINPUT74), .B2(G651), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(KEYINPUT74), .A2(KEYINPUT75), .A3(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n516), .A2(KEYINPUT76), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n523), .B(G543), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n517), .ZN(new_n542));
  AND4_X1   g117(.A1(new_n526), .A2(new_n538), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n537), .B(KEYINPUT6), .C1(KEYINPUT74), .C2(G651), .ZN(new_n544));
  INV_X1    g119(.A(new_n534), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(new_n545), .A3(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n543), .A2(G88), .B1(G50), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n532), .A2(new_n548), .A3(KEYINPUT78), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n530), .B1(new_n527), .B2(new_n528), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n526), .A2(new_n538), .A3(new_n541), .A4(new_n542), .ZN(new_n552));
  INV_X1    g127(.A(G88), .ZN(new_n553));
  INV_X1    g128(.A(G50), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n552), .A2(new_n553), .B1(new_n554), .B2(new_n546), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n549), .A2(new_n556), .ZN(G166));
  AND3_X1   g132(.A1(new_n526), .A2(new_n542), .A3(new_n541), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n558), .A2(G63), .A3(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n543), .A2(G89), .ZN(new_n560));
  NAND3_X1  g135(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT7), .Z(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n547), .B2(G51), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(G286));
  INV_X1    g139(.A(G286), .ZN(G168));
  NAND2_X1  g140(.A1(G77), .A2(G543), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n526), .A2(new_n542), .A3(new_n541), .ZN(new_n567));
  INV_X1    g142(.A(G64), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(new_n531), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT79), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n543), .A2(G90), .B1(G52), .B2(new_n547), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n570), .A2(KEYINPUT79), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(G171));
  NAND3_X1  g150(.A1(new_n524), .A2(G56), .A3(new_n526), .ZN(new_n576));
  NAND2_X1  g151(.A1(G68), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n530), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G81), .ZN(new_n579));
  INV_X1    g154(.A(G43), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n552), .A2(new_n579), .B1(new_n580), .B2(new_n546), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G860), .ZN(G153));
  NAND4_X1  g158(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g159(.A1(G1), .A2(G3), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT80), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT8), .ZN(new_n587));
  NAND4_X1  g162(.A1(G319), .A2(G483), .A3(G661), .A4(new_n587), .ZN(G188));
  INV_X1    g163(.A(G65), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n541), .A2(new_n542), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n522), .A2(new_n523), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n524), .A2(KEYINPUT83), .A3(new_n526), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n589), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G78), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(KEYINPUT81), .A2(G53), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n546), .A2(KEYINPUT9), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT9), .B1(new_n546), .B2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n524), .A2(new_n604), .A3(new_n526), .A4(new_n538), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(G91), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n598), .A2(new_n602), .A3(new_n606), .ZN(G299));
  INV_X1    g182(.A(new_n574), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n608), .A2(new_n571), .A3(new_n572), .ZN(G301));
  INV_X1    g184(.A(G166), .ZN(G303));
  INV_X1    g185(.A(G74), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n567), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G49), .B2(new_n547), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n603), .A2(G87), .A3(new_n605), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(G288));
  NAND2_X1  g190(.A1(new_n547), .A2(G48), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n558), .A2(KEYINPUT84), .A3(G61), .ZN(new_n618));
  NAND2_X1  g193(.A1(G73), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n620));
  INV_X1    g195(.A(G61), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n567), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(new_n531), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n603), .A2(G86), .A3(new_n605), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(G305));
  AOI22_X1  g201(.A1(new_n558), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(new_n530), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n543), .A2(G85), .B1(G47), .B2(new_n547), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(G290));
  NAND2_X1  g205(.A1(G301), .A2(G868), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n603), .A2(G92), .A3(new_n605), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n603), .A2(KEYINPUT10), .A3(G92), .A4(new_n605), .ZN(new_n635));
  AND2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G66), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n593), .B2(new_n594), .ZN(new_n638));
  NAND2_X1  g213(.A1(G79), .A2(G543), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(G651), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n547), .A2(G54), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n631), .B1(new_n644), .B2(G868), .ZN(G284));
  OAI21_X1  g220(.A(new_n631), .B1(new_n644), .B2(G868), .ZN(G321));
  INV_X1    g221(.A(G868), .ZN(new_n647));
  NOR2_X1   g222(.A1(G286), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G299), .B(KEYINPUT85), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(new_n647), .ZN(G297));
  AOI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n647), .ZN(G280));
  XNOR2_X1  g226(.A(KEYINPUT86), .B(G559), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n644), .B1(G860), .B2(new_n652), .ZN(G148));
  NAND2_X1  g228(.A1(new_n644), .A2(new_n652), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT87), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n655), .A2(new_n647), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n647), .B2(new_n582), .ZN(G323));
  XNOR2_X1  g232(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g233(.A1(new_n490), .A2(G123), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n474), .A2(G111), .ZN(new_n660));
  OAI21_X1  g235(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(G135), .B2(new_n470), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT89), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(G2096), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(G2096), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n475), .A2(new_n484), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT12), .ZN(new_n668));
  INV_X1    g243(.A(G2100), .ZN(new_n669));
  OAI22_X1  g244(.A1(new_n668), .A2(KEYINPUT13), .B1(KEYINPUT88), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(KEYINPUT13), .B2(new_n668), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(KEYINPUT88), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n665), .A2(new_n666), .A3(new_n673), .ZN(G156));
  XNOR2_X1  g249(.A(KEYINPUT15), .B(G2435), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2438), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2427), .B(G2430), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(KEYINPUT14), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT90), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n676), .B2(new_n677), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2443), .B(G2446), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1341), .B(G1348), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2451), .B(G2454), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT16), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n687), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n688), .A2(new_n689), .A3(G14), .ZN(G401));
  XOR2_X1   g265(.A(G2072), .B(G2078), .Z(new_n691));
  XOR2_X1   g266(.A(G2084), .B(G2090), .Z(new_n692));
  XNOR2_X1  g267(.A(G2067), .B(G2678), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n691), .B1(new_n694), .B2(KEYINPUT18), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT91), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2100), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT18), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(KEYINPUT17), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n692), .A2(new_n693), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G2096), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n697), .B(new_n702), .ZN(G227));
  XOR2_X1   g278(.A(G1971), .B(G1976), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT19), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1956), .B(G2474), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1961), .B(G1966), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n706), .A2(new_n707), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n705), .A2(new_n710), .A3(new_n708), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n705), .A2(new_n710), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n713));
  AOI211_X1 g288(.A(new_n709), .B(new_n711), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT93), .ZN(new_n716));
  XOR2_X1   g291(.A(G1981), .B(G1986), .Z(new_n717));
  XNOR2_X1  g292(.A(G1991), .B(G1996), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n716), .B(new_n721), .ZN(G229));
  INV_X1    g297(.A(G28), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(KEYINPUT30), .ZN(new_n725));
  OR2_X1    g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n729), .B2(KEYINPUT24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(KEYINPUT24), .B2(new_n729), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n488), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n728), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n664), .A2(new_n732), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n735), .B(new_n736), .C1(new_n734), .C2(new_n733), .ZN(new_n737));
  INV_X1    g312(.A(G16), .ZN(new_n738));
  NOR2_X1   g313(.A1(G168), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(G21), .ZN(new_n740));
  INV_X1    g315(.A(G1966), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n732), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n732), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT29), .B(G2090), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n470), .A2(G140), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n490), .A2(G128), .ZN(new_n748));
  INV_X1    g323(.A(G104), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n749), .A2(new_n474), .A3(KEYINPUT95), .ZN(new_n750));
  AOI21_X1  g325(.A(KEYINPUT95), .B1(new_n749), .B2(new_n474), .ZN(new_n751));
  OAI221_X1 g326(.A(G2104), .B1(G116), .B2(new_n474), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n747), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n732), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n740), .B2(new_n741), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n737), .A2(new_n742), .A3(new_n746), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(G164), .A2(G29), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G27), .B2(G29), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n582), .A2(new_n738), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n738), .B2(G19), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G1341), .ZN(new_n768));
  NAND2_X1  g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  INV_X1    g344(.A(G127), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n484), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n474), .B1(new_n771), .B2(KEYINPUT96), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT96), .B2(new_n771), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT25), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n470), .B2(G139), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT97), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(new_n732), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n732), .B2(G33), .ZN(new_n780));
  INV_X1    g355(.A(G2072), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G1341), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n766), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n760), .A2(new_n764), .A3(new_n768), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n738), .A2(G20), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT23), .Z(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT99), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1956), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n732), .A2(G32), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n470), .A2(G141), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n490), .A2(G129), .ZN(new_n793));
  NAND3_X1  g368(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT26), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  AOI22_X1  g372(.A1(G105), .A2(new_n478), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n792), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n791), .B1(new_n800), .B2(new_n732), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT27), .ZN(new_n802));
  INV_X1    g377(.A(G1996), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n762), .A2(new_n763), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n780), .B2(new_n781), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  NOR2_X1   g382(.A1(G171), .A2(new_n738), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G5), .B2(new_n738), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n804), .B(new_n806), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n785), .A2(new_n790), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n807), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT98), .Z(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G1956), .B2(new_n789), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n738), .A2(G4), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n644), .B2(new_n738), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1348), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n811), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G6), .B(G305), .S(G16), .Z(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT32), .B(G1981), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n738), .A2(G23), .ZN(new_n822));
  INV_X1    g397(.A(G288), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n738), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT33), .B(G1976), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n738), .A2(G22), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G166), .B2(new_n738), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(G1971), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(G1971), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n826), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OR3_X1    g406(.A1(new_n821), .A2(KEYINPUT34), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT34), .B1(new_n821), .B2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n470), .A2(G131), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n490), .A2(G119), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n474), .A2(G107), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  MUX2_X1   g413(.A(G25), .B(new_n838), .S(G29), .Z(new_n839));
  XOR2_X1   g414(.A(KEYINPUT35), .B(G1991), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(G16), .A2(G24), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n628), .A2(new_n629), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(G16), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n841), .B(KEYINPUT94), .C1(G1986), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G1986), .B2(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n832), .A2(new_n833), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n818), .A2(new_n849), .A3(new_n850), .ZN(G311));
  NAND3_X1  g426(.A1(new_n818), .A2(new_n849), .A3(new_n850), .ZN(G150));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n552), .A2(new_n853), .B1(new_n854), .B2(new_n546), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n526), .A2(G67), .A3(new_n541), .A4(new_n542), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n530), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(G860), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n644), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n576), .A2(new_n577), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n531), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n543), .A2(G81), .B1(G43), .B2(new_n547), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n546), .A2(new_n854), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n543), .B2(G93), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n856), .A2(new_n857), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n531), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n864), .A2(new_n865), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n578), .A2(new_n581), .B1(new_n855), .B2(new_n858), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n862), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n875));
  AOI21_X1  g450(.A(G860), .B1(new_n875), .B2(KEYINPUT100), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(KEYINPUT100), .B2(new_n875), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT101), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n860), .B1(new_n877), .B2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(new_n664), .B(new_n488), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n838), .B(KEYINPUT103), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n668), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n490), .A2(G130), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT102), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n470), .A2(G142), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n474), .A2(G118), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n884), .B(new_n890), .Z(new_n891));
  NOR2_X1   g466(.A1(new_n512), .A2(new_n507), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n753), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n778), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n800), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n882), .B1(new_n891), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n897), .B2(new_n891), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n891), .A2(KEYINPUT104), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n896), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n882), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n899), .B(new_n900), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g481(.A(new_n647), .B1(new_n855), .B2(new_n858), .ZN(new_n907));
  OAI21_X1  g482(.A(G299), .B1(new_n636), .B2(new_n643), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n606), .A2(new_n602), .ZN(new_n909));
  AND4_X1   g484(.A1(KEYINPUT83), .A2(new_n526), .A3(new_n542), .A4(new_n541), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT83), .B1(new_n524), .B2(new_n526), .ZN(new_n911));
  OAI21_X1  g486(.A(G65), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n596), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n909), .B1(G651), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n642), .ZN(new_n915));
  OAI21_X1  g490(.A(G66), .B1(new_n910), .B2(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n639), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n917), .B2(G651), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n634), .A2(new_n635), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n908), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n655), .A2(new_n872), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT87), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n654), .B(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(new_n873), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n922), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n923), .A2(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n908), .A2(new_n920), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n908), .B2(new_n920), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n935));
  NOR2_X1   g510(.A1(G166), .A2(new_n823), .ZN(new_n936));
  AOI21_X1  g511(.A(G288), .B1(new_n549), .B2(new_n556), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(G290), .A2(new_n625), .A3(new_n624), .ZN(new_n939));
  NAND2_X1  g514(.A1(G305), .A2(new_n843), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n939), .ZN(new_n942));
  AOI21_X1  g517(.A(G290), .B1(new_n624), .B2(new_n625), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n942), .A2(new_n943), .B1(new_n936), .B2(new_n937), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(KEYINPUT105), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n945), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n935), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n934), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n952), .B(new_n927), .C1(new_n933), .C2(new_n928), .ZN(new_n955));
  OR3_X1    g530(.A1(new_n948), .A2(new_n951), .A3(new_n935), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n907), .B1(new_n957), .B2(new_n647), .ZN(G295));
  OAI21_X1  g533(.A(new_n907), .B1(new_n957), .B2(new_n647), .ZN(G331));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n870), .A2(G286), .A3(new_n871), .ZN(new_n961));
  AOI21_X1  g536(.A(G286), .B1(new_n870), .B2(new_n871), .ZN(new_n962));
  OAI21_X1  g537(.A(G301), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n872), .A2(G168), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n870), .A2(G286), .A3(new_n871), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(G171), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n921), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n930), .A2(KEYINPUT108), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n921), .A2(KEYINPUT41), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n908), .A2(new_n920), .A3(new_n971), .A4(new_n929), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n967), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n968), .B1(new_n974), .B2(KEYINPUT109), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n976), .A3(new_n967), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n945), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT107), .B1(new_n967), .B2(new_n921), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n967), .B1(new_n931), .B2(new_n932), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n963), .A2(new_n966), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n922), .A3(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n979), .A2(new_n980), .A3(new_n945), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n900), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n960), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n984), .A2(new_n985), .A3(new_n900), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n973), .A2(new_n976), .A3(new_n967), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n976), .B1(new_n973), .B2(new_n967), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(new_n968), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n988), .B(KEYINPUT110), .C1(new_n991), .C2(new_n945), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n979), .A2(new_n980), .A3(new_n983), .ZN(new_n993));
  INV_X1    g568(.A(new_n945), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(new_n900), .A3(new_n984), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n987), .A2(new_n992), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n984), .A2(new_n900), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT43), .B1(new_n978), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n999), .B1(new_n988), .B2(new_n995), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT111), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n1002), .A2(KEYINPUT111), .A3(new_n1003), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(G397));
  NOR2_X1   g581(.A1(G290), .A2(G1986), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT112), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(G1986), .B2(G290), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n512), .B2(new_n507), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n471), .A2(new_n480), .A3(G40), .A4(new_n487), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1015), .B(KEYINPUT113), .ZN(new_n1018));
  INV_X1    g593(.A(new_n840), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n838), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n838), .A2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n753), .B(G2067), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT114), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n803), .B2(new_n800), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1016), .A2(G1996), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1025), .A2(new_n1018), .B1(new_n800), .B2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1017), .A2(new_n1022), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n623), .A2(new_n531), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(new_n625), .A3(new_n1030), .A4(new_n616), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n543), .A2(G86), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n617), .B(new_n1032), .C1(new_n623), .C2(new_n531), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1033), .B2(new_n1030), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  AND4_X1   g612(.A1(G40), .A2(new_n471), .A3(new_n480), .A4(new_n487), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1011), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1040), .B1(new_n1044), .B2(G288), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT52), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n823), .B2(G1976), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1046), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1043), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1012), .A2(G1384), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1014), .B1(new_n893), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1384), .B1(new_n509), .B2(new_n513), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(KEYINPUT45), .ZN(new_n1055));
  INV_X1    g630(.A(G1971), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1014), .B1(new_n1039), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2090), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1059), .B(new_n1060), .C1(new_n1054), .C2(new_n1058), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1037), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n549), .A2(G8), .A3(new_n556), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT120), .B1(new_n1051), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT73), .B1(new_n503), .B2(new_n508), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n512), .A2(new_n510), .A3(new_n507), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1068), .B(new_n1052), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1014), .B1(new_n1012), .B2(new_n1011), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1068), .B1(new_n514), .B2(new_n1052), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n741), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT119), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1038), .B1(KEYINPUT50), .B2(new_n1011), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n514), .A2(new_n1010), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(KEYINPUT50), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n734), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n741), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1076), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(G8), .A3(G168), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1049), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1086), .B(new_n1087), .C1(new_n1065), .C2(new_n1062), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1062), .A2(KEYINPUT115), .A3(new_n1065), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1089), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1067), .A2(new_n1085), .A3(new_n1088), .A4(new_n1094), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT50), .B(G1384), .C1(new_n509), .C2(new_n513), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1038), .B1(new_n1039), .B2(new_n1058), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT116), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n514), .A2(new_n1058), .A3(new_n1010), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1014), .B1(KEYINPUT50), .B2(new_n1011), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1102), .A3(new_n1060), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1057), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1037), .B1(new_n1104), .B2(KEYINPUT117), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1106), .A3(new_n1057), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1065), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1062), .A2(KEYINPUT115), .A3(new_n1065), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT115), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1086), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1108), .A2(new_n1111), .A3(new_n1084), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1095), .B1(new_n1112), .B2(KEYINPUT63), .ZN(new_n1113));
  AOI211_X1 g688(.A(G1976), .B(G288), .C1(new_n1036), .C2(new_n1042), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1031), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1040), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1092), .A2(new_n1086), .A3(new_n1093), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT121), .B(G1956), .Z(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(G2072), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1053), .B(new_n1122), .C1(new_n1054), .C2(KEYINPUT45), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n914), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1120), .A2(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(G2067), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1059), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1130));
  INV_X1    g705(.A(G1348), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1127), .B1(new_n644), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1139), .A2(KEYINPUT124), .A3(new_n1123), .A4(new_n1120), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1141), .B1(new_n1137), .B2(new_n1127), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1052), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1038), .B1(new_n892), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1078), .B2(new_n1012), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  AOI22_X1  g727(.A1(new_n1151), .A2(new_n803), .B1(new_n1128), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n582), .B1(KEYINPUT123), .B2(new_n1147), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1148), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1128), .A2(new_n1152), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1055), .B2(G1996), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(KEYINPUT123), .A3(new_n1147), .A4(new_n582), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1145), .A2(new_n1146), .A3(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1132), .A2(KEYINPUT60), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1132), .A2(KEYINPUT60), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(new_n644), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1160), .A2(KEYINPUT125), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1145), .A2(new_n1159), .A3(new_n1146), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1138), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1076), .A2(G168), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT126), .B1(new_n1083), .B2(G8), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT51), .ZN(new_n1170));
  OAI211_X1 g745(.A(G8), .B(new_n1168), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1082), .A2(new_n1080), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1052), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT118), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1081), .B1(new_n1175), .B2(new_n741), .ZN(new_n1176));
  OAI21_X1  g751(.A(G8), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1170), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(G286), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1180), .A2(G8), .A3(new_n1168), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1171), .A2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(G171), .B(KEYINPUT54), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT53), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1055), .B2(G2078), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1130), .A2(new_n807), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n763), .A2(KEYINPUT53), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1187), .B(new_n1188), .C1(new_n1175), .C2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1185), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1014), .B(KEYINPUT127), .Z(new_n1192));
  AOI21_X1  g767(.A(new_n1189), .B1(new_n893), .B2(new_n1052), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1192), .A2(new_n1013), .A3(new_n1193), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1184), .A2(new_n1188), .A3(new_n1187), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1108), .A2(new_n1111), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1183), .A2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1113), .B(new_n1118), .C1(new_n1167), .C2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1171), .A2(new_n1182), .A3(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1202), .A2(G171), .A3(new_n1190), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1200), .B1(new_n1171), .B2(new_n1182), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1028), .B1(new_n1199), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1024), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1018), .B1(new_n1207), .B2(new_n799), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1026), .B(KEYINPUT46), .Z(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT47), .Z(new_n1211));
  NAND2_X1  g786(.A1(new_n1008), .A2(new_n1015), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT48), .ZN(new_n1213));
  AND3_X1   g788(.A1(new_n1213), .A2(new_n1022), .A3(new_n1027), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1027), .A2(new_n1021), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(G2067), .B2(new_n753), .ZN(new_n1216));
  AOI211_X1 g791(.A(new_n1211), .B(new_n1214), .C1(new_n1018), .C2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1206), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g793(.A1(G401), .A2(new_n462), .A3(G227), .A4(G229), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n998), .A2(new_n1220), .A3(new_n905), .ZN(G225));
  INV_X1    g795(.A(G225), .ZN(G308));
endmodule


