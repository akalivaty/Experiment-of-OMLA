//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT72), .B(G237), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT73), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT73), .A2(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G210), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n194), .B(KEYINPUT27), .Z(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G101), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  XOR2_X1   g011(.A(new_n197), .B(KEYINPUT74), .Z(new_n198));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(KEYINPUT11), .B2(G134), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G137), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT11), .A2(G134), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G137), .ZN(new_n211));
  AND4_X1   g025(.A1(new_n205), .A2(new_n209), .A3(new_n211), .A4(new_n207), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n204), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G131), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n216), .B(new_n204), .C1(new_n208), .C2(new_n212), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(KEYINPUT66), .A3(G131), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT0), .A3(G128), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT0), .B(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n218), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT67), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n220), .A2(new_n230), .A3(new_n227), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G143), .ZN(new_n233));
  INV_X1    g047(.A(G143), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n235), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n236), .A2(new_n226), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n229), .A2(new_n231), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n206), .A2(new_n203), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n240), .B(G131), .C1(new_n203), .C2(new_n200), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n217), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n225), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n244));
  INV_X1    g058(.A(G119), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G116), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT68), .A3(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT2), .B(G113), .Z(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n246), .A2(new_n248), .B1(G116), .B2(new_n245), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n252), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(KEYINPUT69), .A3(new_n256), .ZN(new_n257));
  OR3_X1    g071(.A1(new_n255), .A2(KEYINPUT69), .A3(new_n252), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n199), .B1(new_n243), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n243), .A2(new_n260), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n242), .A2(KEYINPUT70), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n217), .A2(new_n239), .A3(new_n264), .A4(new_n241), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n259), .A3(new_n225), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n261), .B(new_n262), .C1(new_n267), .C2(new_n199), .ZN(new_n268));
  INV_X1    g082(.A(new_n267), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n266), .A2(new_n270), .A3(KEYINPUT30), .A4(new_n225), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n225), .A2(KEYINPUT30), .A3(new_n263), .A4(new_n265), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT30), .B1(new_n225), .B2(new_n242), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n269), .B1(new_n275), .B2(new_n260), .ZN(new_n276));
  OAI221_X1 g090(.A(new_n188), .B1(new_n198), .B2(new_n268), .C1(new_n276), .C2(new_n197), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n266), .A2(new_n225), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n260), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n199), .B1(new_n279), .B2(new_n267), .ZN(new_n280));
  INV_X1    g094(.A(new_n261), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n197), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(new_n188), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n187), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n198), .A2(new_n268), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n275), .A2(new_n260), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n197), .A3(new_n267), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n276), .A2(KEYINPUT31), .A3(new_n197), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n287), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT31), .B1(new_n276), .B2(new_n197), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n225), .A2(new_n242), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT71), .B(new_n272), .C1(new_n301), .C2(KEYINPUT30), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n259), .B1(new_n302), .B2(new_n271), .ZN(new_n303));
  NOR4_X1   g117(.A1(new_n303), .A2(new_n292), .A3(new_n283), .A4(new_n269), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n288), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n296), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n298), .A2(new_n299), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n296), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT75), .A3(new_n287), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n286), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n190), .A2(new_n191), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(G221), .A3(G234), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT77), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G137), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n245), .B2(G128), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n226), .A2(KEYINPUT23), .A3(G119), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n317), .B(new_n318), .C1(G119), .C2(new_n226), .ZN(new_n319));
  XNOR2_X1  g133(.A(G119), .B(G128), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT24), .B(G110), .Z(new_n321));
  AOI22_X1  g135(.A1(new_n319), .A2(G110), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G125), .B(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  OR3_X1    g139(.A1(new_n325), .A2(KEYINPUT16), .A3(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(G146), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(G146), .B1(new_n324), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n322), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n319), .A2(G110), .B1(new_n320), .B2(new_n321), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n232), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n315), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G902), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n315), .A2(new_n335), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n339), .B(KEYINPUT25), .Z(new_n340));
  INV_X1    g154(.A(G234), .ZN(new_n341));
  OAI21_X1  g155(.A(G217), .B1(new_n341), .B2(G902), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT76), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n336), .A2(new_n338), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n343), .A2(G902), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT9), .B(G234), .ZN(new_n350));
  OAI21_X1  g164(.A(G221), .B1(new_n350), .B2(G902), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT12), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n218), .A2(new_n219), .ZN(new_n354));
  INV_X1    g168(.A(G104), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(new_n355), .B2(G107), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n357));
  INV_X1    g171(.A(G107), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G104), .ZN(new_n359));
  INV_X1    g173(.A(G101), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(G107), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n356), .A2(new_n359), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n355), .A2(G107), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n358), .A2(G104), .ZN(new_n364));
  OAI21_X1  g178(.A(G101), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n239), .B(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n353), .B1(new_n354), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n366), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n239), .B(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(KEYINPUT12), .A3(new_n219), .A4(new_n218), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n354), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n239), .A2(new_n369), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n356), .A2(new_n359), .A3(new_n361), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G101), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(G101), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n224), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n239), .A2(KEYINPUT10), .A3(new_n369), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n372), .B1(new_n373), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n311), .A2(G227), .ZN(new_n386));
  XOR2_X1   g200(.A(G110), .B(G140), .Z(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n384), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT79), .B1(new_n389), .B2(new_n354), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n373), .A2(new_n391), .A3(new_n384), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n373), .A2(new_n384), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n388), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n385), .A2(new_n388), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G469), .B1(new_n396), .B2(G902), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n372), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n390), .B2(new_n392), .ZN(new_n399));
  INV_X1    g213(.A(new_n388), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G469), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(new_n337), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n352), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G113), .B(G122), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(new_n355), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n323), .B(new_n232), .ZN(new_n408));
  INV_X1    g222(.A(G214), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n234), .B1(new_n192), .B2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n311), .A2(G143), .A3(G214), .A4(new_n189), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(KEYINPUT84), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(KEYINPUT18), .A2(G131), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n408), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n417));
  AOI211_X1 g231(.A(new_n417), .B(new_n216), .C1(new_n410), .C2(new_n411), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(new_n411), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G131), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n410), .A2(new_n216), .A3(new_n411), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n417), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT86), .B1(new_n328), .B2(new_n329), .ZN(new_n426));
  INV_X1    g240(.A(new_n329), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n327), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n426), .B(new_n429), .C1(new_n418), .C2(new_n419), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n407), .B(new_n416), .C1(new_n425), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT88), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT87), .B1(new_n422), .B2(new_n417), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n426), .A2(new_n429), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n420), .A4(new_n424), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n407), .A4(new_n416), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n422), .A2(KEYINPUT85), .A3(new_n423), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n323), .B(KEYINPUT19), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n328), .B1(new_n232), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT85), .B1(new_n422), .B2(new_n423), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n416), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n407), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n448));
  NOR2_X1   g262(.A1(G475), .A2(G902), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n432), .A2(new_n437), .B1(new_n445), .B2(new_n444), .ZN(new_n451));
  INV_X1    g265(.A(new_n449), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT20), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n407), .B1(new_n435), .B2(new_n416), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n432), .B2(new_n437), .ZN(new_n456));
  OAI21_X1  g270(.A(G475), .B1(new_n456), .B2(G902), .ZN(new_n457));
  XNOR2_X1  g271(.A(G128), .B(G143), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n203), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT89), .ZN(new_n460));
  XOR2_X1   g274(.A(G116), .B(G122), .Z(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(G107), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(KEYINPUT13), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n234), .A2(G128), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(G134), .C1(KEYINPUT13), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n458), .B(new_n203), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n247), .A2(KEYINPUT14), .A3(G122), .ZN(new_n468));
  OAI211_X1 g282(.A(G107), .B(new_n468), .C1(new_n461), .C2(KEYINPUT14), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n467), .B(new_n469), .C1(G107), .C2(new_n461), .ZN(new_n470));
  INV_X1    g284(.A(G217), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n350), .A2(new_n471), .A3(G953), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n466), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n472), .B1(new_n466), .B2(new_n470), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n475), .A2(new_n337), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n479));
  OAI21_X1  g293(.A(G478), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n476), .B(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n454), .A2(new_n457), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT5), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n245), .A3(G116), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G113), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n251), .B2(new_n485), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT81), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(new_n369), .A3(new_n490), .A4(new_n256), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n255), .B2(KEYINPUT5), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n252), .A2(new_n249), .A3(new_n250), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n492), .A2(new_n493), .B1(KEYINPUT81), .B2(new_n366), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT8), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n484), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n497), .ZN(new_n499));
  AOI211_X1 g313(.A(KEYINPUT82), .B(new_n499), .C1(new_n491), .C2(new_n494), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n239), .A2(new_n325), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n325), .B2(new_n223), .ZN(new_n503));
  INV_X1    g317(.A(G953), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G224), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(KEYINPUT7), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n257), .A2(new_n258), .A3(new_n379), .A4(new_n381), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n489), .A2(new_n369), .A3(new_n256), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n496), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(KEYINPUT7), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n502), .B(new_n510), .C1(new_n325), .C2(new_n223), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n337), .B1(new_n501), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT83), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n507), .A2(new_n508), .ZN(new_n515));
  INV_X1    g329(.A(new_n496), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT80), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT6), .A4(new_n509), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n503), .B(new_n505), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT83), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n524), .B(new_n337), .C1(new_n501), .C2(new_n512), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n514), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(G210), .B1(G237), .B2(G902), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n514), .A2(new_n527), .A3(new_n523), .A4(new_n525), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(G234), .A2(G237), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n532), .A2(G952), .A3(new_n504), .ZN(new_n533));
  INV_X1    g347(.A(new_n311), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n534), .A2(G902), .A3(new_n532), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT21), .B(G898), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(G214), .B1(G237), .B2(G902), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n405), .A2(new_n483), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n310), .A2(new_n349), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(new_n360), .ZN(G3));
  NAND2_X1  g358(.A1(new_n531), .A2(new_n539), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n531), .A2(new_n547), .A3(new_n539), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n448), .B1(new_n447), .B2(new_n449), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n451), .A2(KEYINPUT20), .A3(new_n452), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n457), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G478), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n337), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n476), .B2(new_n553), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n475), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n557), .B(new_n556), .C1(new_n473), .C2(new_n474), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G478), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n555), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n555), .B2(new_n561), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n552), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n549), .A2(new_n538), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n405), .A2(new_n349), .ZN(new_n569));
  OAI21_X1  g383(.A(G472), .B1(new_n295), .B2(G902), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n308), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n355), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(G6));
  NAND2_X1  g389(.A1(new_n549), .A2(new_n538), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n454), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n450), .A2(new_n453), .A3(KEYINPUT95), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n457), .A2(new_n481), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n571), .A2(new_n576), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT35), .B(G107), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G9));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n315), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(new_n335), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n347), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n344), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n541), .A2(new_n308), .A3(new_n570), .A4(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT37), .B(G110), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G12));
  NAND2_X1  g407(.A1(new_n307), .A2(new_n309), .ZN(new_n594));
  INV_X1    g408(.A(new_n286), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G900), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n533), .B1(new_n535), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n579), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT95), .B1(new_n450), .B2(new_n453), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n581), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT96), .ZN(new_n603));
  INV_X1    g417(.A(new_n590), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n546), .B2(new_n548), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n580), .A2(new_n606), .A3(new_n581), .A4(new_n599), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n596), .A2(new_n404), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT97), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n405), .B1(new_n594), .B2(new_n595), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n608), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G128), .ZN(G30));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n279), .A2(new_n267), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n198), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n291), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n187), .B1(new_n619), .B2(new_n337), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n616), .B1(new_n594), .B2(new_n621), .ZN(new_n622));
  AOI211_X1 g436(.A(KEYINPUT100), .B(new_n620), .C1(new_n307), .C2(new_n309), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT101), .ZN(new_n625));
  INV_X1    g439(.A(new_n552), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n482), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT99), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n531), .B(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n627), .A2(new_n630), .A3(new_n539), .A4(new_n604), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n598), .B(KEYINPUT39), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n404), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT40), .ZN(new_n634));
  OR3_X1    g448(.A1(new_n625), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G143), .ZN(G45));
  NAND3_X1  g450(.A1(new_n552), .A2(new_n565), .A3(new_n599), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n605), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n611), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G146), .ZN(G48));
  NAND2_X1  g455(.A1(new_n401), .A2(new_n337), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n402), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n642), .A2(new_n644), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n645), .A2(new_n646), .A3(new_n352), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n549), .A2(new_n538), .A3(new_n567), .A4(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n310), .A2(new_n648), .A3(new_n349), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT41), .B(G113), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G15));
  INV_X1    g465(.A(new_n539), .ZN(new_n652));
  AOI211_X1 g466(.A(KEYINPUT91), .B(new_n652), .C1(new_n529), .C2(new_n530), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n547), .B1(new_n531), .B2(new_n539), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n647), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n310), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n349), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n580), .A2(new_n657), .A3(new_n538), .A4(new_n581), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G116), .ZN(G18));
  NAND4_X1  g475(.A1(new_n626), .A2(new_n482), .A3(new_n538), .A4(new_n590), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G119), .ZN(G21));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n198), .B1(new_n282), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n280), .A2(KEYINPUT103), .A3(new_n281), .ZN(new_n668));
  OAI22_X1  g482(.A1(new_n300), .A2(new_n304), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n296), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n570), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n349), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n549), .A2(new_n627), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n672), .A2(new_n538), .A3(new_n673), .A4(new_n647), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G122), .ZN(G24));
  NAND3_X1  g489(.A1(new_n570), .A2(new_n670), .A3(new_n590), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n678));
  INV_X1    g492(.A(new_n655), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n677), .A2(new_n678), .A3(new_n638), .A4(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n549), .A2(new_n638), .A3(new_n647), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n681), .B2(new_n676), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  NAND3_X1  g498(.A1(new_n298), .A2(new_n595), .A3(new_n306), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n529), .A2(new_n539), .A3(new_n530), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n404), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n637), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n689), .A3(new_n657), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n685), .A2(new_n689), .A3(new_n692), .A4(new_n657), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n687), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n596), .A2(new_n657), .A3(new_n638), .A4(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n694), .B1(new_n696), .B2(new_n688), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n216), .ZN(G33));
  NOR3_X1   g512(.A1(new_n310), .A2(new_n349), .A3(new_n687), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n603), .A2(new_n607), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G134), .ZN(G36));
  NAND2_X1  g516(.A1(new_n626), .A2(new_n565), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n703), .A2(KEYINPUT43), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(KEYINPUT43), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n570), .A2(new_n308), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n590), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n396), .A2(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n396), .A2(KEYINPUT45), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(G469), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(G469), .A2(G902), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n716), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n403), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n351), .A3(new_n632), .ZN(new_n722));
  INV_X1    g536(.A(new_n686), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n711), .A2(new_n712), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G137), .ZN(G39));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n351), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT47), .ZN(new_n728));
  NOR4_X1   g542(.A1(new_n728), .A2(new_n657), .A3(new_n637), .A4(new_n723), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n310), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT106), .B(G140), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G42));
  NOR4_X1   g546(.A1(new_n703), .A2(new_n349), .A3(new_n652), .A4(new_n352), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n645), .A2(new_n646), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n736), .B(KEYINPUT49), .Z(new_n737));
  NOR3_X1   g551(.A1(new_n735), .A2(new_n630), .A3(new_n737), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n625), .B(new_n738), .C1(new_n734), .C2(new_n733), .ZN(new_n739));
  AOI221_X4 g553(.A(new_n655), .B1(new_n658), .B2(new_n662), .C1(new_n594), .C2(new_n595), .ZN(new_n740));
  INV_X1    g554(.A(new_n674), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n740), .A2(new_n741), .A3(new_n649), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n691), .A2(new_n693), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n310), .A2(new_n349), .A3(new_n637), .A4(new_n687), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n604), .A2(new_n481), .A3(new_n598), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n457), .A3(new_n580), .A4(new_n695), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n638), .A2(new_n695), .ZN(new_n749));
  OAI22_X1  g563(.A1(new_n310), .A2(new_n748), .B1(new_n676), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n700), .B2(new_n699), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  INV_X1    g566(.A(new_n540), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n569), .A2(new_n570), .A3(new_n308), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n566), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n752), .B1(new_n543), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n596), .A2(new_n657), .A3(new_n541), .ZN(new_n757));
  INV_X1    g571(.A(new_n755), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(KEYINPUT108), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n626), .A2(new_n481), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n591), .B1(new_n754), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT109), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n591), .B(new_n763), .C1(new_n754), .C2(new_n760), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n751), .A2(new_n756), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT110), .B1(new_n746), .B2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n756), .A2(new_n759), .A3(new_n765), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n596), .B(new_n679), .C1(new_n659), .C2(new_n663), .ZN(new_n769));
  INV_X1    g583(.A(new_n648), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n596), .A2(new_n657), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n771), .A3(new_n674), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n697), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n768), .A2(new_n773), .A3(new_n774), .A4(new_n751), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n611), .A2(new_n639), .B1(new_n680), .B2(new_n682), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n673), .A2(new_n404), .A3(new_n604), .A4(new_n599), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n622), .B2(new_n623), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n612), .B1(new_n611), .B2(new_n608), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n310), .A2(new_n781), .A3(KEYINPUT97), .A4(new_n405), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n776), .B(new_n779), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n614), .A2(KEYINPUT52), .A3(new_n776), .A4(new_n779), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n767), .A2(new_n775), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n788), .A2(KEYINPUT111), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT111), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT54), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n788), .A2(KEYINPUT112), .A3(new_n789), .ZN(new_n797));
  INV_X1    g611(.A(new_n787), .ZN(new_n798));
  INV_X1    g612(.A(new_n766), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n697), .B2(new_n772), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n742), .A2(new_n745), .A3(KEYINPUT113), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n799), .A2(KEYINPUT53), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n796), .A2(new_n797), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n794), .B1(KEYINPUT54), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n808));
  INV_X1    g622(.A(new_n647), .ZN(new_n809));
  INV_X1    g623(.A(new_n533), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(new_n810), .A3(new_n723), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n625), .A2(new_n657), .A3(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n812), .B(new_n626), .C1(new_n564), .C2(new_n563), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(KEYINPUT115), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(KEYINPUT115), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n706), .A2(new_n349), .A3(new_n810), .A4(new_n671), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n686), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(KEYINPUT114), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n818), .A2(KEYINPUT114), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n736), .A2(new_n352), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n819), .B(new_n820), .C1(new_n728), .C2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n809), .A2(new_n630), .A3(new_n539), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT50), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n707), .A2(new_n811), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n676), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n822), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n808), .B1(new_n816), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n808), .B(new_n828), .C1(new_n814), .C2(new_n815), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n812), .A2(new_n567), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n685), .A2(new_n657), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT48), .Z(new_n834));
  OAI211_X1 g648(.A(new_n504), .B(G952), .C1(KEYINPUT116), .C2(KEYINPUT51), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n817), .B2(new_n679), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n831), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n807), .A2(new_n829), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(G952), .A2(G953), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT117), .Z(new_n840));
  OAI21_X1  g654(.A(new_n739), .B1(new_n838), .B2(new_n840), .ZN(G75));
  NOR2_X1   g655(.A1(new_n311), .A2(G952), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n806), .A2(G902), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(new_n193), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n519), .A2(new_n521), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(new_n522), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT55), .Z(new_n849));
  OAI21_X1  g663(.A(new_n843), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n846), .B2(new_n849), .ZN(G51));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n806), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n716), .B(KEYINPUT57), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n401), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n845), .A2(new_n715), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n842), .B1(new_n855), .B2(new_n856), .ZN(G54));
  NAND4_X1  g671(.A1(new_n806), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n843), .B1(new_n858), .B2(new_n451), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n451), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(KEYINPUT118), .A3(new_n451), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(G60));
  NOR2_X1   g678(.A1(new_n558), .A2(new_n560), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n554), .B(KEYINPUT59), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n843), .B1(new_n853), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n865), .B1(new_n807), .B2(new_n866), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(G63));
  NAND2_X1  g684(.A1(G217), .A2(G902), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT119), .Z(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT60), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n806), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n345), .B(KEYINPUT121), .Z(new_n875));
  AOI21_X1  g689(.A(new_n842), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n877), .A2(new_n806), .A3(new_n588), .A4(new_n873), .ZN(new_n878));
  INV_X1    g692(.A(new_n873), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n804), .B1(new_n792), .B2(new_n795), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n797), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n877), .B1(new_n881), .B2(new_n588), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n876), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(KEYINPUT61), .B(new_n876), .C1(new_n878), .C2(new_n882), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(G66));
  INV_X1    g701(.A(G224), .ZN(new_n888));
  OAI21_X1  g702(.A(G953), .B1(new_n536), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n768), .A2(new_n742), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n891), .B2(new_n534), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n847), .B1(G898), .B2(new_n311), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT122), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n892), .B(new_n894), .ZN(G69));
  XNOR2_X1  g709(.A(new_n275), .B(new_n440), .ZN(new_n896));
  OAI211_X1 g710(.A(G900), .B(new_n534), .C1(new_n896), .C2(G227), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(G227), .B2(new_n896), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n614), .A2(new_n776), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n635), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n902), .B(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n730), .A2(new_n725), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n310), .A2(new_n349), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n633), .B(new_n723), .C1(new_n760), .C2(new_n566), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n896), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n673), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n913), .A2(new_n722), .A3(new_n832), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n906), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n745), .A2(new_n701), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT124), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n901), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n534), .B1(new_n919), .B2(new_n896), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n898), .B1(new_n912), .B2(new_n920), .ZN(G72));
  NAND4_X1  g735(.A1(new_n915), .A2(new_n891), .A3(new_n901), .A4(new_n917), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n187), .A2(new_n337), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n276), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n197), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n843), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n932), .A3(new_n843), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n925), .B1(new_n910), .B2(new_n890), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n197), .A3(new_n927), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT127), .B1(new_n276), .B2(new_n197), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n283), .B2(new_n927), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n276), .A2(KEYINPUT127), .A3(new_n197), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n793), .B(new_n925), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n934), .A2(new_n936), .A3(new_n940), .ZN(G57));
endmodule


