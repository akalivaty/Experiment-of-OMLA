//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT70), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n192), .A2(new_n196), .ZN(new_n197));
  OR3_X1    g011(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT2), .A2(G113), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n192), .A2(new_n196), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(new_n202), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT71), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n206), .A2(new_n209), .B1(new_n202), .B2(new_n207), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G134), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(new_n211), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(G137), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(G131), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT0), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT65), .B1(new_n226), .B2(G143), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(G143), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n225), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n223), .A2(new_n224), .ZN(new_n234));
  XNOR2_X1  g048(.A(G143), .B(G146), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n233), .A2(new_n234), .B1(new_n235), .B2(new_n225), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n228), .B1(new_n229), .B2(G146), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n226), .A2(KEYINPUT65), .A3(G143), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n232), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n224), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n229), .A2(G146), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n232), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n219), .B2(new_n216), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT67), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n247), .B(new_n250), .C1(G131), .C2(new_n221), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n237), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT30), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n210), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n204), .A2(new_n205), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n208), .A2(KEYINPUT71), .ZN(new_n260));
  OAI22_X1  g074(.A1(new_n259), .A2(new_n260), .B1(new_n203), .B2(new_n197), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(new_n252), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G237), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(G210), .ZN(new_n266));
  INV_X1    g080(.A(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n268), .B(new_n269), .Z(new_n270));
  OAI21_X1  g084(.A(new_n188), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n262), .A2(KEYINPUT28), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n270), .B(KEYINPUT72), .Z(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n261), .A2(new_n252), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT73), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n261), .A2(new_n279), .A3(new_n252), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n262), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n274), .B(new_n276), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n270), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT74), .B(new_n284), .C1(new_n258), .C2(new_n262), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n271), .A2(new_n272), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n262), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n277), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n273), .B1(new_n288), .B2(KEYINPUT28), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n284), .A2(new_n272), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n187), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n274), .B1(new_n281), .B2(new_n282), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n275), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n256), .A2(new_n257), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n261), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n287), .A3(new_n270), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT31), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n263), .A2(new_n299), .A3(new_n270), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n294), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n187), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT32), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n301), .A2(new_n305), .A3(new_n187), .A4(new_n302), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n292), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT16), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(G140), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(KEYINPUT75), .A3(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n310), .B1(new_n315), .B2(new_n308), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G146), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n193), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n224), .A2(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT24), .B(G110), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n318), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n326), .B2(G110), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n311), .A2(new_n226), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT76), .Z(new_n330));
  XNOR2_X1  g144(.A(new_n316), .B(new_n226), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n326), .A2(G110), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n320), .A2(new_n321), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT77), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT22), .B(G137), .Z(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n330), .A2(new_n339), .A3(new_n334), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n302), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G217), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(G234), .B2(new_n302), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G902), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n346), .A2(new_n348), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n307), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(KEYINPUT9), .B(G234), .Z(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G221), .B1(new_n354), .B2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n243), .B2(new_n246), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n361));
  OAI211_X1 g175(.A(G104), .B(new_n360), .C1(new_n361), .C2(KEYINPUT3), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT79), .B(new_n363), .C1(new_n364), .C2(G107), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n361), .A2(KEYINPUT3), .B1(new_n364), .B2(G107), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n267), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n360), .A2(G104), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n364), .A2(G107), .ZN(new_n370));
  OAI21_X1  g184(.A(G101), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n246), .B1(new_n241), .B2(new_n235), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n368), .A2(new_n373), .A3(new_n371), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n359), .A2(new_n372), .B1(new_n374), .B2(new_n358), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n366), .A2(new_n367), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n368), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n379), .A3(G101), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n236), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n222), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n375), .A2(new_n381), .A3(new_n382), .A4(KEYINPUT80), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT12), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n374), .B1(new_n372), .B2(new_n247), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n391), .B2(new_n382), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(KEYINPUT12), .A3(new_n222), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n387), .A2(new_n388), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n388), .B1(new_n387), .B2(new_n394), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n265), .A2(G227), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n398), .B(new_n399), .Z(new_n400));
  NOR3_X1   g214(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n387), .B2(new_n400), .ZN(new_n403));
  INV_X1    g217(.A(new_n400), .ZN(new_n404));
  AOI211_X1 g218(.A(KEYINPUT82), .B(new_n404), .C1(new_n385), .C2(new_n386), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n382), .B1(new_n375), .B2(new_n381), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n357), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n403), .ZN(new_n409));
  INV_X1    g223(.A(new_n405), .ZN(new_n410));
  INV_X1    g224(.A(new_n406), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n387), .A2(new_n394), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT81), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n404), .A3(new_n395), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(KEYINPUT83), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n408), .A2(new_n302), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G469), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n387), .A2(new_n400), .A3(new_n394), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n406), .B1(new_n385), .B2(new_n386), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n400), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G469), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT84), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n302), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n422), .A2(KEYINPUT84), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n356), .B1(new_n418), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n264), .A2(new_n265), .A3(G214), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(G143), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n429), .A2(new_n248), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT17), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n429), .B(new_n248), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n331), .B(new_n432), .C1(KEYINPUT17), .C2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G113), .B(G122), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT86), .B(G104), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT18), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n429), .B1(new_n439), .B2(new_n248), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n328), .B1(new_n315), .B2(new_n226), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n440), .B(new_n441), .C1(new_n430), .C2(new_n439), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n434), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n313), .A2(KEYINPUT19), .A3(new_n314), .ZN(new_n444));
  INV_X1    g258(.A(new_n311), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(KEYINPUT19), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n433), .B(new_n317), .C1(G146), .C2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n438), .B1(new_n447), .B2(new_n442), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G475), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n302), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n438), .B1(new_n434), .B2(new_n442), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n302), .B1(new_n443), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G475), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n450), .A4(new_n302), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(G234), .A2(G237), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(G952), .A3(new_n265), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT21), .B(G898), .Z(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(G902), .A3(G953), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n189), .A2(KEYINPUT14), .A3(G122), .ZN(new_n467));
  XOR2_X1   g281(.A(G116), .B(G122), .Z(new_n468));
  OAI211_X1 g282(.A(G107), .B(new_n467), .C1(new_n468), .C2(KEYINPUT14), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n468), .A2(G107), .ZN(new_n472));
  XNOR2_X1  g286(.A(G128), .B(G143), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n212), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(new_n470), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n471), .A2(new_n472), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n468), .A2(G107), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n212), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n212), .B1(new_n473), .B2(KEYINPUT13), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n229), .A2(G128), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(KEYINPUT13), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n353), .A2(G217), .A3(new_n265), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n302), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n487), .B(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n458), .A2(new_n466), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G214), .B1(G237), .B2(G902), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n206), .A2(new_n209), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n197), .B2(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G113), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(new_n372), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n378), .A2(new_n380), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n497), .B1(new_n498), .B2(new_n210), .ZN(new_n499));
  XOR2_X1   g313(.A(G110), .B(G122), .Z(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n500), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n497), .B(new_n502), .C1(new_n498), .C2(new_n210), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n236), .A2(G125), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n247), .A2(new_n309), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n265), .A2(G224), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT85), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n507), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n499), .A2(new_n511), .A3(new_n500), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n504), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n500), .B(KEYINPUT8), .Z(new_n514));
  INV_X1    g328(.A(new_n497), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n372), .B1(new_n493), .B2(new_n496), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n507), .A2(KEYINPUT7), .A3(new_n508), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n508), .A2(KEYINPUT7), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n505), .A2(new_n519), .A3(new_n506), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n503), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n302), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G210), .B1(G237), .B2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n513), .A2(new_n302), .A3(new_n523), .A4(new_n521), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n491), .A2(new_n492), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n352), .A2(new_n427), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(G101), .ZN(G3));
  NAND2_X1  g344(.A1(new_n301), .A2(new_n302), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G472), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n303), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n534), .A2(new_n350), .A3(new_n427), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(new_n536), .A3(new_n526), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n526), .A2(new_n536), .ZN(new_n538));
  INV_X1    g352(.A(new_n466), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n492), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n487), .A2(new_n488), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n487), .A2(KEYINPUT89), .A3(new_n488), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n486), .B(KEYINPUT33), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(G478), .A3(new_n302), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n458), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n540), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n535), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(G104), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(G6));
  INV_X1    g369(.A(new_n458), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n490), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n540), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n535), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G107), .Z(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(G9));
  NAND2_X1  g375(.A1(new_n346), .A2(new_n348), .ZN(new_n562));
  INV_X1    g376(.A(new_n340), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n335), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n349), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n528), .A2(new_n427), .A3(new_n534), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G110), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT91), .B(KEYINPUT37), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(G12));
  INV_X1    g385(.A(new_n307), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n537), .A2(new_n492), .A3(new_n538), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n572), .A2(new_n427), .A3(new_n574), .A4(new_n567), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n464), .A2(G900), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n460), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n575), .A2(new_n557), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(new_n224), .ZN(G30));
  XNOR2_X1  g394(.A(new_n577), .B(KEYINPUT39), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n427), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(KEYINPUT40), .Z(new_n583));
  INV_X1    g397(.A(new_n567), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n458), .A2(new_n490), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n304), .A2(new_n306), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n288), .A2(new_n275), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n297), .A2(G472), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(G472), .A2(G902), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT93), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n585), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n527), .B(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n492), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n583), .A2(new_n584), .A3(new_n592), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G143), .ZN(G45));
  AND3_X1   g412(.A1(new_n572), .A2(new_n427), .A3(new_n567), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT94), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n550), .A2(new_n578), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n574), .A4(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n601), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT94), .B1(new_n575), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G146), .ZN(G48));
  NAND2_X1  g420(.A1(new_n421), .A2(new_n302), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n426), .A2(new_n355), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT95), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n352), .A2(new_n551), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT41), .B(G113), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G15));
  NAND3_X1  g431(.A1(new_n352), .A2(new_n558), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT96), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n352), .A2(new_n620), .A3(new_n558), .A4(new_n614), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G116), .ZN(G18));
  NOR2_X1   g437(.A1(new_n573), .A2(new_n609), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n572), .A2(new_n491), .A3(new_n567), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G119), .ZN(G21));
  OAI211_X1 g440(.A(new_n298), .B(new_n300), .C1(new_n276), .C2(new_n289), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n187), .A3(new_n302), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT97), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n627), .A2(new_n630), .A3(new_n187), .A4(new_n302), .ZN(new_n631));
  AND4_X1   g445(.A1(new_n350), .A2(new_n532), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n540), .B1(new_n611), .B2(new_n613), .ZN(new_n633));
  INV_X1    g447(.A(new_n585), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT98), .A4(new_n634), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G122), .ZN(G24));
  NAND4_X1  g454(.A1(new_n567), .A2(new_n532), .A3(new_n629), .A4(new_n631), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n603), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n624), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G125), .ZN(G27));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n356), .A2(new_n595), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n415), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n414), .A2(KEYINPUT99), .A3(new_n404), .A4(new_n395), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n412), .A2(KEYINPUT100), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n407), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(G469), .B1(new_n654), .B2(G902), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n527), .B1(new_n655), .B2(new_n426), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n352), .A2(new_n646), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n645), .B1(new_n657), .B2(new_n603), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n645), .B(KEYINPUT42), .C1(new_n657), .C2(new_n603), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G131), .ZN(G33));
  NOR2_X1   g477(.A1(new_n557), .A2(new_n578), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n352), .A2(new_n664), .A3(new_n646), .A4(new_n656), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G134), .ZN(G36));
  NOR2_X1   g480(.A1(new_n527), .A2(new_n595), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n458), .A2(new_n548), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT43), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n533), .A3(new_n567), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n670), .A2(new_n673), .A3(new_n671), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n670), .B2(new_n671), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n667), .B(new_n672), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n650), .A2(KEYINPUT45), .A3(new_n651), .A4(new_n653), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n408), .A2(new_n678), .A3(new_n416), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(G469), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n677), .A2(new_n679), .A3(KEYINPUT102), .A4(G469), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n422), .A2(new_n302), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n684), .A2(KEYINPUT46), .A3(new_n686), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n426), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n355), .A3(new_n581), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n691), .A2(KEYINPUT103), .A3(new_n355), .A4(new_n581), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n676), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n215), .ZN(G39));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT46), .B1(new_n684), .B2(new_n686), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n688), .B(new_n685), .C1(new_n682), .C2(new_n683), .ZN(new_n700));
  INV_X1    g514(.A(new_n426), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n698), .B1(new_n702), .B2(new_n356), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n691), .A2(KEYINPUT47), .A3(new_n355), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n572), .A2(new_n350), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n601), .A3(new_n667), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G140), .ZN(G42));
  AND2_X1   g522(.A1(new_n615), .A2(new_n625), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n527), .A2(new_n492), .A3(new_n539), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n490), .B(KEYINPUT106), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n556), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n556), .B2(new_n549), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n535), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n622), .A2(new_n639), .A3(new_n709), .A4(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n599), .A2(new_n577), .A3(new_n667), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n665), .B1(new_n717), .B2(new_n712), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n529), .A2(new_n568), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n579), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n567), .A2(new_n356), .A3(new_n578), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n655), .A2(new_n426), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n592), .A3(new_n574), .A4(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n605), .A2(new_n721), .A3(new_n643), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT52), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n642), .A2(new_n646), .A3(new_n656), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n660), .A2(new_n661), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n579), .B1(new_n602), .B2(new_n604), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n643), .A4(new_n724), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n720), .A2(new_n726), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR4_X1   g549(.A1(new_n728), .A2(new_n716), .A3(new_n719), .A4(new_n718), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT53), .A3(new_n726), .A4(new_n732), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT107), .B(KEYINPUT54), .Z(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n735), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n735), .B2(new_n737), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n352), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n667), .A2(new_n610), .A3(new_n461), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n669), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT48), .Z(new_n750));
  AND3_X1   g564(.A1(new_n632), .A2(new_n461), .A3(new_n669), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n624), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n265), .A2(G952), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n586), .A2(new_n350), .A3(new_n591), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n747), .ZN(new_n755));
  INV_X1    g569(.A(new_n550), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n750), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT112), .ZN(new_n759));
  NOR2_X1   g573(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n751), .A2(new_n667), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT108), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n426), .A2(new_n608), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n355), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n763), .B1(new_n705), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n609), .B1(KEYINPUT109), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n751), .A2(new_n595), .A3(new_n594), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(KEYINPUT109), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n769), .B(new_n770), .Z(new_n771));
  NOR2_X1   g585(.A1(new_n748), .A2(new_n641), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT110), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n755), .A2(new_n556), .A3(new_n548), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n766), .A2(new_n771), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n775), .B(new_n776), .Z(new_n777));
  NAND3_X1  g591(.A1(new_n744), .A2(new_n761), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(G952), .B2(G953), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT105), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT105), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n646), .B(new_n781), .C1(new_n764), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n764), .B2(new_n782), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n754), .A2(new_n594), .A3(new_n668), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n785), .ZN(G75));
  AOI21_X1  g600(.A(new_n302), .B1(new_n735), .B2(new_n737), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(G210), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n504), .A2(new_n512), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT113), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT55), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n510), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n790), .A2(new_n794), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n265), .A2(G952), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(G51));
  NAND2_X1  g612(.A1(new_n735), .A2(new_n737), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n738), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n740), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(new_n685), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n685), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n421), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n787), .A2(new_n682), .A3(new_n683), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n797), .B1(new_n806), .B2(new_n807), .ZN(G54));
  INV_X1    g622(.A(new_n797), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n787), .A2(KEYINPUT58), .A3(G475), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n449), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n449), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT115), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n810), .A2(new_n814), .A3(new_n449), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n811), .B1(new_n813), .B2(new_n815), .ZN(G60));
  NAND2_X1  g630(.A1(G478), .A2(G902), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT59), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n741), .B2(new_n743), .ZN(new_n819));
  INV_X1    g633(.A(new_n546), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n797), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n739), .B1(new_n735), .B2(new_n737), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n546), .B(new_n818), .C1(new_n741), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n801), .A2(KEYINPUT116), .A3(new_n546), .A4(new_n818), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(G63));
  NAND2_X1  g641(.A1(G217), .A2(G902), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT60), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n735), .B2(new_n737), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n797), .B1(new_n830), .B2(new_n565), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n832));
  OAI221_X1 g646(.A(new_n831), .B1(KEYINPUT117), .B2(new_n832), .C1(new_n343), .C2(new_n830), .ZN(new_n833));
  INV_X1    g647(.A(new_n829), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n799), .A2(new_n565), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(KEYINPUT117), .A3(new_n809), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n809), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n830), .A2(new_n343), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n836), .B(KEYINPUT61), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n833), .A2(new_n839), .ZN(G66));
  OAI21_X1  g654(.A(new_n265), .B1(new_n716), .B2(new_n719), .ZN(new_n841));
  INV_X1    g655(.A(G224), .ZN(new_n842));
  OAI21_X1  g656(.A(G953), .B1(new_n463), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(KEYINPUT118), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(KEYINPUT118), .B2(new_n841), .ZN(new_n845));
  INV_X1    g659(.A(G898), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n792), .B1(new_n846), .B2(G953), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n845), .B(new_n847), .ZN(G69));
  NOR2_X1   g662(.A1(new_n573), .A2(new_n585), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n699), .A2(new_n700), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n356), .B1(new_n850), .B2(new_n426), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT103), .B1(new_n851), .B2(new_n581), .ZN(new_n852));
  INV_X1    g666(.A(new_n695), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n352), .B(new_n849), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n707), .A3(new_n662), .A4(new_n665), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n730), .A2(new_n643), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT122), .B1(new_n696), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n676), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n852), .B2(new_n853), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n862));
  INV_X1    g676(.A(new_n858), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n856), .A2(new_n857), .A3(new_n859), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n859), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT123), .B1(new_n866), .B2(new_n855), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n867), .A3(new_n265), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n295), .B(KEYINPUT119), .Z(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n446), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(G900), .B2(G953), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n870), .B(KEYINPUT120), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n707), .A2(new_n861), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n730), .A2(new_n597), .A3(new_n643), .ZN(new_n876));
  AND2_X1   g690(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n877));
  NOR2_X1   g691(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n745), .A2(new_n582), .A3(new_n713), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n875), .B(new_n880), .C1(new_n667), .C2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n874), .B1(new_n882), .B2(G953), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n873), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n874), .A2(KEYINPUT124), .ZN(new_n885));
  NAND2_X1  g699(.A1(G227), .A2(G900), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(G953), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n873), .A2(new_n883), .A3(new_n887), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(G72));
  NAND3_X1  g705(.A1(new_n271), .A2(new_n297), .A3(new_n285), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n589), .B(KEYINPUT63), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT126), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n799), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n809), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n716), .A2(new_n719), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n263), .B(KEYINPUT125), .Z(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n882), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n899), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n865), .B2(new_n867), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n893), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n899), .B(new_n284), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n897), .B1(new_n903), .B2(new_n904), .ZN(G57));
endmodule


