//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT64), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G127gat), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G134gat), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n209), .A2(new_n210), .A3(new_n212), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n214), .ZN(new_n216));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(G176gat), .ZN(new_n226));
  OR2_X1    g025(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT24), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT24), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(G183gat), .A3(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n225), .B(new_n229), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(new_n226), .B2(new_n220), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n225), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT66), .B(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n234), .B1(new_n242), .B2(G183gat), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n237), .A2(new_n238), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT26), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n230), .B(new_n245), .C1(new_n247), .C2(new_n223), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT27), .B(G183gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT28), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n241), .A2(new_n249), .A3(KEYINPUT28), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n219), .B1(new_n244), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n243), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n225), .A2(new_n229), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n236), .B1(new_n231), .B2(new_n233), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n238), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n254), .ZN(new_n261));
  INV_X1    g060(.A(new_n219), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n204), .B1(new_n255), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT32), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G15gat), .B(G43gat), .Z(new_n267));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n244), .A2(new_n219), .A3(new_n254), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n262), .B1(new_n260), .B2(new_n261), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n203), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT33), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n255), .A2(new_n263), .A3(new_n204), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT34), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT34), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n255), .A2(new_n263), .A3(new_n278), .A4(new_n204), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n269), .B1(new_n264), .B2(KEYINPUT33), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n277), .A3(new_n279), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n266), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n283), .A3(new_n266), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT36), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT36), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n281), .A2(new_n283), .A3(new_n266), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(new_n284), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n292));
  XNOR2_X1  g091(.A(G78gat), .B(G106gat), .ZN(new_n293));
  INV_X1    g092(.A(G50gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G228gat), .A2(G233gat), .ZN(new_n296));
  XOR2_X1   g095(.A(G155gat), .B(G162gat), .Z(new_n297));
  INV_X1    g096(.A(G141gat), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(KEYINPUT2), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT68), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n300), .A2(new_n307), .A3(new_n301), .ZN(new_n308));
  XNOR2_X1  g107(.A(G155gat), .B(G162gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n311));
  INV_X1    g110(.A(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT69), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n311), .B1(new_n316), .B2(G155gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n303), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(G211gat), .A2(G218gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G197gat), .A2(G204gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(G197gat), .A2(G204gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n325), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT29), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n318), .B1(new_n331), .B2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(new_n303), .C1(new_n310), .C2(new_n317), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT67), .B(new_n321), .C1(new_n324), .C2(new_n325), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n326), .A2(new_n330), .A3(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n334), .A2(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n339), .B2(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n335), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n336), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n341), .A2(KEYINPUT73), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n296), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G22gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(KEYINPUT74), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n334), .A2(new_n347), .A3(new_n335), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n342), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n338), .A2(new_n336), .A3(new_n335), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n333), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n296), .B1(new_n351), .B2(new_n318), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n344), .A2(new_n345), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n345), .B1(new_n344), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n295), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n296), .ZN(new_n357));
  INV_X1    g156(.A(new_n332), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n342), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT73), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n339), .A2(KEYINPUT73), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n349), .A2(new_n352), .ZN(new_n364));
  OAI21_X1  g163(.A(G22gat), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n295), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n344), .A2(new_n345), .A3(new_n353), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n292), .B1(new_n356), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n356), .A2(new_n368), .A3(new_n292), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G1gat), .B(G29gat), .Z(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT0), .ZN(new_n374));
  XNOR2_X1  g173(.A(G57gat), .B(G85gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n304), .A2(new_n305), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n309), .B1(new_n311), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT69), .B(G162gat), .ZN(new_n383));
  INV_X1    g182(.A(G155gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT2), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n381), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n262), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n318), .A2(new_n219), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n379), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT5), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n385), .A2(new_n309), .A3(new_n308), .A4(new_n306), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n262), .A2(new_n391), .A3(KEYINPUT4), .A4(new_n303), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n318), .B2(new_n219), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT70), .B1(new_n386), .B2(new_n333), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT70), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n318), .A2(new_n397), .A3(KEYINPUT3), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n334), .A2(new_n219), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n390), .B1(new_n401), .B2(new_n378), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n318), .A2(new_n397), .A3(KEYINPUT3), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n318), .B2(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n392), .A2(new_n394), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .A4(new_n378), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n377), .B1(new_n402), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT71), .B(KEYINPUT6), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(new_n406), .A3(new_n378), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n318), .B(new_n219), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n407), .B1(new_n415), .B2(new_n379), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n376), .A3(new_n408), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n418), .A2(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n410), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  INV_X1    g223(.A(G226gat), .ZN(new_n425));
  INV_X1    g224(.A(G233gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n260), .A2(new_n261), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n335), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n427), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n342), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  INV_X1    g232(.A(new_n342), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n433), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n421), .B(new_n424), .C1(new_n432), .C2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n424), .B1(new_n432), .B2(new_n435), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n430), .A2(new_n342), .A3(new_n431), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n434), .B1(new_n433), .B2(new_n429), .ZN(new_n439));
  INV_X1    g238(.A(new_n424), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT30), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n413), .A2(new_n420), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n291), .B1(new_n372), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT75), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n376), .B(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n417), .B2(new_n408), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT76), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI211_X1 g248(.A(KEYINPUT76), .B(new_n446), .C1(new_n417), .C2(new_n408), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n419), .B(KEYINPUT77), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n413), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT77), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n449), .A2(new_n450), .ZN(new_n455));
  INV_X1    g254(.A(new_n419), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT37), .B1(new_n432), .B2(new_n435), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n438), .A2(new_n439), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n424), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT38), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n437), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n453), .A2(new_n457), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n356), .A2(new_n368), .A3(new_n292), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(new_n369), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n405), .A2(new_n406), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n379), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(KEYINPUT39), .C1(new_n379), .C2(new_n415), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n472), .B(new_n446), .C1(KEYINPUT39), .C2(new_n471), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT40), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n442), .A2(new_n436), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(new_n455), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n469), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n444), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT78), .B(KEYINPUT35), .ZN(new_n480));
  INV_X1    g279(.A(new_n446), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n402), .B2(new_n409), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT76), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n447), .A2(new_n448), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT77), .B1(new_n485), .B2(new_n419), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n480), .B1(new_n452), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n289), .A2(new_n284), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(new_n475), .C1(new_n468), .C2(new_n369), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n479), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n489), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n457), .A2(new_n413), .A3(new_n451), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT79), .A4(new_n480), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n372), .A2(new_n443), .A3(new_n488), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n478), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n498));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(G197gat), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT11), .B(G169gat), .Z(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT81), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n502), .A2(new_n503), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT81), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n503), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n511), .B(KEYINPUT13), .Z(new_n512));
  OAI21_X1  g311(.A(KEYINPUT85), .B1(new_n294), .B2(G43gat), .ZN(new_n513));
  INV_X1    g312(.A(G43gat), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT84), .B1(new_n514), .B2(G50gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(new_n514), .A3(G50gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(new_n294), .A3(G43gat), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n513), .A2(new_n515), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT83), .B(KEYINPUT15), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT14), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(new_n523), .A3(new_n524), .A4(new_n525), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT15), .B1(new_n514), .B2(G50gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n294), .A2(G43gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n522), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(KEYINPUT82), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT82), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n539), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n540), .A3(new_n526), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n532), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n533), .A2(new_n534), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G1gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT16), .ZN(new_n547));
  INV_X1    g346(.A(G15gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G22gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n345), .A2(G15gat), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(G1gat), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g351(.A(G8gat), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n546), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n556));
  INV_X1    g355(.A(G8gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n545), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n535), .B1(new_n520), .B2(new_n521), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n561), .A2(new_n531), .B1(new_n542), .B2(new_n543), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n553), .A2(new_n558), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n512), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n545), .A2(KEYINPUT17), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n559), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT18), .B(new_n511), .C1(new_n562), .C2(new_n563), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n565), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n537), .A2(new_n567), .A3(new_n544), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n567), .B1(new_n537), .B2(new_n544), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n563), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n545), .A2(new_n559), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n511), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n571), .A2(KEYINPUT87), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n511), .A2(KEYINPUT18), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n545), .B2(new_n559), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT87), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n565), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n510), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n581), .A2(new_n504), .A3(new_n565), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n572), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n498), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n566), .A2(new_n568), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n570), .B1(new_n590), .B2(new_n563), .ZN(new_n591));
  INV_X1    g390(.A(new_n512), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n562), .A2(new_n563), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n592), .B1(new_n576), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT87), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n586), .A3(new_n583), .ZN(new_n596));
  INV_X1    g395(.A(new_n510), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(KEYINPUT88), .A3(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n589), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n497), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT92), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n607), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(G57gat), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n612), .A2(G64gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(G64gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT9), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G71gat), .A2(G78gat), .ZN(new_n616));
  INV_X1    g415(.A(G71gat), .ZN(new_n617));
  INV_X1    g416(.A(G78gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT89), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT89), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(G71gat), .B2(G78gat), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n615), .A2(new_n616), .A3(new_n619), .A4(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT91), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT9), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n612), .A2(KEYINPUT90), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT90), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(G57gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n627), .A3(G64gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n614), .ZN(new_n629));
  AOI221_X4 g428(.A(new_n623), .B1(new_n624), .B2(new_n616), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n624), .A2(new_n616), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT91), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n622), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT21), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n634), .B2(new_n636), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n611), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n637), .A3(new_n610), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n634), .A2(KEYINPUT94), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n644), .B(new_n622), .C1(new_n630), .C2(new_n633), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(KEYINPUT21), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n563), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n640), .B2(new_n642), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n604), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n640), .A2(new_n642), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(new_n603), .A3(new_n648), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(G85gat), .ZN(new_n657));
  INV_X1    g456(.A(G92gat), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT7), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT7), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(G85gat), .A3(G92gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G99gat), .B(G106gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(G99gat), .A2(G106gat), .ZN(new_n664));
  AOI22_X1  g463(.A1(KEYINPUT8), .A2(new_n664), .B1(new_n657), .B2(new_n658), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n662), .B2(new_n665), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n634), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n668), .B(new_n622), .C1(new_n633), .C2(new_n630), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n666), .A2(new_n667), .A3(new_n672), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n643), .A2(new_n645), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(G230gat), .A2(G233gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n670), .A2(new_n671), .ZN(new_n679));
  INV_X1    g478(.A(new_n677), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(G120gat), .B(G148gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(G176gat), .B(G204gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n683), .B(new_n684), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n678), .A2(new_n681), .A3(new_n685), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n669), .B1(new_n573), .B2(new_n574), .ZN(new_n690));
  NAND2_X1  g489(.A1(G232gat), .A2(G233gat), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT95), .Z(new_n692));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n545), .B2(new_n668), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(G190gat), .B(G218gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT96), .ZN(new_n699));
  INV_X1    g498(.A(new_n697), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n690), .A2(new_n700), .A3(new_n695), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n692), .A2(new_n693), .ZN(new_n702));
  XOR2_X1   g501(.A(G134gat), .B(G162gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(KEYINPUT96), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n707), .A2(new_n704), .B1(new_n698), .B2(new_n701), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n656), .A2(new_n689), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n602), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n413), .A2(new_n420), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n546), .ZN(G1324gat));
  INV_X1    g513(.A(new_n475), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT16), .B(G8gat), .Z(new_n716));
  NAND4_X1  g515(.A1(new_n602), .A2(new_n715), .A3(new_n710), .A4(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G8gat), .B1(new_n711), .B2(new_n475), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n717), .ZN(new_n719));
  MUX2_X1   g518(.A(new_n717), .B(new_n719), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g519(.A(KEYINPUT98), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT97), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n287), .A2(new_n290), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n287), .B2(new_n290), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n725), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(KEYINPUT98), .A3(new_n723), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G15gat), .B1(new_n711), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n488), .A2(new_n548), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n711), .B2(new_n732), .ZN(G1326gat));
  NAND3_X1  g532(.A1(new_n602), .A2(new_n469), .A3(new_n710), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT99), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(KEYINPUT99), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT43), .B(G22gat), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n736), .B2(new_n737), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(G1327gat));
  NOR2_X1   g540(.A1(new_n584), .A2(new_n588), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n656), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n744), .A3(new_n689), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT44), .B1(new_n497), .B2(new_n709), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT101), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n706), .B2(new_n708), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n707), .A2(new_n704), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n698), .A2(new_n701), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(KEYINPUT101), .A3(new_n705), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n467), .A2(new_n477), .ZN(new_n758));
  INV_X1    g557(.A(new_n712), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n469), .B1(new_n759), .B2(new_n715), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n724), .A2(new_n725), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n490), .A2(new_n493), .B1(new_n495), .B2(KEYINPUT35), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n745), .B1(new_n746), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G29gat), .B1(new_n767), .B2(new_n712), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n769));
  INV_X1    g568(.A(new_n709), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n744), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n689), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n602), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n524), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n769), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n774), .A2(new_n769), .A3(new_n775), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n768), .A2(new_n776), .A3(new_n777), .ZN(G1328gat));
  OAI21_X1  g577(.A(G36gat), .B1(new_n767), .B2(new_n475), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n715), .A2(new_n525), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT46), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n780), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(G1329gat));
  OAI21_X1  g582(.A(G43gat), .B1(new_n767), .B2(new_n761), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n602), .A2(new_n514), .A3(new_n488), .A4(new_n773), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G43gat), .B1(new_n767), .B2(new_n730), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n785), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n788), .B2(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g588(.A(new_n294), .B1(new_n766), .B2(new_n469), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT48), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n469), .A2(new_n294), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n791), .A2(KEYINPUT102), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n792), .A2(KEYINPUT102), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n792), .A2(KEYINPUT102), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n797), .B(new_n798), .C1(new_n790), .C2(new_n794), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n796), .A2(new_n799), .ZN(G1331gat));
  INV_X1    g599(.A(new_n764), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n762), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n743), .A2(new_n689), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n709), .A3(new_n656), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT103), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT103), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(new_n808), .A3(new_n805), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n759), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT104), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n625), .A2(new_n627), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT104), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n807), .A2(new_n813), .A3(new_n759), .A4(new_n809), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n811), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(G1332gat));
  AOI21_X1  g616(.A(new_n475), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n807), .A2(new_n809), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT105), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n819), .B(new_n821), .ZN(G1333gat));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n729), .A3(new_n809), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G71gat), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n617), .A3(new_n488), .A4(new_n809), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(KEYINPUT50), .A3(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1334gat));
  NAND3_X1  g629(.A1(new_n807), .A2(new_n469), .A3(new_n809), .ZN(new_n831));
  XOR2_X1   g630(.A(KEYINPUT106), .B(G78gat), .Z(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(G1335gat));
  NAND2_X1  g632(.A1(new_n803), .A2(new_n744), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT107), .Z(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n746), .B2(new_n765), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n759), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G85gat), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n771), .A2(new_n743), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n802), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT51), .B(new_n841), .C1(new_n763), .C2(new_n764), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n759), .A2(new_n657), .A3(new_n772), .ZN(new_n846));
  OAI22_X1  g645(.A1(new_n839), .A2(new_n840), .B1(new_n845), .B2(new_n846), .ZN(G1336gat));
  INV_X1    g646(.A(KEYINPUT109), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n475), .B(new_n835), .C1(new_n746), .C2(new_n765), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n658), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n475), .A2(new_n689), .A3(G92gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n842), .B2(new_n844), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n849), .B2(new_n658), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI221_X1 g654(.A(new_n852), .B1(new_n848), .B2(KEYINPUT52), .C1(new_n849), .C2(new_n658), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(G1337gat));
  INV_X1    g656(.A(G99gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n488), .A2(new_n772), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n845), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n836), .B2(new_n729), .ZN(new_n861));
  OR3_X1    g660(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT110), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT110), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1338gat));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n372), .B(new_n835), .C1(new_n746), .C2(new_n765), .ZN(new_n866));
  INV_X1    g665(.A(G106gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n372), .A2(G106gat), .A3(new_n689), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n842), .B2(new_n844), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n866), .B2(new_n867), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n868), .A2(new_n871), .A3(KEYINPUT53), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n873));
  OAI221_X1 g672(.A(new_n870), .B1(new_n865), .B2(new_n873), .C1(new_n866), .C2(new_n867), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1339gat));
  NAND3_X1  g674(.A1(new_n656), .A2(new_n689), .A3(new_n709), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n876), .A2(new_n743), .A3(KEYINPUT112), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT112), .B1(new_n876), .B2(new_n743), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n673), .A2(new_n675), .A3(new_n680), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n678), .A2(KEYINPUT54), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n680), .B1(new_n673), .B2(new_n675), .ZN(new_n883));
  XNOR2_X1  g682(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n685), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(KEYINPUT55), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n688), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n576), .A2(new_n593), .A3(new_n592), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n569), .A2(new_n564), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n511), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n502), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n587), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT55), .B1(new_n882), .B2(new_n885), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n887), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n748), .A2(new_n752), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n880), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n891), .A2(new_n587), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n885), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT55), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n897), .A2(new_n900), .A3(new_n688), .A4(new_n886), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n753), .A3(KEYINPUT114), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n689), .A2(new_n892), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n893), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n743), .B2(new_n904), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n896), .A2(new_n902), .B1(new_n905), .B2(new_n895), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n879), .B1(new_n906), .B2(new_n744), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n712), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n491), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT115), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n207), .A3(new_n743), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n907), .A2(new_n469), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(new_n759), .A3(new_n475), .A4(new_n488), .ZN(new_n913));
  OAI21_X1  g712(.A(G113gat), .B1(new_n913), .B2(new_n601), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT116), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n911), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1340gat));
  NAND3_X1  g718(.A1(new_n910), .A2(new_n205), .A3(new_n772), .ZN(new_n920));
  OAI21_X1  g719(.A(G120gat), .B1(new_n913), .B2(new_n689), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1341gat));
  INV_X1    g721(.A(new_n909), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n213), .A3(new_n656), .ZN(new_n924));
  OAI21_X1  g723(.A(G127gat), .B1(new_n913), .B2(new_n744), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1342gat));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n211), .A3(new_n770), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT56), .ZN(new_n928));
  OAI21_X1  g727(.A(G134gat), .B1(new_n913), .B2(new_n709), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(KEYINPUT56), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(G1343gat));
  NOR4_X1   g730(.A1(new_n724), .A2(new_n725), .A3(new_n712), .A4(new_n715), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n469), .A2(KEYINPUT57), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n896), .A2(new_n902), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT88), .B1(new_n598), .B2(new_n587), .ZN(new_n935));
  AOI221_X4 g734(.A(new_n498), .B1(new_n586), .B2(new_n585), .C1(new_n596), .C2(new_n597), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n904), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n903), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT117), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n709), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n903), .B1(new_n600), .B2(new_n904), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT117), .B1(new_n942), .B2(new_n770), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n934), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n744), .ZN(new_n945));
  INV_X1    g744(.A(new_n879), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n933), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n906), .A2(new_n744), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n946), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT57), .B1(new_n949), .B2(new_n469), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n932), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT118), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT57), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n907), .B2(new_n372), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n879), .B1(new_n944), .B2(new_n744), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n933), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n957), .A3(new_n932), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n952), .A2(new_n743), .A3(new_n958), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n729), .A2(new_n372), .A3(new_n715), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n908), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n601), .A2(G141gat), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n959), .A2(G141gat), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT58), .ZN(new_n964));
  OAI21_X1  g763(.A(G141gat), .B1(new_n951), .B2(new_n601), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT58), .B1(new_n961), .B2(new_n962), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT119), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n967), .B1(new_n965), .B2(new_n966), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n963), .A2(new_n964), .B1(new_n968), .B2(new_n969), .ZN(G1344gat));
  INV_X1    g769(.A(new_n958), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n957), .B1(new_n956), .B2(new_n932), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n971), .A2(new_n972), .A3(new_n689), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n299), .A2(KEYINPUT59), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n770), .B1(new_n937), .B2(new_n938), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n901), .A2(new_n709), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n744), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n601), .A2(KEYINPUT121), .A3(new_n710), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n980), .B1(new_n600), .B2(new_n876), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n372), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n975), .B1(new_n983), .B2(KEYINPUT57), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n979), .A2(new_n981), .ZN(new_n985));
  INV_X1    g784(.A(new_n977), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n986), .B1(new_n942), .B2(new_n770), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n985), .B1(new_n987), .B2(new_n744), .ZN(new_n988));
  OAI211_X1 g787(.A(KEYINPUT122), .B(new_n953), .C1(new_n988), .C2(new_n372), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n949), .A2(KEYINPUT57), .A3(new_n469), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n984), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n932), .A2(new_n772), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n299), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g792(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n994));
  OAI22_X1  g793(.A1(new_n973), .A2(new_n974), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n961), .A2(new_n299), .A3(new_n772), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1345gat));
  NAND3_X1  g796(.A1(new_n961), .A2(new_n384), .A3(new_n656), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n971), .A2(new_n972), .A3(new_n744), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n999), .B2(new_n384), .ZN(G1346gat));
  AOI21_X1  g799(.A(new_n316), .B1(new_n961), .B2(new_n770), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n971), .A2(new_n972), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n753), .A2(new_n383), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(G1347gat));
  NOR2_X1   g803(.A1(new_n907), .A2(new_n759), .ZN(new_n1005));
  AND4_X1   g804(.A1(new_n372), .A2(new_n1005), .A3(new_n715), .A4(new_n488), .ZN(new_n1006));
  NAND4_X1  g805(.A1(new_n1006), .A2(new_n227), .A3(new_n228), .A4(new_n743), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n759), .A2(new_n475), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n1008), .A2(new_n488), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n912), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g809(.A(G169gat), .B1(new_n1010), .B2(new_n601), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1007), .A2(new_n1011), .ZN(G1348gat));
  NAND3_X1  g811(.A1(new_n1006), .A2(new_n221), .A3(new_n772), .ZN(new_n1013));
  OAI21_X1  g812(.A(G176gat), .B1(new_n1010), .B2(new_n689), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(G1349gat));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n912), .A2(new_n656), .A3(new_n1009), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n1016), .B1(new_n1017), .B2(G183gat), .ZN(new_n1018));
  AND2_X1   g817(.A1(new_n656), .A2(new_n249), .ZN(new_n1019));
  AND3_X1   g818(.A1(new_n1006), .A2(KEYINPUT123), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g819(.A(KEYINPUT123), .B1(new_n1006), .B2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1022), .A2(KEYINPUT60), .ZN(new_n1023));
  INV_X1    g822(.A(KEYINPUT60), .ZN(new_n1024));
  OAI211_X1 g823(.A(new_n1024), .B(new_n1018), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1023), .A2(new_n1025), .ZN(G1350gat));
  OAI21_X1  g825(.A(G190gat), .B1(new_n1010), .B2(new_n709), .ZN(new_n1027));
  XNOR2_X1  g826(.A(new_n1027), .B(KEYINPUT61), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1006), .A2(new_n241), .A3(new_n895), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1028), .A2(new_n1029), .ZN(G1351gat));
  NOR3_X1   g829(.A1(new_n729), .A2(new_n372), .A3(new_n475), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1005), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g831(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g832(.A(G197gat), .B1(new_n1033), .B2(new_n743), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n726), .A2(new_n728), .A3(new_n1008), .ZN(new_n1035));
  XOR2_X1   g834(.A(new_n1035), .B(KEYINPUT125), .Z(new_n1036));
  AND2_X1   g835(.A1(new_n991), .A2(new_n1036), .ZN(new_n1037));
  AND2_X1   g836(.A1(new_n600), .A2(G197gat), .ZN(new_n1038));
  AOI21_X1  g837(.A(new_n1034), .B1(new_n1037), .B2(new_n1038), .ZN(G1352gat));
  NOR3_X1   g838(.A1(new_n1032), .A2(G204gat), .A3(new_n689), .ZN(new_n1040));
  XNOR2_X1  g839(.A(new_n1040), .B(KEYINPUT62), .ZN(new_n1041));
  AND2_X1   g840(.A1(new_n1037), .A2(new_n772), .ZN(new_n1042));
  INV_X1    g841(.A(G204gat), .ZN(new_n1043));
  OAI21_X1  g842(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(G1353gat));
  NAND3_X1  g843(.A1(new_n991), .A2(new_n656), .A3(new_n1036), .ZN(new_n1045));
  INV_X1    g844(.A(KEYINPUT63), .ZN(new_n1046));
  NAND3_X1  g845(.A1(new_n1045), .A2(new_n1046), .A3(G211gat), .ZN(new_n1047));
  NOR2_X1   g846(.A1(new_n744), .A2(G211gat), .ZN(new_n1048));
  NAND3_X1  g847(.A1(new_n1005), .A2(new_n1031), .A3(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g848(.A(new_n1049), .B(KEYINPUT126), .ZN(new_n1050));
  NAND2_X1  g849(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g850(.A(new_n1046), .B1(new_n1045), .B2(G211gat), .ZN(new_n1052));
  OAI21_X1  g851(.A(KEYINPUT127), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g852(.A1(new_n1045), .A2(G211gat), .ZN(new_n1054));
  NAND2_X1  g853(.A1(new_n1054), .A2(KEYINPUT63), .ZN(new_n1055));
  INV_X1    g854(.A(KEYINPUT127), .ZN(new_n1056));
  NAND4_X1  g855(.A1(new_n1055), .A2(new_n1056), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1057));
  NAND2_X1  g856(.A1(new_n1053), .A2(new_n1057), .ZN(G1354gat));
  INV_X1    g857(.A(G218gat), .ZN(new_n1059));
  NAND3_X1  g858(.A1(new_n1033), .A2(new_n1059), .A3(new_n895), .ZN(new_n1060));
  AND2_X1   g859(.A1(new_n1037), .A2(new_n770), .ZN(new_n1061));
  OAI21_X1  g860(.A(new_n1060), .B1(new_n1061), .B2(new_n1059), .ZN(G1355gat));
endmodule


