

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761;

  XNOR2_X1 U373 ( .A(n727), .B(n728), .ZN(n349) );
  OR2_X1 U374 ( .A1(n704), .A2(n587), .ZN(n461) );
  BUF_X1 U375 ( .A(n681), .Z(n418) );
  XNOR2_X1 U376 ( .A(n472), .B(KEYINPUT66), .ZN(n528) );
  INV_X1 U377 ( .A(KEYINPUT4), .ZN(n472) );
  NOR2_X2 U378 ( .A1(G902), .A2(n649), .ZN(n545) );
  XNOR2_X2 U379 ( .A(n471), .B(n397), .ZN(n745) );
  NOR2_X1 U380 ( .A1(n349), .A2(n731), .ZN(G63) );
  XNOR2_X1 U381 ( .A(n444), .B(n526), .ZN(n602) );
  NOR2_X1 U382 ( .A1(n591), .A2(n590), .ZN(n660) );
  XNOR2_X2 U383 ( .A(n745), .B(n530), .ZN(n387) );
  XNOR2_X2 U384 ( .A(n633), .B(KEYINPUT86), .ZN(n661) );
  NOR2_X2 U385 ( .A1(n443), .A2(n632), .ZN(n633) );
  INV_X1 U386 ( .A(n385), .ZN(n384) );
  OR2_X1 U387 ( .A1(n483), .A2(KEYINPUT44), .ZN(n422) );
  XNOR2_X1 U388 ( .A(n392), .B(n365), .ZN(n758) );
  XNOR2_X1 U389 ( .A(n469), .B(n468), .ZN(n757) );
  NAND2_X1 U390 ( .A1(n396), .A2(n393), .ZN(n587) );
  XNOR2_X1 U391 ( .A(n415), .B(KEYINPUT82), .ZN(n629) );
  AND2_X1 U392 ( .A1(n431), .A2(n350), .ZN(n440) );
  AND2_X1 U393 ( .A1(n675), .A2(n674), .ZN(n586) );
  XNOR2_X1 U394 ( .A(n626), .B(KEYINPUT38), .ZN(n689) );
  XNOR2_X1 U395 ( .A(n411), .B(n732), .ZN(n391) );
  XNOR2_X1 U396 ( .A(n428), .B(n427), .ZN(n411) );
  OR2_X1 U397 ( .A1(n730), .A2(G902), .ZN(n444) );
  XNOR2_X1 U398 ( .A(n527), .B(G134), .ZN(n397) );
  XNOR2_X2 U399 ( .A(n624), .B(n459), .ZN(n609) );
  NOR2_X2 U400 ( .A1(n678), .A2(n677), .ZN(n675) );
  INV_X1 U401 ( .A(KEYINPUT48), .ZN(n465) );
  NAND2_X1 U402 ( .A1(n391), .A2(n644), .ZN(n506) );
  XNOR2_X1 U403 ( .A(n528), .B(G137), .ZN(n471) );
  XNOR2_X1 U404 ( .A(n353), .B(n493), .ZN(n467) );
  INV_X1 U405 ( .A(KEYINPUT3), .ZN(n493) );
  XNOR2_X1 U406 ( .A(n746), .B(KEYINPUT80), .ZN(n377) );
  OR2_X1 U407 ( .A1(n718), .A2(G902), .ZN(n398) );
  NOR2_X1 U408 ( .A1(n507), .A2(n358), .ZN(n435) );
  INV_X1 U409 ( .A(n507), .ZN(n436) );
  NAND2_X1 U410 ( .A1(n373), .A2(n726), .ZN(n372) );
  INV_X1 U411 ( .A(n386), .ZN(n373) );
  INV_X1 U412 ( .A(KEYINPUT81), .ZN(n464) );
  XNOR2_X1 U413 ( .A(n367), .B(KEYINPUT91), .ZN(n389) );
  XNOR2_X1 U414 ( .A(n547), .B(n462), .ZN(n704) );
  XNOR2_X1 U415 ( .A(n463), .B(KEYINPUT33), .ZN(n462) );
  INV_X1 U416 ( .A(KEYINPUT112), .ZN(n463) );
  OR2_X1 U417 ( .A1(n663), .A2(n622), .ZN(n604) );
  XNOR2_X1 U418 ( .A(n606), .B(KEYINPUT85), .ZN(n580) );
  XNOR2_X1 U419 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n631) );
  XOR2_X1 U420 ( .A(G131), .B(G140), .Z(n555) );
  XNOR2_X2 U421 ( .A(G146), .B(G125), .ZN(n502) );
  AND2_X1 U422 ( .A1(n758), .A2(n655), .ZN(n483) );
  XNOR2_X1 U423 ( .A(n502), .B(KEYINPUT10), .ZN(n556) );
  XNOR2_X1 U424 ( .A(n457), .B(n456), .ZN(n531) );
  XNOR2_X1 U425 ( .A(G110), .B(KEYINPUT96), .ZN(n456) );
  XNOR2_X1 U426 ( .A(n458), .B(G107), .ZN(n457) );
  INV_X1 U427 ( .A(G104), .ZN(n458) );
  INV_X1 U428 ( .A(n555), .ZN(n455) );
  AND2_X1 U429 ( .A1(n739), .A2(n647), .ZN(n378) );
  AND2_X1 U430 ( .A1(n673), .A2(n646), .ZN(n403) );
  AND2_X1 U431 ( .A1(n479), .A2(n359), .ZN(n476) );
  XNOR2_X1 U432 ( .A(n408), .B(n543), .ZN(n649) );
  XNOR2_X1 U433 ( .A(n387), .B(n537), .ZN(n408) );
  XNOR2_X1 U434 ( .A(G131), .B(KEYINPUT5), .ZN(n541) );
  XNOR2_X1 U435 ( .A(n537), .B(n426), .ZN(n732) );
  XNOR2_X1 U436 ( .A(n531), .B(n494), .ZN(n426) );
  XOR2_X1 U437 ( .A(G122), .B(KEYINPUT16), .Z(n494) );
  XNOR2_X1 U438 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n510) );
  XNOR2_X1 U439 ( .A(G116), .B(G107), .ZN(n562) );
  XOR2_X1 U440 ( .A(KEYINPUT107), .B(G122), .Z(n563) );
  INV_X1 U441 ( .A(n748), .ZN(n532) );
  INV_X1 U442 ( .A(n609), .ZN(n674) );
  XNOR2_X1 U443 ( .A(n628), .B(KEYINPUT115), .ZN(n703) );
  XNOR2_X1 U444 ( .A(n410), .B(n409), .ZN(n641) );
  INV_X1 U445 ( .A(KEYINPUT39), .ZN(n409) );
  NOR2_X1 U446 ( .A1(n629), .A2(n689), .ZN(n410) );
  INV_X1 U447 ( .A(KEYINPUT1), .ZN(n459) );
  INV_X1 U448 ( .A(KEYINPUT34), .ZN(n460) );
  XNOR2_X1 U449 ( .A(n578), .B(n577), .ZN(n581) );
  XNOR2_X1 U450 ( .A(n576), .B(KEYINPUT76), .ZN(n577) );
  NAND2_X1 U451 ( .A1(n575), .A2(n574), .ZN(n578) );
  NOR2_X1 U452 ( .A1(n622), .A2(n621), .ZN(n623) );
  AND2_X1 U453 ( .A1(n394), .A2(n437), .ZN(n393) );
  NAND2_X1 U454 ( .A1(n440), .A2(n351), .ZN(n396) );
  NOR2_X1 U455 ( .A1(n674), .A2(n581), .ZN(n583) );
  INV_X1 U456 ( .A(KEYINPUT6), .ZN(n407) );
  NAND2_X1 U457 ( .A1(n368), .A2(n379), .ZN(n450) );
  AND2_X1 U458 ( .A1(n386), .A2(G472), .ZN(n368) );
  AND2_X1 U459 ( .A1(n374), .A2(n371), .ZN(n370) );
  AND2_X1 U460 ( .A1(n372), .A2(n424), .ZN(n371) );
  INV_X1 U461 ( .A(KEYINPUT47), .ZN(n414) );
  XNOR2_X1 U462 ( .A(G143), .B(G113), .ZN(n548) );
  OR2_X1 U463 ( .A1(G237), .A2(G902), .ZN(n503) );
  XOR2_X1 U464 ( .A(KEYINPUT78), .B(KEYINPUT105), .Z(n539) );
  NOR2_X1 U465 ( .A1(n643), .A2(n405), .ZN(n404) );
  INV_X1 U466 ( .A(n673), .ZN(n405) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n485) );
  XOR2_X1 U468 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n486) );
  XNOR2_X1 U469 ( .A(n586), .B(n536), .ZN(n546) );
  INV_X1 U470 ( .A(KEYINPUT111), .ZN(n536) );
  NOR2_X1 U471 ( .A1(n690), .A2(n689), .ZN(n693) );
  INV_X1 U472 ( .A(n587), .ZN(n575) );
  XNOR2_X1 U473 ( .A(KEYINPUT75), .B(KEYINPUT102), .ZN(n514) );
  XNOR2_X1 U474 ( .A(G128), .B(G137), .ZN(n512) );
  XNOR2_X1 U475 ( .A(G119), .B(KEYINPUT103), .ZN(n518) );
  XNOR2_X1 U476 ( .A(n531), .B(n455), .ZN(n534) );
  NAND2_X2 U477 ( .A1(n390), .A2(n648), .ZN(n386) );
  NAND2_X1 U478 ( .A1(n378), .A2(n377), .ZN(n390) );
  XNOR2_X1 U479 ( .A(n495), .B(n355), .ZN(n427) );
  BUF_X1 U480 ( .A(n746), .Z(n413) );
  NOR2_X1 U481 ( .A1(n474), .A2(n475), .ZN(n473) );
  NOR2_X1 U482 ( .A1(n690), .A2(n441), .ZN(n439) );
  NAND2_X1 U483 ( .A1(n434), .A2(n441), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n566), .B(n420), .ZN(n728) );
  NAND2_X1 U485 ( .A1(n382), .A2(n399), .ZN(n381) );
  NOR2_X1 U486 ( .A1(n400), .A2(n731), .ZN(n399) );
  NOR2_X1 U487 ( .A1(n402), .A2(G210), .ZN(n400) );
  XNOR2_X1 U488 ( .A(KEYINPUT42), .B(KEYINPUT116), .ZN(n468) );
  XNOR2_X1 U489 ( .A(n630), .B(KEYINPUT40), .ZN(n761) );
  NOR2_X1 U490 ( .A1(n637), .A2(n434), .ZN(n607) );
  XNOR2_X1 U491 ( .A(n461), .B(n460), .ZN(n570) );
  NOR2_X1 U492 ( .A1(n581), .A2(n442), .ZN(n392) );
  NAND2_X1 U493 ( .A1(n580), .A2(n354), .ZN(n442) );
  NAND2_X1 U494 ( .A1(n583), .A2(n357), .ZN(n655) );
  XNOR2_X1 U495 ( .A(n450), .B(n363), .ZN(n449) );
  INV_X1 U496 ( .A(KEYINPUT60), .ZN(n423) );
  NAND2_X1 U497 ( .A1(n370), .A2(n369), .ZN(n376) );
  OR2_X1 U498 ( .A1(n383), .A2(n425), .ZN(n369) );
  OR2_X1 U499 ( .A1(n614), .A2(KEYINPUT19), .ZN(n350) );
  AND2_X1 U500 ( .A1(n438), .A2(n435), .ZN(n351) );
  XNOR2_X1 U501 ( .A(n467), .B(n492), .ZN(n537) );
  XOR2_X1 U502 ( .A(n505), .B(n504), .Z(n352) );
  XOR2_X1 U503 ( .A(KEYINPUT74), .B(G119), .Z(n353) );
  XNOR2_X1 U504 ( .A(KEYINPUT110), .B(n579), .ZN(n354) );
  XOR2_X1 U505 ( .A(n502), .B(KEYINPUT17), .Z(n355) );
  AND2_X1 U506 ( .A1(n453), .A2(n422), .ZN(n356) );
  AND2_X1 U507 ( .A1(n621), .A2(n677), .ZN(n357) );
  XOR2_X1 U508 ( .A(KEYINPUT0), .B(KEYINPUT93), .Z(n358) );
  OR2_X1 U509 ( .A1(n614), .A2(n480), .ZN(n359) );
  INV_X1 U510 ( .A(n615), .ZN(n480) );
  AND2_X1 U511 ( .A1(n432), .A2(n358), .ZN(n360) );
  INV_X1 U512 ( .A(KEYINPUT19), .ZN(n441) );
  AND2_X1 U513 ( .A1(n402), .A2(G210), .ZN(n361) );
  NOR2_X1 U514 ( .A1(n532), .A2(G952), .ZN(n731) );
  INV_X1 U515 ( .A(n731), .ZN(n424) );
  XNOR2_X1 U516 ( .A(KEYINPUT90), .B(KEYINPUT45), .ZN(n362) );
  XOR2_X1 U517 ( .A(KEYINPUT62), .B(n649), .Z(n363) );
  INV_X1 U518 ( .A(KEYINPUT44), .ZN(n454) );
  XOR2_X1 U519 ( .A(n730), .B(KEYINPUT122), .Z(n364) );
  XOR2_X1 U520 ( .A(KEYINPUT32), .B(KEYINPUT84), .Z(n365) );
  INV_X1 U521 ( .A(n726), .ZN(n425) );
  XNOR2_X1 U522 ( .A(n725), .B(n724), .ZN(n726) );
  INV_X1 U523 ( .A(n716), .ZN(n402) );
  XNOR2_X1 U524 ( .A(G902), .B(KEYINPUT15), .ZN(n644) );
  XOR2_X1 U525 ( .A(KEYINPUT63), .B(KEYINPUT95), .Z(n366) );
  NOR2_X1 U526 ( .A1(n381), .A2(n401), .ZN(n380) );
  NAND2_X1 U527 ( .A1(n640), .A2(n404), .ZN(n367) );
  NAND2_X1 U528 ( .A1(n383), .A2(n375), .ZN(n374) );
  AND2_X1 U529 ( .A1(n386), .A2(n425), .ZN(n375) );
  XNOR2_X1 U530 ( .A(n376), .B(n423), .ZN(G60) );
  AND2_X1 U531 ( .A1(n640), .A2(n403), .ZN(n746) );
  XNOR2_X2 U532 ( .A(n595), .B(n362), .ZN(n739) );
  NAND2_X1 U533 ( .A1(n386), .A2(n379), .ZN(n385) );
  AND2_X1 U534 ( .A1(n379), .A2(G475), .ZN(n383) );
  NAND2_X1 U535 ( .A1(n379), .A2(n709), .ZN(n712) );
  NAND2_X1 U536 ( .A1(n470), .A2(n379), .ZN(n447) );
  XNOR2_X2 U537 ( .A(n388), .B(n464), .ZN(n379) );
  XNOR2_X1 U538 ( .A(n380), .B(n717), .ZN(G51) );
  NAND2_X1 U539 ( .A1(n384), .A2(n361), .ZN(n382) );
  NAND2_X1 U540 ( .A1(n384), .A2(G469), .ZN(n721) );
  NAND2_X1 U541 ( .A1(n384), .A2(G478), .ZN(n727) );
  AND2_X1 U542 ( .A1(n385), .A2(n716), .ZN(n401) );
  AND2_X1 U543 ( .A1(n386), .A2(G217), .ZN(n470) );
  XNOR2_X1 U544 ( .A(n387), .B(n535), .ZN(n718) );
  NAND2_X1 U545 ( .A1(n389), .A2(n739), .ZN(n388) );
  XNOR2_X1 U546 ( .A(n391), .B(n481), .ZN(n716) );
  NAND2_X1 U547 ( .A1(n395), .A2(n358), .ZN(n394) );
  NAND2_X1 U548 ( .A1(n438), .A2(n436), .ZN(n395) );
  XNOR2_X1 U549 ( .A(n397), .B(n567), .ZN(n420) );
  XNOR2_X2 U550 ( .A(n398), .B(G469), .ZN(n624) );
  XNOR2_X1 U551 ( .A(n625), .B(KEYINPUT114), .ZN(n443) );
  XNOR2_X1 U552 ( .A(n661), .B(n414), .ZN(n635) );
  AND2_X1 U553 ( .A1(n635), .A2(n634), .ZN(n448) );
  NAND2_X1 U554 ( .A1(n757), .A2(n761), .ZN(n416) );
  XNOR2_X1 U555 ( .A(n406), .B(n465), .ZN(n640) );
  NAND2_X1 U556 ( .A1(n419), .A2(n466), .ZN(n406) );
  XNOR2_X2 U557 ( .A(n418), .B(n407), .ZN(n606) );
  NOR2_X1 U558 ( .A1(n690), .A2(n615), .ZN(n478) );
  NAND2_X1 U559 ( .A1(n412), .A2(n624), .ZN(n625) );
  XNOR2_X1 U560 ( .A(n623), .B(KEYINPUT28), .ZN(n412) );
  NOR2_X1 U561 ( .A1(n636), .A2(n448), .ZN(n419) );
  NAND2_X1 U562 ( .A1(n501), .A2(n500), .ZN(n430) );
  NAND2_X1 U563 ( .A1(n626), .A2(n350), .ZN(n433) );
  NAND2_X1 U564 ( .A1(n421), .A2(n482), .ZN(n595) );
  NAND2_X1 U565 ( .A1(n473), .A2(n616), .ZN(n415) );
  XNOR2_X1 U566 ( .A(n416), .B(n631), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n417), .B(n366), .ZN(G57) );
  NAND2_X1 U568 ( .A1(n449), .A2(n424), .ZN(n417) );
  NAND2_X1 U569 ( .A1(n605), .A2(n606), .ZN(n637) );
  NAND2_X1 U570 ( .A1(n356), .A2(n451), .ZN(n421) );
  NAND2_X1 U571 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U572 ( .A1(n499), .A2(KEYINPUT94), .ZN(n429) );
  NAND2_X1 U573 ( .A1(n433), .A2(n360), .ZN(n437) );
  NAND2_X1 U574 ( .A1(n350), .A2(KEYINPUT19), .ZN(n432) );
  INV_X1 U575 ( .A(n626), .ZN(n434) );
  NAND2_X1 U576 ( .A1(n440), .A2(n438), .ZN(n632) );
  NAND2_X1 U577 ( .A1(n626), .A2(n439), .ZN(n438) );
  OR2_X1 U578 ( .A1(n703), .A2(n443), .ZN(n469) );
  NOR2_X1 U579 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U580 ( .A(n521), .B(n522), .ZN(n730) );
  XNOR2_X1 U581 ( .A(n445), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U582 ( .A1(n446), .A2(n424), .ZN(n445) );
  XNOR2_X1 U583 ( .A(n447), .B(n364), .ZN(n446) );
  NAND2_X1 U584 ( .A1(n452), .A2(n483), .ZN(n451) );
  NOR2_X1 U585 ( .A1(n759), .A2(n454), .ZN(n452) );
  NAND2_X1 U586 ( .A1(n759), .A2(n454), .ZN(n453) );
  XNOR2_X2 U587 ( .A(n571), .B(KEYINPUT35), .ZN(n759) );
  NOR2_X1 U588 ( .A1(n681), .A2(n480), .ZN(n474) );
  NAND2_X1 U589 ( .A1(n477), .A2(n476), .ZN(n475) );
  NAND2_X1 U590 ( .A1(n681), .A2(n478), .ZN(n477) );
  INV_X1 U591 ( .A(n617), .ZN(n479) );
  XNOR2_X1 U592 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n481) );
  AND2_X1 U593 ( .A1(n594), .A2(n593), .ZN(n482) );
  INV_X1 U594 ( .A(n681), .ZN(n621) );
  INV_X1 U595 ( .A(n756), .ZN(n594) );
  INV_X1 U596 ( .A(n690), .ZN(n614) );
  XNOR2_X1 U597 ( .A(n529), .B(G146), .ZN(n530) );
  INV_X1 U598 ( .A(G472), .ZN(n544) );
  INV_X1 U599 ( .A(G953), .ZN(n484) );
  XNOR2_X1 U600 ( .A(KEYINPUT64), .B(n484), .ZN(n496) );
  INV_X1 U601 ( .A(n496), .ZN(n748) );
  INV_X1 U602 ( .A(G953), .ZN(n738) );
  XNOR2_X1 U603 ( .A(n486), .B(n485), .ZN(n488) );
  NAND2_X1 U604 ( .A1(n488), .A2(G952), .ZN(n487) );
  XNOR2_X1 U605 ( .A(n487), .B(KEYINPUT100), .ZN(n702) );
  NOR2_X1 U606 ( .A1(G953), .A2(n702), .ZN(n599) );
  NOR2_X1 U607 ( .A1(G898), .A2(n738), .ZN(n734) );
  AND2_X1 U608 ( .A1(G902), .A2(n488), .ZN(n596) );
  NAND2_X1 U609 ( .A1(n734), .A2(n596), .ZN(n489) );
  XNOR2_X1 U610 ( .A(KEYINPUT101), .B(n489), .ZN(n490) );
  NOR2_X1 U611 ( .A1(n599), .A2(n490), .ZN(n507) );
  NAND2_X1 U612 ( .A1(n503), .A2(G214), .ZN(n491) );
  XNOR2_X1 U613 ( .A(n491), .B(KEYINPUT99), .ZN(n690) );
  XNOR2_X1 U614 ( .A(G116), .B(G113), .ZN(n492) );
  XOR2_X1 U615 ( .A(KEYINPUT70), .B(G101), .Z(n529) );
  XNOR2_X1 U616 ( .A(n528), .B(n529), .ZN(n495) );
  XNOR2_X2 U617 ( .A(G143), .B(G128), .ZN(n527) );
  XNOR2_X1 U618 ( .A(n527), .B(KEYINPUT18), .ZN(n498) );
  NAND2_X1 U619 ( .A1(G224), .A2(n496), .ZN(n497) );
  XNOR2_X1 U620 ( .A(n498), .B(n497), .ZN(n499) );
  INV_X1 U621 ( .A(n499), .ZN(n501) );
  INV_X1 U622 ( .A(KEYINPUT94), .ZN(n500) );
  XOR2_X1 U623 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n505) );
  NAND2_X1 U624 ( .A1(G210), .A2(n503), .ZN(n504) );
  XNOR2_X2 U625 ( .A(n506), .B(n352), .ZN(n626) );
  NAND2_X1 U626 ( .A1(n644), .A2(G234), .ZN(n508) );
  XNOR2_X1 U627 ( .A(n508), .B(KEYINPUT20), .ZN(n523) );
  NAND2_X1 U628 ( .A1(G221), .A2(n523), .ZN(n509) );
  XNOR2_X1 U629 ( .A(KEYINPUT21), .B(n509), .ZN(n678) );
  NAND2_X1 U630 ( .A1(n496), .A2(G234), .ZN(n511) );
  XNOR2_X1 U631 ( .A(n511), .B(n510), .ZN(n561) );
  NAND2_X1 U632 ( .A1(n561), .A2(G221), .ZN(n522) );
  XOR2_X1 U633 ( .A(G140), .B(G110), .Z(n513) );
  XNOR2_X1 U634 ( .A(n513), .B(n512), .ZN(n517) );
  XOR2_X1 U635 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n515) );
  XNOR2_X1 U636 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U637 ( .A(n517), .B(n516), .ZN(n520) );
  XNOR2_X1 U638 ( .A(n518), .B(n556), .ZN(n519) );
  XNOR2_X1 U639 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U640 ( .A(KEYINPUT104), .B(KEYINPUT25), .Z(n525) );
  NAND2_X1 U641 ( .A1(G217), .A2(n523), .ZN(n524) );
  XNOR2_X1 U642 ( .A(n525), .B(n524), .ZN(n526) );
  INV_X1 U643 ( .A(n602), .ZN(n677) );
  NAND2_X1 U644 ( .A1(G227), .A2(n532), .ZN(n533) );
  XNOR2_X1 U645 ( .A(n534), .B(n533), .ZN(n535) );
  NOR2_X1 U646 ( .A1(G953), .A2(G237), .ZN(n550) );
  NAND2_X1 U647 ( .A1(n550), .A2(G210), .ZN(n538) );
  XNOR2_X1 U648 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U649 ( .A(n540), .B(KEYINPUT79), .Z(n542) );
  XNOR2_X1 U650 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X2 U651 ( .A(n545), .B(n544), .ZN(n681) );
  NAND2_X1 U652 ( .A1(n546), .A2(n606), .ZN(n547) );
  XOR2_X1 U653 ( .A(G122), .B(G104), .Z(n549) );
  XNOR2_X1 U654 ( .A(n549), .B(n548), .ZN(n554) );
  XOR2_X1 U655 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n552) );
  NAND2_X1 U656 ( .A1(G214), .A2(n550), .ZN(n551) );
  XNOR2_X1 U657 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U658 ( .A(n554), .B(n553), .ZN(n557) );
  XNOR2_X1 U659 ( .A(n556), .B(n555), .ZN(n744) );
  XNOR2_X1 U660 ( .A(n557), .B(n744), .ZN(n725) );
  NOR2_X1 U661 ( .A1(G902), .A2(n725), .ZN(n559) );
  XNOR2_X1 U662 ( .A(KEYINPUT106), .B(KEYINPUT13), .ZN(n558) );
  XNOR2_X1 U663 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U664 ( .A(G475), .B(n560), .Z(n591) );
  INV_X1 U665 ( .A(n591), .ZN(n572) );
  XNOR2_X1 U666 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n567) );
  NAND2_X1 U667 ( .A1(n561), .A2(G217), .ZN(n565) );
  XNOR2_X1 U668 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U669 ( .A(n565), .B(n564), .ZN(n566) );
  NOR2_X1 U670 ( .A1(G902), .A2(n728), .ZN(n568) );
  XOR2_X1 U671 ( .A(G478), .B(n568), .Z(n590) );
  NAND2_X1 U672 ( .A1(n572), .A2(n590), .ZN(n618) );
  XNOR2_X1 U673 ( .A(KEYINPUT83), .B(n618), .ZN(n569) );
  NAND2_X1 U674 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U675 ( .A1(n590), .A2(n572), .ZN(n691) );
  INV_X1 U676 ( .A(n678), .ZN(n573) );
  AND2_X1 U677 ( .A1(n691), .A2(n573), .ZN(n574) );
  XOR2_X1 U678 ( .A(KEYINPUT67), .B(KEYINPUT22), .Z(n576) );
  NOR2_X1 U679 ( .A1(n602), .A2(n609), .ZN(n579) );
  NOR2_X1 U680 ( .A1(n677), .A2(n606), .ZN(n582) );
  NAND2_X1 U681 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U682 ( .A(KEYINPUT109), .B(n584), .ZN(n756) );
  NAND2_X1 U683 ( .A1(n624), .A2(n675), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n587), .A2(n613), .ZN(n585) );
  NAND2_X1 U685 ( .A1(n585), .A2(n621), .ZN(n651) );
  NAND2_X1 U686 ( .A1(n418), .A2(n586), .ZN(n686) );
  NOR2_X1 U687 ( .A1(n686), .A2(n587), .ZN(n588) );
  XNOR2_X1 U688 ( .A(n588), .B(KEYINPUT31), .ZN(n665) );
  NAND2_X1 U689 ( .A1(n651), .A2(n665), .ZN(n592) );
  NAND2_X1 U690 ( .A1(n591), .A2(n590), .ZN(n589) );
  XOR2_X1 U691 ( .A(KEYINPUT108), .B(n589), .Z(n656) );
  NOR2_X1 U692 ( .A1(n656), .A2(n660), .ZN(n610) );
  INV_X1 U693 ( .A(n610), .ZN(n694) );
  NAND2_X1 U694 ( .A1(n592), .A2(n694), .ZN(n593) );
  INV_X1 U695 ( .A(n660), .ZN(n663) );
  NAND2_X1 U696 ( .A1(n596), .A2(n748), .ZN(n597) );
  NOR2_X1 U697 ( .A1(G900), .A2(n597), .ZN(n598) );
  NOR2_X1 U698 ( .A1(n599), .A2(n598), .ZN(n617) );
  NOR2_X1 U699 ( .A1(n678), .A2(n617), .ZN(n600) );
  XNOR2_X1 U700 ( .A(n600), .B(KEYINPUT73), .ZN(n601) );
  XOR2_X1 U701 ( .A(KEYINPUT72), .B(n603), .Z(n622) );
  NOR2_X1 U702 ( .A1(n690), .A2(n604), .ZN(n605) );
  XOR2_X1 U703 ( .A(KEYINPUT36), .B(n607), .Z(n608) );
  NOR2_X1 U704 ( .A1(n609), .A2(n608), .ZN(n668) );
  NAND2_X1 U705 ( .A1(n610), .A2(KEYINPUT47), .ZN(n611) );
  XOR2_X1 U706 ( .A(KEYINPUT88), .B(n611), .Z(n612) );
  NOR2_X1 U707 ( .A1(n668), .A2(n612), .ZN(n620) );
  INV_X1 U708 ( .A(n613), .ZN(n616) );
  XOR2_X1 U709 ( .A(KEYINPUT113), .B(KEYINPUT30), .Z(n615) );
  NOR2_X1 U710 ( .A1(n629), .A2(n618), .ZN(n619) );
  NAND2_X1 U711 ( .A1(n619), .A2(n626), .ZN(n659) );
  NAND2_X1 U712 ( .A1(n620), .A2(n659), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n693), .A2(n691), .ZN(n627) );
  XNOR2_X1 U714 ( .A(n627), .B(KEYINPUT41), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n641), .A2(n660), .ZN(n630) );
  OR2_X1 U716 ( .A1(KEYINPUT47), .A2(n694), .ZN(n634) );
  OR2_X1 U717 ( .A1(n674), .A2(n637), .ZN(n638) );
  XNOR2_X1 U718 ( .A(KEYINPUT43), .B(n638), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n639), .A2(n434), .ZN(n673) );
  NAND2_X1 U720 ( .A1(n641), .A2(n656), .ZN(n646) );
  NAND2_X1 U721 ( .A1(KEYINPUT2), .A2(n646), .ZN(n642) );
  XOR2_X1 U722 ( .A(KEYINPUT87), .B(n642), .Z(n643) );
  INV_X1 U723 ( .A(n644), .ZN(n647) );
  NAND2_X1 U724 ( .A1(KEYINPUT2), .A2(n647), .ZN(n645) );
  XOR2_X1 U725 ( .A(n645), .B(KEYINPUT69), .Z(n648) );
  INV_X1 U726 ( .A(n646), .ZN(n671) );
  NOR2_X1 U727 ( .A1(n663), .A2(n651), .ZN(n650) );
  XOR2_X1 U728 ( .A(G104), .B(n650), .Z(G6) );
  INV_X1 U729 ( .A(n656), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n666), .A2(n651), .ZN(n653) );
  XNOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U733 ( .A(G107), .B(n654), .ZN(G9) );
  XNOR2_X1 U734 ( .A(G110), .B(n655), .ZN(G12) );
  XOR2_X1 U735 ( .A(G128), .B(KEYINPUT29), .Z(n658) );
  NAND2_X1 U736 ( .A1(n661), .A2(n656), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n658), .B(n657), .ZN(G30) );
  XNOR2_X1 U738 ( .A(G143), .B(n659), .ZN(G45) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(G146), .ZN(G48) );
  NOR2_X1 U741 ( .A1(n663), .A2(n665), .ZN(n664) );
  XOR2_X1 U742 ( .A(G113), .B(n664), .Z(G15) );
  NOR2_X1 U743 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U744 ( .A(G116), .B(n667), .Z(G18) );
  XOR2_X1 U745 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n670) );
  XNOR2_X1 U746 ( .A(G125), .B(n668), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n670), .B(n669), .ZN(G27) );
  XNOR2_X1 U748 ( .A(G134), .B(KEYINPUT118), .ZN(n672) );
  XOR2_X1 U749 ( .A(n672), .B(n671), .Z(G36) );
  XNOR2_X1 U750 ( .A(G140), .B(n673), .ZN(G42) );
  NOR2_X1 U751 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U752 ( .A(KEYINPUT50), .B(n676), .Z(n684) );
  XOR2_X1 U753 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n680) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n680), .B(n679), .ZN(n682) );
  NOR2_X1 U756 ( .A1(n682), .A2(n418), .ZN(n683) );
  NAND2_X1 U757 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U758 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U759 ( .A(KEYINPUT51), .B(n687), .ZN(n688) );
  NOR2_X1 U760 ( .A1(n703), .A2(n688), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U765 ( .A1(n704), .A2(n697), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(KEYINPUT52), .ZN(n701) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U771 ( .A(n707), .B(KEYINPUT120), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n708), .A2(n738), .ZN(n714) );
  OR2_X1 U773 ( .A1(n739), .A2(KEYINPUT2), .ZN(n709) );
  NOR2_X1 U774 ( .A1(KEYINPUT2), .A2(n413), .ZN(n710) );
  XOR2_X1 U775 ( .A(KEYINPUT89), .B(n710), .Z(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U778 ( .A(n715), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U779 ( .A(KEYINPUT92), .B(KEYINPUT56), .ZN(n717) );
  XNOR2_X1 U780 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n720) );
  XNOR2_X1 U781 ( .A(n718), .B(KEYINPUT57), .ZN(n719) );
  XNOR2_X1 U782 ( .A(n720), .B(n719), .ZN(n722) );
  XNOR2_X1 U783 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U784 ( .A1(n731), .A2(n723), .ZN(G54) );
  XOR2_X1 U785 ( .A(KEYINPUT59), .B(KEYINPUT68), .Z(n724) );
  XNOR2_X1 U786 ( .A(G101), .B(n732), .ZN(n733) );
  XNOR2_X1 U787 ( .A(n733), .B(KEYINPUT124), .ZN(n735) );
  NOR2_X1 U788 ( .A1(n735), .A2(n734), .ZN(n743) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n736) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U791 ( .A1(n737), .A2(G898), .ZN(n741) );
  NAND2_X1 U792 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U794 ( .A(n743), .B(n742), .ZN(G69) );
  XOR2_X1 U795 ( .A(n745), .B(n744), .Z(n750) );
  XNOR2_X1 U796 ( .A(n750), .B(n413), .ZN(n747) );
  NOR2_X1 U797 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U798 ( .A(KEYINPUT125), .B(n749), .ZN(n754) );
  XNOR2_X1 U799 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U800 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U801 ( .A1(n752), .A2(G953), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U803 ( .A(KEYINPUT126), .B(n755), .ZN(G72) );
  XOR2_X1 U804 ( .A(G101), .B(n756), .Z(G3) );
  XNOR2_X1 U805 ( .A(G137), .B(n757), .ZN(G39) );
  XNOR2_X1 U806 ( .A(G119), .B(n758), .ZN(G21) );
  XNOR2_X1 U807 ( .A(n759), .B(G122), .ZN(n760) );
  XNOR2_X1 U808 ( .A(n760), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U809 ( .A(G131), .B(n761), .ZN(G33) );
endmodule

