

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(n712), .ZN(n696) );
  BUF_X1 U554 ( .A(n712), .Z(n720) );
  OR2_X1 U555 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U556 ( .A(KEYINPUT32), .B(KEYINPUT98), .ZN(n516) );
  OR2_X1 U557 ( .A1(n739), .A2(n738), .ZN(n517) );
  XNOR2_X1 U558 ( .A(n691), .B(n690), .ZN(n695) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n708) );
  XNOR2_X1 U560 ( .A(n719), .B(KEYINPUT31), .ZN(n734) );
  AND2_X1 U561 ( .A1(n728), .A2(n727), .ZN(n730) );
  AND2_X1 U562 ( .A1(n740), .A2(n517), .ZN(n757) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NOR2_X1 U564 ( .A1(n521), .A2(n520), .ZN(n890) );
  NOR2_X1 U565 ( .A1(n527), .A2(n526), .ZN(G164) );
  AND2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U567 ( .A1(G114), .A2(n889), .ZN(n519) );
  INV_X1 U568 ( .A(G2105), .ZN(n521) );
  XNOR2_X1 U569 ( .A(KEYINPUT64), .B(G2104), .ZN(n520) );
  AND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(n886) );
  NAND2_X1 U571 ( .A1(G102), .A2(n886), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n519), .A2(n518), .ZN(n527) );
  NAND2_X1 U573 ( .A1(G126), .A2(n890), .ZN(n522) );
  XNOR2_X1 U574 ( .A(n522), .B(KEYINPUT86), .ZN(n525) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n523), .Z(n885) );
  NAND2_X1 U576 ( .A1(n885), .A2(G138), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U578 ( .A1(G137), .A2(n885), .ZN(n528) );
  XOR2_X1 U579 ( .A(n528), .B(KEYINPUT65), .Z(n531) );
  NAND2_X1 U580 ( .A1(G101), .A2(n886), .ZN(n529) );
  XOR2_X1 U581 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U583 ( .A1(G113), .A2(n889), .ZN(n533) );
  NAND2_X1 U584 ( .A1(G125), .A2(n890), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X2 U586 ( .A1(n535), .A2(n534), .ZN(G160) );
  NOR2_X1 U587 ( .A1(G543), .A2(G651), .ZN(n640) );
  NAND2_X1 U588 ( .A1(G85), .A2(n640), .ZN(n537) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n637) );
  INV_X1 U590 ( .A(G651), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n637), .A2(n538), .ZN(n644) );
  NAND2_X1 U592 ( .A1(G72), .A2(n644), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n543) );
  NOR2_X1 U594 ( .A1(G651), .A2(n637), .ZN(n641) );
  NAND2_X1 U595 ( .A1(G47), .A2(n641), .ZN(n541) );
  NOR2_X1 U596 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n539), .Z(n648) );
  NAND2_X1 U598 ( .A1(G60), .A2(n648), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U600 ( .A1(n543), .A2(n542), .ZN(G290) );
  NAND2_X1 U601 ( .A1(G52), .A2(n641), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G64), .A2(n648), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U604 ( .A(KEYINPUT66), .B(n546), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G90), .A2(n640), .ZN(n548) );
  NAND2_X1 U606 ( .A1(G77), .A2(n644), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U609 ( .A1(n551), .A2(n550), .ZN(G171) );
  XOR2_X1 U610 ( .A(G860), .B(KEYINPUT70), .Z(n598) );
  NAND2_X1 U611 ( .A1(G56), .A2(n648), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT14), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G43), .A2(n641), .ZN(n553) );
  XOR2_X1 U614 ( .A(KEYINPUT69), .B(n553), .Z(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n640), .A2(G81), .ZN(n556) );
  XNOR2_X1 U617 ( .A(n556), .B(KEYINPUT12), .ZN(n558) );
  NAND2_X1 U618 ( .A1(G68), .A2(n644), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U620 ( .A(KEYINPUT13), .B(n559), .Z(n560) );
  NOR2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n972) );
  INV_X1 U622 ( .A(n972), .ZN(n693) );
  OR2_X1 U623 ( .A1(n598), .A2(n693), .ZN(G153) );
  INV_X1 U624 ( .A(G82), .ZN(G220) );
  INV_X1 U625 ( .A(G108), .ZN(G238) );
  NAND2_X1 U626 ( .A1(G51), .A2(n641), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G63), .A2(n648), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(KEYINPUT6), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT73), .ZN(n572) );
  XNOR2_X1 U631 ( .A(KEYINPUT5), .B(KEYINPUT72), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n640), .A2(G89), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT4), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G76), .A2(n644), .ZN(n567) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT7), .B(n573), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT74), .B(n574), .ZN(G286) );
  NAND2_X1 U641 ( .A1(G94), .A2(G452), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n833) );
  NAND2_X1 U646 ( .A1(n833), .A2(G567), .ZN(n577) );
  XOR2_X1 U647 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G92), .A2(n640), .ZN(n579) );
  NAND2_X1 U651 ( .A1(G79), .A2(n644), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G54), .A2(n641), .ZN(n581) );
  NAND2_X1 U654 ( .A1(G66), .A2(n648), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U657 ( .A(KEYINPUT15), .B(n584), .Z(n585) );
  XNOR2_X1 U658 ( .A(KEYINPUT71), .B(n585), .ZN(n961) );
  INV_X1 U659 ( .A(G868), .ZN(n658) );
  NAND2_X1 U660 ( .A1(n961), .A2(n658), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U662 ( .A1(G53), .A2(n641), .ZN(n589) );
  NAND2_X1 U663 ( .A1(G65), .A2(n648), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G91), .A2(n640), .ZN(n591) );
  NAND2_X1 U666 ( .A1(G78), .A2(n644), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n971) );
  INV_X1 U669 ( .A(n971), .ZN(G299) );
  XNOR2_X1 U670 ( .A(KEYINPUT75), .B(G868), .ZN(n594) );
  NOR2_X1 U671 ( .A1(G286), .A2(n594), .ZN(n596) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U674 ( .A(KEYINPUT76), .B(n597), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n598), .A2(G559), .ZN(n599) );
  INV_X1 U676 ( .A(n961), .ZN(n615) );
  NAND2_X1 U677 ( .A1(n599), .A2(n615), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G559), .A2(n658), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n615), .A2(n601), .ZN(n602) );
  XNOR2_X1 U681 ( .A(n602), .B(KEYINPUT77), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n693), .A2(G868), .ZN(n603) );
  NOR2_X1 U683 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G135), .A2(n885), .ZN(n606) );
  NAND2_X1 U685 ( .A1(G111), .A2(n889), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G123), .A2(n890), .ZN(n607) );
  XNOR2_X1 U688 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n886), .A2(G99), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n918) );
  XNOR2_X1 U692 ( .A(n918), .B(G2096), .ZN(n612) );
  XNOR2_X1 U693 ( .A(n612), .B(KEYINPUT78), .ZN(n614) );
  INV_X1 U694 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G559), .A2(n615), .ZN(n616) );
  XNOR2_X1 U697 ( .A(n616), .B(n693), .ZN(n656) );
  NOR2_X1 U698 ( .A1(n656), .A2(G860), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G80), .A2(n644), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G55), .A2(n641), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U702 ( .A1(G93), .A2(n640), .ZN(n619) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n619), .ZN(n620) );
  NOR2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n648), .A2(G67), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n659) );
  XOR2_X1 U707 ( .A(n659), .B(KEYINPUT80), .Z(n624) );
  XNOR2_X1 U708 ( .A(n625), .B(n624), .ZN(G145) );
  NAND2_X1 U709 ( .A1(G88), .A2(n640), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G75), .A2(n644), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U712 ( .A(KEYINPUT82), .B(n628), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G50), .A2(n641), .ZN(n630) );
  NAND2_X1 U714 ( .A1(G62), .A2(n648), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U716 ( .A1(n632), .A2(n631), .ZN(G166) );
  NAND2_X1 U717 ( .A1(G49), .A2(n641), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U720 ( .A(KEYINPUT81), .B(n635), .Z(n636) );
  NOR2_X1 U721 ( .A1(n648), .A2(n636), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n637), .A2(G87), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G86), .A2(n640), .ZN(n643) );
  NAND2_X1 U725 ( .A1(G48), .A2(n641), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n644), .A2(G73), .ZN(n645) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n645), .Z(n646) );
  NOR2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n648), .A2(G61), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(G305) );
  XNOR2_X1 U732 ( .A(G166), .B(G288), .ZN(n655) );
  XNOR2_X1 U733 ( .A(KEYINPUT19), .B(G290), .ZN(n651) );
  XNOR2_X1 U734 ( .A(n651), .B(G305), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n971), .B(n652), .ZN(n653) );
  XNOR2_X1 U736 ( .A(n653), .B(n659), .ZN(n654) );
  XNOR2_X1 U737 ( .A(n655), .B(n654), .ZN(n901) );
  XOR2_X1 U738 ( .A(n656), .B(n901), .Z(n657) );
  NAND2_X1 U739 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U748 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  NAND2_X1 U749 ( .A1(G120), .A2(G69), .ZN(n666) );
  XOR2_X1 U750 ( .A(KEYINPUT83), .B(n666), .Z(n667) );
  NOR2_X1 U751 ( .A1(G238), .A2(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(G57), .A2(n668), .ZN(n838) );
  NAND2_X1 U753 ( .A1(G567), .A2(n838), .ZN(n673) );
  NOR2_X1 U754 ( .A1(G219), .A2(G220), .ZN(n669) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U756 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U757 ( .A1(G96), .A2(n671), .ZN(n839) );
  NAND2_X1 U758 ( .A1(G2106), .A2(n839), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U760 ( .A(KEYINPUT84), .B(n674), .Z(G319) );
  INV_X1 U761 ( .A(G319), .ZN(n676) );
  NAND2_X1 U762 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n835) );
  NAND2_X1 U764 ( .A1(n835), .A2(G36), .ZN(n677) );
  XOR2_X1 U765 ( .A(KEYINPUT85), .B(n677), .Z(G176) );
  XNOR2_X1 U766 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NAND2_X1 U768 ( .A1(G40), .A2(G160), .ZN(n678) );
  XNOR2_X1 U769 ( .A(KEYINPUT89), .B(n678), .ZN(n769) );
  NAND2_X1 U770 ( .A1(n771), .A2(n769), .ZN(n712) );
  OR2_X1 U771 ( .A1(n696), .A2(G1961), .ZN(n680) );
  XNOR2_X1 U772 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NAND2_X1 U773 ( .A1(n696), .A2(n943), .ZN(n679) );
  NAND2_X1 U774 ( .A1(n680), .A2(n679), .ZN(n716) );
  AND2_X1 U775 ( .A1(n716), .A2(G171), .ZN(n681) );
  XOR2_X1 U776 ( .A(KEYINPUT94), .B(n681), .Z(n711) );
  NAND2_X1 U777 ( .A1(G1956), .A2(n720), .ZN(n682) );
  XNOR2_X1 U778 ( .A(KEYINPUT95), .B(n682), .ZN(n685) );
  NAND2_X1 U779 ( .A1(n696), .A2(G2072), .ZN(n683) );
  XNOR2_X1 U780 ( .A(KEYINPUT27), .B(n683), .ZN(n684) );
  NOR2_X1 U781 ( .A1(n685), .A2(n684), .ZN(n703) );
  NOR2_X1 U782 ( .A1(n971), .A2(n703), .ZN(n686) );
  XOR2_X1 U783 ( .A(n686), .B(KEYINPUT28), .Z(n707) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n696), .ZN(n687) );
  XNOR2_X1 U785 ( .A(n687), .B(KEYINPUT26), .ZN(n689) );
  NAND2_X1 U786 ( .A1(G1341), .A2(n720), .ZN(n688) );
  NAND2_X1 U787 ( .A1(n689), .A2(n688), .ZN(n691) );
  INV_X1 U788 ( .A(KEYINPUT96), .ZN(n690) );
  NAND2_X1 U789 ( .A1(n695), .A2(n972), .ZN(n692) );
  NAND2_X1 U790 ( .A1(n692), .A2(n961), .ZN(n702) );
  NOR2_X1 U791 ( .A1(n961), .A2(n693), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n695), .A2(n694), .ZN(n700) );
  NOR2_X1 U793 ( .A1(G2067), .A2(n720), .ZN(n698) );
  NOR2_X1 U794 ( .A1(n696), .A2(G1348), .ZN(n697) );
  NOR2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n971), .A2(n703), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U801 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n733) );
  NAND2_X1 U803 ( .A1(G8), .A2(n712), .ZN(n764) );
  NOR2_X1 U804 ( .A1(G1966), .A2(n764), .ZN(n739) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n720), .ZN(n735) );
  NOR2_X1 U806 ( .A1(n739), .A2(n735), .ZN(n713) );
  NAND2_X1 U807 ( .A1(G8), .A2(n713), .ZN(n714) );
  XNOR2_X1 U808 ( .A(KEYINPUT30), .B(n714), .ZN(n715) );
  NOR2_X1 U809 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U810 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n764), .ZN(n722) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n723), .A2(G303), .ZN(n725) );
  AND2_X1 U815 ( .A1(n734), .A2(n725), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n733), .A2(n724), .ZN(n728) );
  INV_X1 U817 ( .A(n725), .ZN(n726) );
  OR2_X1 U818 ( .A1(n726), .A2(G286), .ZN(n727) );
  INV_X1 U819 ( .A(KEYINPUT97), .ZN(n729) );
  XNOR2_X1 U820 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U821 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U822 ( .A(n732), .B(n516), .ZN(n740) );
  NAND2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n737) );
  NAND2_X1 U824 ( .A1(G8), .A2(n735), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n741) );
  XOR2_X1 U828 ( .A(n741), .B(KEYINPUT99), .Z(n742) );
  NOR2_X1 U829 ( .A1(n974), .A2(n742), .ZN(n743) );
  XOR2_X1 U830 ( .A(KEYINPUT100), .B(n743), .Z(n744) );
  NOR2_X1 U831 ( .A1(n757), .A2(n744), .ZN(n747) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NOR2_X1 U833 ( .A1(KEYINPUT101), .A2(n764), .ZN(n745) );
  NAND2_X1 U834 ( .A1(n966), .A2(n745), .ZN(n746) );
  NOR2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U836 ( .A1(KEYINPUT33), .A2(n748), .ZN(n756) );
  INV_X1 U837 ( .A(KEYINPUT101), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n974), .A2(KEYINPUT33), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n974), .A2(KEYINPUT101), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  OR2_X1 U842 ( .A1(n764), .A2(n753), .ZN(n754) );
  XOR2_X1 U843 ( .A(G1981), .B(G305), .Z(n977) );
  NAND2_X1 U844 ( .A1(n754), .A2(n977), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n768) );
  INV_X1 U846 ( .A(n757), .ZN(n760) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U848 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n761), .A2(n764), .ZN(n766) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U852 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  OR2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n783) );
  INV_X1 U856 ( .A(n769), .ZN(n770) );
  NOR2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n819) );
  NAND2_X1 U858 ( .A1(G140), .A2(n885), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G104), .A2(n886), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n774), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G116), .A2(n889), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G128), .A2(n890), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n777), .Z(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U867 ( .A(KEYINPUT36), .B(n780), .Z(n897) );
  XOR2_X1 U868 ( .A(KEYINPUT37), .B(G2067), .Z(n816) );
  AND2_X1 U869 ( .A1(n897), .A2(n816), .ZN(n923) );
  NAND2_X1 U870 ( .A1(n819), .A2(n923), .ZN(n781) );
  XNOR2_X1 U871 ( .A(KEYINPUT90), .B(n781), .ZN(n814) );
  INV_X1 U872 ( .A(n814), .ZN(n782) );
  NOR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n805) );
  NAND2_X1 U874 ( .A1(G141), .A2(n885), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G117), .A2(n889), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G105), .A2(n886), .ZN(n786) );
  XOR2_X1 U878 ( .A(KEYINPUT93), .B(n786), .Z(n787) );
  XNOR2_X1 U879 ( .A(n787), .B(KEYINPUT38), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G129), .A2(n890), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n882) );
  AND2_X1 U883 ( .A1(n882), .A2(G1996), .ZN(n801) );
  NAND2_X1 U884 ( .A1(G95), .A2(n886), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G119), .A2(n890), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U887 ( .A1(G131), .A2(n885), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G107), .A2(n889), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U891 ( .A(n798), .B(KEYINPUT91), .ZN(n866) );
  NAND2_X1 U892 ( .A1(G1991), .A2(n866), .ZN(n799) );
  XOR2_X1 U893 ( .A(KEYINPUT92), .B(n799), .Z(n800) );
  NOR2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n920) );
  XOR2_X1 U895 ( .A(G1986), .B(KEYINPUT88), .Z(n802) );
  XNOR2_X1 U896 ( .A(G290), .B(n802), .ZN(n962) );
  NAND2_X1 U897 ( .A1(n920), .A2(n962), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n803), .A2(n819), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n822) );
  NOR2_X1 U900 ( .A1(n882), .A2(G1996), .ZN(n806) );
  XNOR2_X1 U901 ( .A(n806), .B(KEYINPUT102), .ZN(n926) );
  INV_X1 U902 ( .A(n920), .ZN(n809) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n866), .ZN(n919) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n919), .A2(n807), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n926), .A2(n810), .ZN(n811) );
  XOR2_X1 U908 ( .A(n811), .B(KEYINPUT103), .Z(n812) );
  XNOR2_X1 U909 ( .A(KEYINPUT39), .B(n812), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n815), .B(KEYINPUT104), .ZN(n818) );
  NOR2_X1 U912 ( .A1(n816), .A2(n897), .ZN(n817) );
  XNOR2_X1 U913 ( .A(n817), .B(KEYINPUT105), .ZN(n931) );
  NAND2_X1 U914 ( .A1(n818), .A2(n931), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U917 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U918 ( .A(G1341), .B(G2454), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n824), .B(G2430), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n825), .B(G1348), .ZN(n831) );
  XOR2_X1 U921 ( .A(G2443), .B(G2427), .Z(n827) );
  XNOR2_X1 U922 ( .A(G2438), .B(G2446), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n827), .B(n826), .ZN(n829) );
  XOR2_X1 U924 ( .A(G2451), .B(G2435), .Z(n828) );
  XNOR2_X1 U925 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U926 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n832), .A2(G14), .ZN(n906) );
  XOR2_X1 U928 ( .A(KEYINPUT106), .B(n906), .Z(G401) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U931 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U934 ( .A(KEYINPUT107), .B(n837), .Z(G188) );
  XOR2_X1 U935 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  NOR2_X1 U939 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  XOR2_X1 U941 ( .A(G2100), .B(G2096), .Z(n841) );
  XNOR2_X1 U942 ( .A(KEYINPUT42), .B(G2678), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U944 ( .A(KEYINPUT43), .B(G2090), .Z(n843) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U947 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U950 ( .A(G1976), .B(G1961), .Z(n849) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1956), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U953 ( .A(G1981), .B(G1971), .Z(n851) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1966), .ZN(n850) );
  XNOR2_X1 U955 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U956 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U957 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n857) );
  XOR2_X1 U959 ( .A(G1991), .B(G2474), .Z(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U961 ( .A1(n890), .A2(G124), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G136), .A2(n885), .ZN(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U965 ( .A(KEYINPUT110), .B(n861), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G112), .A2(n889), .ZN(n863) );
  NAND2_X1 U967 ( .A1(G100), .A2(n886), .ZN(n862) );
  NAND2_X1 U968 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U969 ( .A1(n865), .A2(n864), .ZN(G162) );
  XNOR2_X1 U970 ( .A(n866), .B(n918), .ZN(n868) );
  XNOR2_X1 U971 ( .A(G160), .B(G164), .ZN(n867) );
  XNOR2_X1 U972 ( .A(n868), .B(n867), .ZN(n881) );
  XOR2_X1 U973 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U974 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n869) );
  XNOR2_X1 U975 ( .A(n870), .B(n869), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G118), .A2(n889), .ZN(n872) );
  NAND2_X1 U977 ( .A1(G130), .A2(n890), .ZN(n871) );
  NAND2_X1 U978 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G142), .A2(n885), .ZN(n874) );
  NAND2_X1 U980 ( .A1(G106), .A2(n886), .ZN(n873) );
  NAND2_X1 U981 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U982 ( .A(n875), .B(KEYINPUT45), .Z(n876) );
  NOR2_X1 U983 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U984 ( .A(n879), .B(n878), .Z(n880) );
  XOR2_X1 U985 ( .A(n881), .B(n880), .Z(n884) );
  XOR2_X1 U986 ( .A(n882), .B(G162), .Z(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n899) );
  NAND2_X1 U988 ( .A1(G139), .A2(n885), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G115), .A2(n889), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G127), .A2(n890), .ZN(n891) );
  NAND2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U996 ( .A(KEYINPUT113), .B(n896), .ZN(n913) );
  XOR2_X1 U997 ( .A(n913), .B(n897), .Z(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U999 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(G171), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n961), .B(n972), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n904), .B(G286), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n905), .ZN(G397) );
  NAND2_X1 U1005 ( .A1(n906), .A2(G319), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n907), .B(KEYINPUT49), .ZN(n908) );
  NOR2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(KEYINPUT114), .B(n910), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1014 ( .A(G164), .B(G2078), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(G2072), .B(KEYINPUT115), .ZN(n914) );
  XNOR2_X1 U1016 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n917), .B(KEYINPUT50), .ZN(n934) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n930) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(KEYINPUT51), .B(n928), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n935), .ZN(n937) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n938), .A2(G29), .ZN(n1020) );
  XOR2_X1 U1034 ( .A(G29), .B(KEYINPUT118), .Z(n959) );
  XOR2_X1 U1035 ( .A(G2084), .B(G34), .Z(n939) );
  XNOR2_X1 U1036 ( .A(KEYINPUT54), .B(n939), .ZN(n955) );
  XNOR2_X1 U1037 ( .A(G2090), .B(G35), .ZN(n953) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n948) );
  XOR2_X1 U1041 ( .A(G1991), .B(G25), .Z(n942) );
  NAND2_X1 U1042 ( .A1(n942), .A2(G28), .ZN(n946) );
  XOR2_X1 U1043 ( .A(G27), .B(n943), .Z(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT116), .B(n944), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G32), .B(G1996), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n951), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(KEYINPUT117), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT55), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(G11), .A2(n960), .ZN(n1018) );
  XNOR2_X1 U1056 ( .A(G16), .B(KEYINPUT56), .ZN(n986) );
  XNOR2_X1 U1057 ( .A(G1348), .B(n961), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(G171), .B(G1961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G303), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(KEYINPUT120), .B(n968), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n984) );
  XNOR2_X1 U1065 ( .A(n971), .B(G1956), .ZN(n976) );
  XOR2_X1 U1066 ( .A(G1341), .B(n972), .Z(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(G168), .B(G1966), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n979), .B(KEYINPUT57), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n980), .B(KEYINPUT119), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n1016) );
  INV_X1 U1076 ( .A(G16), .ZN(n1014) );
  XOR2_X1 U1077 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n1012) );
  XNOR2_X1 U1078 ( .A(G1961), .B(G5), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G21), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n1010) );
  XOR2_X1 U1081 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n999) );
  XOR2_X1 U1082 ( .A(KEYINPUT122), .B(G4), .Z(n990) );
  XNOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(n990), .B(n989), .ZN(n993) );
  XOR2_X1 U1085 ( .A(KEYINPUT121), .B(G1956), .Z(n991) );
  XNOR2_X1 U1086 ( .A(G20), .B(n991), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(G1341), .B(G19), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(G1981), .B(G6), .ZN(n994) );
  NOR2_X1 U1090 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1092 ( .A(n999), .B(n998), .ZN(n1008) );
  XOR2_X1 U1093 ( .A(G1986), .B(G24), .Z(n1004) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1096 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1097 ( .A(n1002), .B(KEYINPUT124), .ZN(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1099 ( .A(n1005), .B(KEYINPUT125), .Z(n1006) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1021), .B(KEYINPUT127), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1022), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

