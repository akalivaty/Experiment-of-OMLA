//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT94), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n203), .A2(KEYINPUT94), .ZN(new_n208));
  OAI21_X1  g007(.A(G8gat), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n206), .A2(KEYINPUT95), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(KEYINPUT95), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n203), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT15), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n222), .A2(KEYINPUT15), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n224), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n228), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT17), .B1(new_n228), .B2(KEYINPUT93), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n215), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n228), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n214), .B(new_n228), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n232), .B(KEYINPUT13), .Z(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n232), .A4(new_n233), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G141gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT92), .B(G197gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT11), .B(G169gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT12), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT96), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n234), .B2(new_n235), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n240), .A2(new_n239), .A3(new_n247), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n250), .A3(new_n235), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(KEYINPUT97), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT97), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n234), .A2(new_n250), .A3(new_n235), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(new_n251), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n259), .B2(new_n253), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n249), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265));
  INV_X1    g064(.A(G113gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G120gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT69), .B(G120gat), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n265), .B(new_n267), .C1(new_n268), .C2(new_n266), .ZN(new_n269));
  INV_X1    g068(.A(G134gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G127gat), .ZN(new_n271));
  INV_X1    g070(.A(G127gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G134gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n277), .A2(new_n278), .A3(new_n266), .ZN(new_n279));
  INV_X1    g078(.A(new_n267), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT70), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n282));
  XNOR2_X1  g081(.A(G113gat), .B(G120gat), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n283), .A2(KEYINPUT1), .B1(KEYINPUT67), .B2(new_n271), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n271), .A2(new_n273), .A3(KEYINPUT67), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n272), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n291), .B2(new_n274), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(KEYINPUT68), .A3(new_n285), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n276), .A2(new_n281), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G155gat), .B(G162gat), .ZN(new_n295));
  XOR2_X1   g094(.A(G141gat), .B(G148gat), .Z(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G141gat), .ZN(new_n300));
  AND2_X1   g099(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n300), .B1(new_n303), .B2(G141gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n295), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT80), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n299), .ZN(new_n310));
  NAND2_X1  g109(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(G141gat), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n300), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G155gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G162gat), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n306), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT80), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n298), .B1(new_n308), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n294), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n281), .A2(new_n269), .A3(new_n275), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n284), .A2(new_n286), .A3(new_n282), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT68), .B1(new_n292), .B2(new_n285), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n322), .A2(new_n324), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n264), .B(new_n323), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n333));
  INV_X1    g132(.A(new_n298), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n314), .A2(new_n320), .A3(new_n319), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n320), .B1(new_n314), .B2(new_n319), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n333), .B1(new_n329), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n287), .A2(new_n293), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n322), .A2(KEYINPUT81), .A3(new_n340), .A4(new_n326), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n337), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n338), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n264), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT83), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n352));
  AOI211_X1 g151(.A(new_n352), .B(new_n349), .C1(new_n346), .C2(new_n347), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n344), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n264), .B(new_n349), .C1(new_n330), .C2(new_n331), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n322), .A2(new_n339), .A3(new_n340), .A4(new_n326), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT84), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n294), .A2(new_n359), .A3(new_n339), .A4(new_n322), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n341), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n361), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n356), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n354), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT0), .ZN(new_n369));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n371), .B1(new_n354), .B2(new_n366), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(new_n371), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n348), .A2(new_n350), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n352), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n348), .A2(KEYINPUT83), .A3(new_n350), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n343), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n374), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT86), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n376), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n354), .A2(new_n366), .A3(new_n371), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(KEYINPUT86), .A3(new_n374), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n375), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT28), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT27), .B(G183gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n392), .B2(G190gat), .ZN(new_n393));
  INV_X1    g192(.A(G190gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(KEYINPUT28), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n398), .A2(KEYINPUT26), .ZN(new_n399));
  NAND2_X1  g198(.A1(G169gat), .A2(G176gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n398), .B2(KEYINPUT26), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n399), .A2(new_n402), .B1(G183gat), .B2(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G183gat), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT24), .B1(new_n406), .B2(new_n394), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT24), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(G183gat), .A3(G190gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n394), .A3(KEYINPUT64), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT64), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(G183gat), .B2(G190gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n397), .A2(KEYINPUT23), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n397), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n397), .A2(KEYINPUT23), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n401), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n415), .A2(new_n418), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT25), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n400), .A2(KEYINPUT66), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n400), .A2(KEYINPUT66), .ZN(new_n426));
  NOR4_X1   g225(.A1(new_n425), .A2(new_n420), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n410), .B1(G183gat), .B2(G190gat), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n422), .A2(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT74), .B1(new_n405), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n428), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT23), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n398), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n418), .A2(new_n435), .A3(new_n400), .A4(new_n419), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n407), .A2(new_n409), .B1(new_n411), .B2(new_n413), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n423), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n404), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n430), .A2(new_n432), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G197gat), .B(G204gat), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT22), .ZN(new_n444));
  INV_X1    g243(.A(G211gat), .ZN(new_n445));
  INV_X1    g244(.A(G218gat), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(G211gat), .B(G218gat), .Z(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT73), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n449), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT72), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n453), .A2(new_n454), .B1(new_n447), .B2(new_n443), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n454), .B2(new_n453), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n404), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n432), .A2(KEYINPUT29), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n430), .A2(new_n441), .ZN(new_n463));
  INV_X1    g262(.A(new_n459), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n463), .A2(new_n460), .B1(new_n432), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT75), .B(new_n462), .C1(new_n465), .C2(new_n458), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n442), .A2(new_n467), .A3(new_n458), .A4(new_n461), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n388), .B(new_n389), .C1(new_n469), .C2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n466), .B2(new_n468), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT76), .B1(new_n475), .B2(KEYINPUT30), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n462), .A2(KEYINPUT75), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n463), .A2(new_n460), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n464), .A2(new_n432), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n458), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n468), .B(new_n473), .C1(new_n477), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(KEYINPUT30), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n474), .A2(new_n476), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n263), .B1(new_n387), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n483), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n385), .A2(KEYINPUT86), .A3(new_n374), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT86), .B1(new_n385), .B2(new_n374), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n486), .A2(new_n487), .A3(new_n376), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT87), .B(new_n485), .C1(new_n488), .C2(new_n375), .ZN(new_n489));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT3), .B1(new_n457), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT88), .B1(new_n494), .B2(new_n322), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n325), .A2(new_n493), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n458), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n494), .A2(KEYINPUT88), .A3(new_n322), .ZN(new_n499));
  OAI211_X1 g298(.A(G228gat), .B(G233gat), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n448), .A2(new_n449), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n452), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n324), .B1(new_n502), .B2(KEYINPUT29), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n503), .A2(new_n337), .B1(G228gat), .B2(G233gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n497), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT31), .B(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n500), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n500), .B2(new_n505), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n492), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n510), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(new_n491), .A3(new_n508), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G43gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(G71gat), .B(G99gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n459), .B(new_n329), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(G227gat), .A3(G233gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT33), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(KEYINPUT32), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n519), .B(KEYINPUT32), .C1(new_n520), .C2(new_n517), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT34), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n518), .ZN(new_n530));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n530), .A2(new_n531), .B1(new_n526), .B2(new_n527), .ZN(new_n532));
  INV_X1    g331(.A(new_n528), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n523), .A2(new_n533), .A3(new_n524), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n529), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n532), .ZN(new_n536));
  INV_X1    g335(.A(new_n534), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n533), .B1(new_n523), .B2(new_n524), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n514), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n484), .A2(new_n489), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT89), .B1(new_n367), .B2(new_n372), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n544), .B(new_n371), .C1(new_n354), .C2(new_n366), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n382), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n375), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n542), .B1(new_n548), .B2(new_n483), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n373), .A2(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n376), .A2(KEYINPUT89), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n375), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT90), .A3(new_n485), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n535), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n558), .A2(KEYINPUT35), .A3(new_n514), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT35), .A2(new_n541), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n514), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n484), .B2(new_n489), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT38), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n473), .A2(KEYINPUT37), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n481), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n466), .A2(KEYINPUT37), .A3(new_n468), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n465), .A2(new_n457), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n442), .A2(new_n457), .A3(new_n461), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT37), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n563), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n481), .B2(new_n564), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n567), .A2(new_n475), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n552), .A3(new_n553), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT39), .B1(new_n346), .B2(new_n347), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n330), .A2(new_n331), .ZN(new_n577));
  INV_X1    g376(.A(new_n365), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n576), .B1(new_n580), .B2(new_n264), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n364), .A2(new_n365), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n582), .B(new_n347), .C1(new_n583), .C2(new_n577), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n371), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT40), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n581), .A2(KEYINPUT40), .A3(new_n371), .A4(new_n584), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n483), .A2(new_n587), .A3(new_n546), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n589), .A3(new_n561), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n539), .A2(new_n535), .A3(KEYINPUT36), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT36), .B1(new_n539), .B2(new_n535), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n562), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT91), .B1(new_n560), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n556), .A2(new_n559), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT91), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n484), .A2(new_n489), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n514), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n590), .A2(new_n593), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n262), .B1(new_n596), .B2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G190gat), .B(G218gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT102), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT103), .ZN(new_n609));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT41), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT98), .Z(new_n613));
  XOR2_X1   g412(.A(new_n609), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n608), .A2(KEYINPUT103), .ZN(new_n616));
  NAND2_X1  g415(.A1(G85gat), .A2(G92gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT99), .A3(KEYINPUT7), .ZN(new_n618));
  NAND2_X1  g417(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(G85gat), .A3(G92gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G92gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT100), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(G92gat), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(G99gat), .ZN(new_n628));
  INV_X1    g427(.A(G106gat), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT8), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n621), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G99gat), .B(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n621), .A2(new_n632), .A3(new_n627), .A4(new_n630), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(KEYINPUT101), .A3(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n230), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n228), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n228), .A2(new_n639), .ZN(new_n643));
  NAND3_X1  g442(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n616), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n615), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n648), .A3(new_n614), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G57gat), .B(G64gat), .Z(new_n655));
  OR2_X1    g454(.A1(G71gat), .A2(G78gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(G71gat), .A2(G78gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT9), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G57gat), .B(G64gat), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n657), .B(new_n656), .C1(new_n662), .C2(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT21), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G231gat), .A2(G233gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G127gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n215), .B1(new_n665), .B2(new_n664), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(new_n317), .ZN(new_n673));
  XOR2_X1   g472(.A(G183gat), .B(G211gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n671), .B(new_n675), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n654), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n661), .A2(new_n663), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(KEYINPUT10), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n639), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n678), .A2(new_n634), .A3(new_n636), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT104), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n637), .A2(new_n664), .A3(new_n638), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n678), .A2(new_n686), .A3(new_n634), .A4(new_n636), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT105), .B(KEYINPUT10), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n639), .A2(KEYINPUT106), .A3(new_n679), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n682), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(G230gat), .A2(G233gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT107), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n695));
  INV_X1    g494(.A(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(G120gat), .B(G148gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT108), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n691), .A2(new_n702), .A3(new_n692), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n694), .A2(new_n697), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n701), .ZN(new_n705));
  INV_X1    g504(.A(new_n693), .ZN(new_n706));
  INV_X1    g505(.A(new_n697), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n677), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n606), .A2(new_n387), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g511(.A1(new_n596), .A2(new_n605), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n713), .A2(new_n261), .A3(new_n483), .A4(new_n710), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT16), .B(G8gat), .Z(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n714), .A2(KEYINPUT42), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT42), .B1(new_n714), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n714), .A2(KEYINPUT109), .A3(G8gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n714), .A2(G8gat), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(G1325gat));
  INV_X1    g523(.A(new_n593), .ZN(new_n725));
  AND4_X1   g524(.A1(G15gat), .A2(new_n606), .A3(new_n725), .A4(new_n710), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n606), .A2(new_n557), .A3(new_n710), .ZN(new_n727));
  INV_X1    g526(.A(G15gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(KEYINPUT110), .A3(new_n728), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(G1326gat));
  NAND3_X1  g532(.A1(new_n606), .A2(new_n514), .A3(new_n710), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT43), .B(G22gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1327gat));
  NOR2_X1   g535(.A1(new_n676), .A2(new_n709), .ZN(new_n737));
  INV_X1    g536(.A(new_n654), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT111), .ZN(new_n740));
  INV_X1    g539(.A(new_n387), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(G29gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n606), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n738), .A2(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n596), .B2(new_n605), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n599), .A2(new_n604), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT44), .B1(new_n749), .B2(new_n738), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n261), .A2(new_n737), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(new_n387), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n745), .B(new_n746), .C1(new_n753), .C2(new_n220), .ZN(G1328gat));
  NOR2_X1   g553(.A1(new_n485), .A2(G36gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n606), .A2(new_n740), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n752), .A2(new_n483), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n216), .ZN(G1329gat));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  INV_X1    g560(.A(G43gat), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n752), .B2(new_n725), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n558), .A2(G43gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n606), .A2(new_n740), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n761), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NOR4_X1   g566(.A1(new_n748), .A2(new_n750), .A3(new_n593), .A4(new_n751), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n765), .B(KEYINPUT47), .C1(new_n768), .C2(new_n762), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1330gat));
  NOR2_X1   g569(.A1(new_n748), .A2(new_n750), .ZN(new_n771));
  INV_X1    g570(.A(new_n751), .ZN(new_n772));
  INV_X1    g571(.A(G50gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n561), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n606), .A2(new_n514), .A3(new_n740), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT48), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n775), .A2(new_n780), .A3(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1331gat));
  INV_X1    g581(.A(new_n709), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n261), .A2(new_n677), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n749), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n387), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n483), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT49), .B(G64gat), .Z(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n788), .B2(new_n790), .ZN(G1333gat));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n725), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n558), .A2(G71gat), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n792), .A2(G71gat), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n785), .A2(new_n514), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g596(.A(new_n654), .B1(new_n599), .B2(new_n604), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n261), .A2(new_n676), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(KEYINPUT51), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT112), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n749), .A2(new_n738), .A3(new_n799), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n798), .A2(new_n805), .A3(KEYINPUT51), .A4(new_n799), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n801), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n626), .A3(new_n387), .A4(new_n709), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n799), .A2(new_n709), .ZN(new_n809));
  NOR4_X1   g608(.A1(new_n748), .A2(new_n750), .A3(new_n741), .A4(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n626), .B2(new_n810), .ZN(G1336gat));
  NOR3_X1   g610(.A1(new_n485), .A2(G92gat), .A3(new_n783), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  NOR4_X1   g613(.A1(new_n748), .A2(new_n750), .A3(new_n485), .A4(new_n809), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n623), .A2(new_n625), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n812), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n804), .B2(new_n800), .ZN(new_n820));
  INV_X1    g619(.A(new_n748), .ZN(new_n821));
  INV_X1    g620(.A(new_n750), .ZN(new_n822));
  INV_X1    g621(.A(new_n809), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n821), .A2(new_n483), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n820), .B1(new_n824), .B2(new_n816), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n813), .A2(new_n818), .B1(new_n825), .B2(new_n814), .ZN(G1337gat));
  NAND3_X1  g625(.A1(new_n771), .A2(new_n725), .A3(new_n823), .ZN(new_n827));
  XOR2_X1   g626(.A(KEYINPUT113), .B(G99gat), .Z(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n558), .A2(new_n783), .A3(new_n828), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n807), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1338gat));
  NOR3_X1   g631(.A1(new_n561), .A2(G106gat), .A3(new_n783), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n807), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g633(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n835));
  NOR4_X1   g634(.A1(new_n748), .A2(new_n750), .A3(new_n561), .A4(new_n809), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n629), .ZN(new_n837));
  INV_X1    g636(.A(new_n833), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n804), .B2(new_n800), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n514), .A3(new_n822), .A4(new_n823), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(G106gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n834), .A2(new_n837), .B1(new_n841), .B2(new_n842), .ZN(G1339gat));
  NOR3_X1   g642(.A1(new_n261), .A2(new_n677), .A3(new_n709), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n682), .A2(new_n689), .A3(new_n696), .A4(new_n690), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n694), .A2(new_n848), .A3(new_n703), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT115), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n694), .A2(new_n848), .A3(new_n851), .A4(new_n703), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n701), .B1(new_n706), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n850), .A2(KEYINPUT55), .A3(new_n852), .A4(new_n854), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n704), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n857), .A2(KEYINPUT116), .A3(new_n704), .A4(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n255), .A2(KEYINPUT97), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n259), .A2(new_n257), .A3(new_n253), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n231), .A2(new_n233), .ZN(new_n867));
  OAI22_X1  g666(.A1(new_n867), .A2(new_n232), .B1(new_n237), .B2(new_n238), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n246), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n738), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n846), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n738), .A2(new_n866), .A3(new_n869), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n861), .A3(KEYINPUT117), .A4(new_n862), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n866), .A2(new_n709), .A3(new_n869), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n863), .B2(new_n262), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n871), .A2(new_n873), .B1(new_n875), .B2(new_n654), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n845), .B1(new_n876), .B2(new_n676), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n540), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n741), .A2(new_n483), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n262), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(new_n266), .ZN(G1340gat));
  OAI21_X1  g681(.A(new_n289), .B1(new_n880), .B2(new_n783), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n878), .A2(new_n268), .A3(new_n709), .A4(new_n879), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(G1341gat));
  INV_X1    g684(.A(new_n676), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(new_n272), .ZN(G1342gat));
  NOR3_X1   g687(.A1(new_n741), .A2(new_n483), .A3(new_n654), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n878), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT56), .B1(new_n891), .B2(new_n270), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n890), .A2(new_n893), .A3(G134gat), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n892), .A2(new_n894), .B1(new_n270), .B2(new_n891), .ZN(G1343gat));
  NOR2_X1   g694(.A1(new_n725), .A2(new_n741), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n485), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT118), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n877), .B2(new_n514), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n514), .A2(KEYINPUT57), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n871), .A2(new_n873), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n261), .A2(new_n704), .A3(new_n858), .A4(new_n857), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n738), .B1(new_n903), .B2(new_n874), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n886), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n905), .B2(new_n845), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n261), .B(new_n898), .C1(new_n899), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G141gat), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n877), .A2(new_n514), .A3(new_n896), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n483), .B1(new_n910), .B2(KEYINPUT119), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n262), .A2(G141gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n877), .A2(new_n913), .A3(new_n514), .A4(new_n896), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n908), .A2(new_n909), .A3(new_n915), .ZN(new_n916));
  NOR4_X1   g715(.A1(new_n910), .A2(G141gat), .A3(new_n262), .A4(new_n483), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n907), .B2(G141gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n918), .B2(new_n909), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n910), .A2(KEYINPUT119), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n920), .A2(new_n485), .A3(new_n709), .A4(new_n914), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT59), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n303), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n898), .B1(new_n899), .B2(new_n906), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n783), .A2(KEYINPUT59), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n870), .A2(new_n859), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n886), .B1(new_n904), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n844), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n561), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n930), .A3(KEYINPUT121), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT57), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n871), .A2(new_n873), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n875), .A2(new_n654), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n844), .B1(new_n938), .B2(new_n886), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n901), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n709), .B(new_n898), .C1(new_n935), .C2(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n925), .A2(new_n926), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n943), .ZN(G1345gat));
  XNOR2_X1  g743(.A(KEYINPUT79), .B(G155gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n924), .B2(new_n886), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n886), .A2(new_n945), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n911), .A2(new_n914), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1346gat));
  OAI21_X1  g748(.A(G162gat), .B1(new_n924), .B2(new_n654), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n654), .A2(G162gat), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n920), .A2(new_n485), .A3(new_n914), .A4(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(G1347gat));
  NOR2_X1   g755(.A1(new_n387), .A2(new_n485), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n877), .A2(new_n540), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n877), .A2(KEYINPUT123), .A3(new_n540), .A4(new_n957), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(G169gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n962), .A2(new_n963), .A3(new_n261), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n878), .A2(new_n261), .A3(new_n957), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(G169gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n965), .B2(G169gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1348gat));
  INV_X1    g768(.A(G176gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n962), .A2(new_n970), .A3(new_n709), .ZN(new_n971));
  OAI21_X1  g770(.A(G176gat), .B1(new_n958), .B2(new_n783), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  NAND4_X1  g772(.A1(new_n878), .A2(new_n392), .A3(new_n676), .A4(new_n957), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n406), .B1(new_n958), .B2(new_n886), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT60), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(G1350gat));
  OAI21_X1  g777(.A(G190gat), .B1(new_n958), .B2(new_n654), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT61), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n960), .A2(new_n394), .A3(new_n738), .A4(new_n961), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(G1351gat));
  NAND3_X1  g784(.A1(new_n593), .A2(new_n514), .A3(new_n957), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n939), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(G197gat), .B1(new_n987), .B2(new_n261), .ZN(new_n988));
  INV_X1    g787(.A(new_n957), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n725), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n990), .B1(new_n935), .B2(new_n940), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n261), .A2(G197gat), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(G1352gat));
  AOI21_X1  g793(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n987), .A2(new_n709), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g795(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n996), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g797(.A(G204gat), .B1(new_n991), .B2(new_n783), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1353gat));
  NAND3_X1  g799(.A1(new_n987), .A2(new_n445), .A3(new_n676), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n676), .B(new_n990), .C1(new_n935), .C2(new_n940), .ZN(new_n1002));
  AND3_X1   g801(.A1(new_n1002), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n1002), .B2(G211gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1354gat));
  AOI21_X1  g804(.A(G218gat), .B1(new_n987), .B2(new_n738), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n738), .A2(G218gat), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT127), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1006), .B1(new_n992), .B2(new_n1008), .ZN(G1355gat));
endmodule


