//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1189,
    new_n1190, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1243, new_n1244, new_n1245;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G50), .ZN(new_n203));
  INV_X1    g0003(.A(G226), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  INV_X1    g0005(.A(G244), .ZN(new_n206));
  OAI22_X1  g0006(.A1(new_n203), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n207), .B(new_n213), .C1(G116), .C2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT65), .Z(new_n221));
  NOR2_X1   g0021(.A1(G58), .A2(G68), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n223), .A2(G50), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n218), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NAND4_X1  g0034(.A1(new_n221), .A2(new_n230), .A3(new_n231), .A4(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G107), .ZN(new_n250));
  INV_X1    g0050(.A(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n248), .B(new_n252), .Z(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n227), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT69), .A2(G58), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n256), .B(KEYINPUT8), .Z(new_n257));
  NAND2_X1  g0057(.A1(new_n228), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n228), .B1(new_n222), .B2(new_n203), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT70), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n255), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n255), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n265), .B(new_n271), .C1(G50), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT67), .ZN(new_n278));
  AND2_X1   g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n227), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n281), .A2(KEYINPUT67), .A3(G1), .A4(G13), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G41), .A2(G45), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G1), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(G274), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT68), .B1(new_n284), .B2(G1), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT68), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n288), .B(new_n267), .C1(G41), .C2(G45), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n280), .A2(new_n282), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G223), .ZN(new_n297));
  OR2_X1    g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  AOI21_X1  g0099(.A(G1698), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n300), .A2(G222), .B1(new_n294), .B2(G77), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n279), .A2(new_n227), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n286), .B1(new_n204), .B2(new_n291), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G200), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n305), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n277), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT18), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  INV_X1    g0113(.A(G274), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n280), .B2(new_n282), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n290), .A2(G232), .B1(new_n315), .B2(new_n285), .ZN(new_n316));
  OAI211_X1 g0116(.A(G226), .B(G1698), .C1(new_n292), .C2(new_n293), .ZN(new_n317));
  OAI211_X1 g0117(.A(G223), .B(new_n295), .C1(new_n292), .C2(new_n293), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G87), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n303), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n313), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n287), .A2(new_n289), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n283), .A2(new_n323), .A3(G232), .ZN(new_n324));
  AND4_X1   g0124(.A1(G179), .A2(new_n321), .A3(new_n286), .A4(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT16), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT7), .B1(new_n294), .B2(new_n228), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n298), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n299), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n298), .A2(new_n228), .A3(new_n299), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n209), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n215), .A2(new_n209), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n338), .B2(new_n222), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n260), .A2(G159), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n327), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n333), .A2(new_n334), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n330), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n341), .B1(new_n344), .B2(G68), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n266), .B1(new_n345), .B2(KEYINPUT16), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n257), .A2(new_n269), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n273), .B2(new_n257), .ZN(new_n349));
  AOI211_X1 g0149(.A(new_n312), .B(new_n326), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT76), .B1(new_n343), .B2(new_n330), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n351), .B2(new_n335), .ZN(new_n352));
  INV_X1    g0152(.A(new_n341), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT16), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n344), .A2(G68), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT16), .A3(new_n353), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n255), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n349), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n322), .A2(new_n325), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT18), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n321), .A2(new_n286), .A3(new_n324), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT77), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n362), .A2(new_n363), .A3(G190), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT77), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n316), .A2(new_n307), .A3(new_n321), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g0169(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n370));
  OR3_X1    g0170(.A1(new_n369), .A2(new_n358), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n358), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n361), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n305), .A2(new_n313), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n275), .B1(new_n305), .B2(G179), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT8), .B(G58), .Z(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n260), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  OAI221_X1 g0183(.A(new_n382), .B1(new_n228), .B2(new_n205), .C1(new_n258), .C2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n255), .B1(new_n205), .B2(new_n273), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n205), .B2(new_n269), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n298), .A2(new_n299), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(G232), .A3(new_n295), .ZN(new_n388));
  INV_X1    g0188(.A(G107), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(G1698), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n388), .B1(new_n389), .B2(new_n387), .C1(new_n390), .C2(new_n210), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n303), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(new_n286), .C1(new_n206), .C2(new_n291), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n386), .B1(new_n393), .B2(G179), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(new_n313), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n311), .A2(new_n376), .A3(new_n380), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n290), .A2(G238), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n300), .A2(G226), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G97), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n387), .A2(G232), .A3(G1698), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n303), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT72), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n315), .A2(new_n405), .A3(new_n285), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n405), .B1(new_n315), .B2(new_n285), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n399), .B(new_n404), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT13), .ZN(new_n410));
  INV_X1    g0210(.A(new_n408), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n406), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n399), .A4(new_n404), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G200), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n410), .A2(new_n414), .A3(G190), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n270), .A2(G68), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT73), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n273), .A2(new_n209), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT12), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n261), .A2(new_n203), .B1(new_n258), .B2(new_n205), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n228), .A2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n255), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT11), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n419), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n416), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT74), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n415), .B2(G200), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT74), .A3(new_n417), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n410), .A2(new_n414), .A3(G179), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n313), .B1(new_n410), .B2(new_n414), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT75), .B(KEYINPUT14), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT75), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT14), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n415), .A2(G169), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n426), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n386), .B1(G200), .B2(new_n393), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n307), .B2(new_n393), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n433), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n398), .A2(new_n444), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n255), .B(new_n273), .C1(new_n267), .C2(G33), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(new_n389), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT23), .B1(new_n228), .B2(G107), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT23), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n389), .A3(G20), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n228), .A2(G33), .A3(G116), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT84), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT84), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n449), .A2(new_n451), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n387), .A2(new_n228), .A3(G87), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT22), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n387), .A2(KEYINPUT22), .A3(new_n228), .A4(G87), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT24), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n457), .A2(new_n464), .A3(new_n460), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n448), .B1(new_n466), .B2(new_n255), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n273), .A2(new_n389), .ZN(new_n468));
  XOR2_X1   g0268(.A(new_n468), .B(KEYINPUT25), .Z(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n300), .A2(G250), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G294), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n212), .C2(new_n390), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n303), .ZN(new_n474));
  INV_X1    g0274(.A(G41), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n267), .B(G45), .C1(new_n475), .C2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT5), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(G41), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G264), .A3(new_n283), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT79), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n476), .A2(new_n481), .B1(KEYINPUT5), .B2(new_n475), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n315), .B(new_n482), .C1(new_n481), .C2(new_n476), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n474), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n365), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n484), .A2(new_n307), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n470), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G179), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n484), .A2(KEYINPUT85), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n484), .A2(G169), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(KEYINPUT85), .C1(new_n489), .C2(new_n484), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n470), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n490), .B1(new_n467), .B2(new_n469), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT86), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n493), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n488), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(G107), .B1(new_n351), .B2(new_n335), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n389), .A2(KEYINPUT6), .A3(G97), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n211), .A2(new_n389), .ZN(new_n502));
  NOR2_X1   g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n501), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n260), .A2(G77), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n500), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n255), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n273), .A2(new_n211), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n446), .A2(G97), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT4), .ZN(new_n513));
  INV_X1    g0313(.A(new_n300), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n206), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n296), .A2(G250), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n300), .A2(KEYINPUT4), .A3(G244), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n515), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n303), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n479), .A2(G257), .A3(new_n283), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n483), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n313), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n520), .A2(new_n489), .A3(new_n483), .A4(new_n521), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n512), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(G200), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n508), .A2(new_n255), .B1(new_n211), .B2(new_n273), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n520), .A2(G190), .A3(new_n483), .A4(new_n521), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n511), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n251), .A2(G20), .ZN(new_n532));
  AOI21_X1  g0332(.A(G20), .B1(G33), .B2(G283), .ZN(new_n533));
  INV_X1    g0333(.A(G33), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G97), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT81), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT81), .B1(new_n533), .B2(new_n535), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n255), .B(new_n532), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT20), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT82), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n538), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n266), .B1(new_n542), .B2(new_n536), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT20), .A4(new_n532), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n539), .A2(new_n540), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n274), .A2(G116), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n446), .A2(G116), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n387), .A2(G264), .A3(G1698), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n294), .A2(G303), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(new_n553), .C1(new_n514), .C2(new_n212), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n303), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n479), .A2(G270), .A3(new_n283), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n483), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n557), .A2(G169), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT83), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n557), .A2(KEYINPUT21), .A3(G169), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n557), .A2(new_n489), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n551), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(KEYINPUT83), .A3(new_n560), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n557), .A2(G200), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n307), .B2(new_n557), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n569), .A2(new_n551), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n563), .A2(new_n566), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n300), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n387), .A2(G244), .A3(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n304), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n267), .A2(G45), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n283), .A2(G250), .A3(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n575), .A2(KEYINPUT67), .A3(new_n314), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  OAI21_X1  g0381(.A(G200), .B1(new_n574), .B2(new_n579), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n583), .A2(new_n228), .A3(G33), .A4(G97), .ZN(new_n584));
  INV_X1    g0384(.A(G87), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n503), .A2(new_n585), .B1(new_n401), .B2(new_n228), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n586), .B2(new_n583), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n228), .B(G68), .C1(new_n292), .C2(new_n293), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n387), .A2(KEYINPUT80), .A3(new_n228), .A4(G68), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n255), .B1(new_n273), .B2(new_n383), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n446), .A2(G87), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n581), .A2(new_n582), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n383), .B2(new_n447), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n580), .A2(new_n489), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n387), .A2(G238), .A3(new_n295), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G116), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n573), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n303), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n280), .A2(new_n282), .B1(new_n267), .B2(G45), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n577), .B1(new_n602), .B2(G250), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n313), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n596), .A2(new_n597), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n595), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n571), .A2(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n445), .A2(new_n499), .A3(new_n531), .A4(new_n608), .ZN(G372));
  INV_X1    g0409(.A(KEYINPUT26), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n592), .A2(new_n255), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n273), .A2(new_n383), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n594), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n365), .B1(new_n601), .B2(new_n603), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n582), .A2(KEYINPUT87), .A3(new_n593), .A4(new_n594), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n581), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n606), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n610), .B1(new_n619), .B2(new_n525), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT88), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n525), .A2(new_n607), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT88), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n610), .C1(new_n619), .C2(new_n525), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n563), .A2(new_n494), .A3(new_n566), .A4(new_n567), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n530), .A2(new_n619), .ZN(new_n628));
  INV_X1    g0428(.A(new_n488), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n626), .A2(new_n606), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n445), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n397), .B1(new_n430), .B2(new_n432), .ZN(new_n633));
  INV_X1    g0433(.A(new_n441), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n374), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n361), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n379), .B1(new_n636), .B2(new_n311), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n632), .A2(new_n637), .ZN(G369));
  NAND3_X1  g0438(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n272), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n267), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n551), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n639), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n571), .B2(new_n648), .ZN(new_n650));
  MUX2_X1   g0450(.A(new_n649), .B(new_n650), .S(KEYINPUT89), .Z(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  INV_X1    g0452(.A(new_n646), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n494), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT90), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n470), .A2(new_n646), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n499), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n639), .A2(new_n653), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n655), .B2(new_n657), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n494), .A2(new_n646), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n232), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n503), .A2(new_n585), .A3(new_n251), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n666), .A2(new_n667), .A3(new_n267), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n226), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT91), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT28), .Z(new_n671));
  NAND2_X1  g0471(.A1(new_n631), .A2(new_n653), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(KEYINPUT29), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT29), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n530), .A2(new_n488), .A3(new_n619), .ZN(new_n675));
  INV_X1    g0475(.A(new_n498), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n497), .B1(new_n496), .B2(new_n493), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n675), .B1(new_n678), .B2(new_n639), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n622), .A2(new_n610), .ZN(new_n680));
  INV_X1    g0480(.A(new_n606), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n619), .A2(new_n525), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n674), .B1(new_n684), .B2(new_n653), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n673), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n520), .A2(new_n483), .A3(new_n521), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n580), .A2(new_n474), .A3(new_n480), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n565), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT30), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n688), .A2(new_n485), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n489), .A3(new_n604), .A4(new_n557), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n653), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n608), .A2(new_n499), .A3(new_n531), .A4(new_n653), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(KEYINPUT31), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(KEYINPUT31), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n686), .B1(new_n687), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n671), .B1(new_n701), .B2(G1), .ZN(G364));
  INV_X1    g0502(.A(new_n666), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n640), .A2(G45), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n652), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(G330), .B2(new_n651), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n228), .A2(G190), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G179), .A2(G200), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT95), .Z(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n489), .A3(G200), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT93), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(G329), .A2(new_n713), .B1(new_n719), .B2(G283), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n228), .A2(new_n307), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n489), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n387), .B1(new_n724), .B2(G322), .ZN(new_n725));
  INV_X1    g0525(.A(G303), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n721), .A2(new_n489), .A3(G200), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G190), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G317), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(KEYINPUT33), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(KEYINPUT33), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n728), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n722), .A2(new_n709), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G311), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n228), .B1(new_n710), .B2(G190), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n729), .A2(new_n307), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n740), .A2(G294), .B1(G326), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT94), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n720), .A2(new_n735), .A3(new_n738), .A4(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n387), .B1(new_n736), .B2(new_n205), .ZN(new_n745));
  INV_X1    g0545(.A(new_n711), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G159), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT32), .ZN(new_n748));
  INV_X1    g0548(.A(new_n727), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n745), .B(new_n748), .C1(G87), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n739), .A2(new_n211), .ZN(new_n751));
  INV_X1    g0551(.A(new_n741), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n203), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n751), .B(new_n753), .C1(G68), .C2(new_n730), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n723), .B(KEYINPUT92), .Z(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n750), .B(new_n754), .C1(new_n215), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n718), .A2(new_n389), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n744), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n227), .B1(G20), .B2(new_n313), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n760), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n248), .A2(G45), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n665), .A2(new_n387), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n765), .B(new_n766), .C1(G45), .C2(new_n225), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n387), .A2(G355), .A3(new_n232), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(G116), .C2(new_n232), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n759), .A2(new_n760), .B1(new_n764), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n763), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n651), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n708), .B1(new_n705), .B2(new_n772), .ZN(G396));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n712), .A2(new_n774), .B1(new_n718), .B2(new_n585), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n752), .A2(new_n726), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n294), .B1(new_n736), .B2(new_n251), .C1(new_n727), .C2(new_n389), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n775), .A2(new_n751), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G294), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n778), .B1(new_n779), .B2(new_n782), .C1(new_n783), .C2(new_n723), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n730), .A2(G150), .B1(new_n741), .B2(G137), .ZN(new_n785));
  INV_X1    g0585(.A(G159), .ZN(new_n786));
  INV_X1    g0586(.A(G143), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n785), .B1(new_n786), .B2(new_n736), .C1(new_n756), .C2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT34), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n789), .B1(new_n215), .B2(new_n739), .C1(new_n209), .C2(new_n718), .ZN(new_n790));
  INV_X1    g0590(.A(G132), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n387), .B1(new_n203), .B2(new_n727), .C1(new_n712), .C2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n784), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n760), .A2(new_n761), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(new_n760), .B1(new_n205), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n386), .A2(new_n646), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n443), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n396), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n397), .A2(new_n646), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n795), .B(new_n706), .C1(new_n762), .C2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n672), .B(new_n800), .Z(new_n802));
  NOR2_X1   g0602(.A1(new_n699), .A2(new_n687), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n802), .B(new_n803), .Z(new_n804));
  OAI21_X1  g0604(.A(new_n801), .B1(new_n804), .B2(new_n706), .ZN(G384));
  XNOR2_X1  g0605(.A(new_n644), .B(KEYINPUT99), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n347), .A2(new_n349), .B1(new_n326), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(KEYINPUT37), .B1(new_n372), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT101), .ZN(new_n809));
  OR3_X1    g0609(.A1(new_n372), .A2(new_n807), .A3(KEYINPUT37), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT101), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n811), .B(KEYINPUT37), .C1(new_n372), .C2(new_n807), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT102), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n806), .B1(new_n347), .B2(new_n349), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n375), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT102), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n809), .A2(new_n810), .A3(new_n817), .A4(new_n812), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT103), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT39), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  INV_X1    g0625(.A(new_n372), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n345), .A2(KEYINPUT16), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n349), .B1(new_n357), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n644), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n359), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n825), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n372), .A2(new_n807), .A3(KEYINPUT37), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n828), .A2(new_n829), .ZN(new_n835));
  OAI211_X1 g0635(.A(KEYINPUT38), .B(new_n834), .C1(new_n376), .C2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n819), .A2(KEYINPUT103), .A3(new_n820), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n823), .A2(new_n824), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n835), .B1(new_n361), .B2(new_n374), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n820), .B1(new_n839), .B2(new_n833), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(new_n824), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n634), .A2(new_n653), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n631), .A2(new_n653), .A3(new_n800), .ZN(new_n846));
  INV_X1    g0646(.A(new_n799), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n426), .A2(new_n646), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n433), .A2(new_n849), .A3(new_n441), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n415), .A2(G169), .A3(new_n439), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n852), .B(new_n434), .C1(new_n435), .C2(new_n436), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n430), .B2(new_n432), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT98), .B1(new_n854), .B2(new_n850), .ZN(new_n855));
  INV_X1    g0655(.A(new_n432), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT74), .B1(new_n431), .B2(new_n417), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n441), .B(new_n850), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n851), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n848), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n806), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n862), .A2(new_n841), .B1(new_n361), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT100), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n843), .A2(new_n845), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n445), .B1(new_n673), .B2(new_n685), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n637), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n868), .B(new_n870), .Z(new_n871));
  NAND3_X1  g0671(.A1(new_n823), .A2(new_n836), .A3(new_n837), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n697), .B(KEYINPUT104), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n873), .A2(new_n696), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n860), .A2(new_n799), .A3(new_n798), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n872), .A2(new_n875), .A3(KEYINPUT40), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n861), .B(new_n800), .C1(new_n873), .C2(new_n696), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(new_n841), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n445), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n881), .B(new_n882), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(G330), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n871), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n267), .B2(new_n640), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n251), .B1(new_n505), .B2(KEYINPUT35), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n229), .C1(KEYINPUT35), .C2(new_n505), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT36), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n225), .A2(new_n205), .A3(new_n338), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n203), .B2(G68), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n891), .A2(new_n267), .A3(G13), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT97), .Z(new_n893));
  NAND3_X1  g0693(.A1(new_n886), .A2(new_n889), .A3(new_n893), .ZN(G367));
  NAND2_X1  g0694(.A1(new_n512), .A2(new_n646), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n531), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n525), .A2(new_n653), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n661), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT42), .Z(new_n900));
  NAND3_X1  g0700(.A1(new_n678), .A2(new_n531), .A3(new_n895), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(new_n525), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n646), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n614), .A2(new_n646), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n618), .A2(new_n606), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n606), .B2(new_n904), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n898), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n659), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n903), .B(new_n907), .C1(new_n659), .C2(new_n909), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT105), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n704), .A2(G1), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n666), .B(KEYINPUT41), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n663), .A2(new_n898), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT45), .Z(new_n921));
  NOR2_X1   g0721(.A1(new_n663), .A2(new_n898), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(new_n652), .A3(new_n658), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n658), .B(new_n660), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n652), .B(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n700), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n659), .A3(new_n923), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n919), .B1(new_n930), .B2(new_n701), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n916), .B1(new_n917), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT106), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT106), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n916), .B(new_n934), .C1(new_n917), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n294), .B1(new_n711), .B2(new_n732), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n755), .B2(G303), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n211), .B2(new_n718), .C1(new_n779), .C2(new_n736), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n740), .A2(G107), .B1(G311), .B2(new_n741), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n782), .B2(new_n783), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n727), .A2(new_n251), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT46), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n939), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n749), .A2(G58), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n739), .A2(new_n209), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n741), .B2(G143), .ZN(new_n947));
  INV_X1    g0747(.A(G137), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n947), .B(new_n387), .C1(new_n948), .C2(new_n711), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G150), .A2(new_n724), .B1(new_n737), .B2(G50), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n718), .B2(new_n205), .ZN(new_n951));
  INV_X1    g0751(.A(new_n782), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n949), .B(new_n951), .C1(new_n952), .C2(G159), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n944), .B1(new_n945), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT47), .Z(new_n955));
  AOI21_X1  g0755(.A(new_n705), .B1(new_n955), .B2(new_n760), .ZN(new_n956));
  INV_X1    g0756(.A(new_n766), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n764), .B1(new_n232), .B2(new_n383), .C1(new_n239), .C2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n906), .A2(new_n771), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n936), .A2(new_n960), .ZN(G387));
  XOR2_X1   g0761(.A(KEYINPUT110), .B(G322), .Z(new_n962));
  AOI22_X1  g0762(.A1(new_n755), .A2(G317), .B1(new_n741), .B2(new_n962), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n726), .B2(new_n736), .C1(new_n782), .C2(new_n774), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT48), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n727), .A2(new_n783), .B1(new_n739), .B2(new_n779), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT109), .Z(new_n967));
  AND2_X1   g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT49), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n746), .A2(G326), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(KEYINPUT49), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n387), .B1(new_n719), .B2(G116), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n257), .A2(new_n731), .B1(new_n209), .B2(new_n736), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT108), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n749), .A2(G77), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n739), .A2(new_n383), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n741), .B2(G159), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n387), .B1(new_n711), .B2(new_n259), .C1(new_n203), .C2(new_n723), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n719), .B2(G97), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n975), .A2(new_n976), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n381), .A2(new_n203), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT50), .Z(new_n984));
  INV_X1    g0784(.A(G45), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n667), .B1(G68), .B2(G77), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n766), .C1(new_n985), .C2(new_n244), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n387), .A2(new_n667), .A3(new_n232), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G107), .C2(new_n232), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT107), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(KEYINPUT107), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n992), .A2(new_n763), .A3(new_n760), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n982), .A2(new_n760), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n994), .B(new_n706), .C1(new_n658), .C2(new_n771), .ZN(new_n995));
  INV_X1    g0795(.A(new_n917), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n928), .A2(new_n703), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT111), .Z(new_n998));
  AND2_X1   g0798(.A1(new_n927), .A2(new_n700), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n995), .B1(new_n996), .B2(new_n927), .C1(new_n998), .C2(new_n999), .ZN(G393));
  NAND3_X1  g0800(.A1(new_n925), .A2(KEYINPUT112), .A3(new_n929), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(KEYINPUT112), .B2(new_n925), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n666), .B(new_n930), .C1(new_n1002), .C2(new_n928), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n909), .A2(new_n763), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n764), .B1(new_n211), .B2(new_n232), .C1(new_n252), .C2(new_n957), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n739), .A2(new_n205), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n387), .B1(new_n711), .B2(new_n787), .C1(new_n727), .C2(new_n209), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n381), .C2(new_n737), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G50), .A2(new_n952), .B1(new_n719), .B2(G87), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n752), .A2(new_n259), .B1(new_n723), .B2(new_n786), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT51), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT113), .Z(new_n1013));
  INV_X1    g0813(.A(new_n962), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n294), .B1(new_n727), .B2(new_n779), .C1(new_n1014), .C2(new_n711), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1015), .B(new_n758), .C1(G116), .C2(new_n740), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n783), .B2(new_n736), .C1(new_n726), .C2(new_n782), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n724), .A2(G311), .B1(G317), .B2(new_n741), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT52), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1013), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n705), .B1(new_n1020), .B2(new_n760), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n1004), .A2(new_n1005), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n1002), .B2(new_n917), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1003), .A2(new_n1023), .ZN(G390));
  AOI21_X1  g0824(.A(new_n705), .B1(new_n257), .B2(new_n794), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT117), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n294), .B1(new_n723), .B2(new_n251), .C1(new_n585), .C2(new_n727), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n752), .A2(new_n779), .B1(new_n739), .B2(new_n205), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n782), .B2(new_n389), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G294), .A2(new_n713), .B1(new_n719), .B2(G68), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1030), .B1(new_n1032), .B2(KEYINPUT118), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(KEYINPUT118), .B2(new_n1032), .C1(new_n211), .C2(new_n736), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n723), .A2(new_n791), .ZN(new_n1035));
  INV_X1    g0835(.A(G128), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n752), .A2(new_n1036), .B1(new_n739), .B2(new_n786), .ZN(new_n1037));
  XOR2_X1   g0837(.A(KEYINPUT54), .B(G143), .Z(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n387), .B1(new_n1039), .B2(new_n736), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(new_n952), .C2(G137), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT53), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n727), .B2(new_n259), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n749), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n713), .A2(G125), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1041), .B(new_n1045), .C1(new_n203), .C2(new_n718), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1034), .B1(new_n1035), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1026), .B1(new_n1047), .B2(new_n760), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT119), .Z(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n843), .B2(new_n762), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT120), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n862), .A2(new_n844), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n838), .A3(new_n842), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT114), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n851), .C1(new_n855), .C2(new_n859), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n798), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n684), .A2(new_n653), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n847), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n872), .A3(new_n844), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1053), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n800), .A2(G330), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n861), .B(new_n1065), .C1(new_n873), .C2(new_n696), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n861), .B(new_n1065), .C1(new_n696), .C2(new_n698), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1053), .A2(new_n1062), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1051), .B1(new_n917), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n445), .B(G330), .C1(new_n873), .C2(new_n696), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n869), .A2(new_n1073), .A3(new_n637), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n695), .A2(KEYINPUT31), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n694), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1064), .B1(new_n1077), .B2(new_n697), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1066), .B1(new_n1078), .B2(new_n861), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n848), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1060), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n873), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1064), .B1(new_n1082), .B2(new_n1077), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1081), .B(new_n1068), .C1(new_n1083), .C2(new_n1057), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1074), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1071), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(KEYINPUT115), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT115), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1053), .A2(new_n1062), .A3(new_n1069), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1066), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1085), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n703), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1085), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1093), .A2(KEYINPUT116), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT116), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1072), .B1(new_n1096), .B2(new_n1097), .ZN(G378));
  XOR2_X1   g0898(.A(new_n1074), .B(KEYINPUT123), .Z(new_n1099));
  AOI21_X1  g0899(.A(new_n1088), .B1(new_n1071), .B2(new_n1085), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1092), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n311), .A2(new_n380), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n275), .A2(new_n829), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT55), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT56), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n877), .A2(G330), .A3(new_n880), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n866), .A2(new_n867), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n866), .B2(new_n867), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1108), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n868), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1107), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n866), .A2(new_n867), .A3(new_n1108), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1102), .A2(KEYINPUT57), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n666), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT124), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT57), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1102), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1117), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1118), .A2(KEYINPUT124), .A3(new_n666), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1121), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1124), .A2(new_n996), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1114), .A2(new_n761), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n794), .A2(new_n203), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n749), .A2(new_n1038), .B1(new_n724), .B2(G128), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT122), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n741), .A2(G125), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n948), .B2(new_n736), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G150), .B2(new_n740), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1132), .B(new_n1135), .C1(new_n791), .C2(new_n731), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT59), .Z(new_n1137));
  AOI21_X1  g0937(.A(G41), .B1(new_n719), .B2(G159), .ZN(new_n1138));
  AOI21_X1  g0938(.A(G33), .B1(new_n746), .B2(G124), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n719), .A2(G58), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT121), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n976), .B1(new_n389), .B2(new_n723), .C1(new_n383), .C2(new_n736), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n712), .A2(new_n779), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1143), .A2(new_n1144), .A3(G41), .A4(new_n387), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n752), .A2(new_n251), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n946), .B(new_n1146), .C1(G97), .C2(new_n730), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT58), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n203), .B1(new_n292), .B2(G41), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1140), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n705), .B1(new_n1151), .B2(new_n760), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1129), .A2(new_n1130), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1128), .A2(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1127), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(G375));
  NAND3_X1  g0957(.A1(new_n1080), .A2(new_n1084), .A3(new_n1074), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1094), .A2(new_n918), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n996), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1054), .A2(new_n761), .A3(new_n1056), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n712), .A2(new_n726), .B1(new_n718), .B2(new_n205), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n752), .A2(new_n783), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n294), .B1(new_n723), .B2(new_n779), .C1(new_n211), .C2(new_n727), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1162), .A2(new_n977), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n389), .B2(new_n736), .C1(new_n251), .C2(new_n782), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n756), .A2(new_n948), .B1(new_n712), .B2(new_n1036), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n752), .A2(new_n791), .B1(new_n739), .B2(new_n203), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n387), .B1(new_n736), .B2(new_n259), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n1142), .C1(new_n782), .C2(new_n1039), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n727), .A2(new_n786), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1166), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1173), .A2(new_n760), .B1(new_n209), .B2(new_n794), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1161), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1160), .B1(new_n706), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1159), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT125), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1159), .A2(KEYINPUT125), .A3(new_n1176), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(G381));
  NAND2_X1  g0981(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1182), .A2(new_n1072), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1156), .A2(new_n1183), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n960), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1186), .B(G390), .C1(new_n933), .C2(new_n935), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(G407));
  INV_X1    g0988(.A(G213), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1184), .B2(new_n645), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(G407), .ZN(G409));
  INV_X1    g0991(.A(KEYINPUT127), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(G387), .A2(G390), .ZN(new_n1193));
  INV_X1    g0993(.A(G390), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n936), .A2(new_n960), .A3(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(G393), .B(G396), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  XOR2_X1   g0997(.A(G393), .B(G396), .Z(new_n1198));
  AOI21_X1  g0998(.A(new_n1194), .B1(new_n936), .B2(new_n960), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1187), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1189), .A2(G343), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1127), .A2(G378), .A3(new_n1155), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT126), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1128), .B2(new_n1154), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1102), .A2(new_n918), .A3(new_n1117), .ZN(new_n1207));
  OAI211_X1 g1007(.A(KEYINPUT126), .B(new_n1153), .C1(new_n1124), .C2(new_n996), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1183), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1203), .B1(new_n1204), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT62), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT60), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n703), .B1(new_n1158), .B2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1214), .B(new_n1094), .C1(new_n1213), .C2(new_n1158), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(G384), .A3(new_n1176), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G384), .B1(new_n1215), .B2(new_n1176), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1211), .A2(new_n1212), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1212), .B1(new_n1211), .B2(new_n1219), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1203), .A2(G2897), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1219), .B(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1204), .A2(new_n1210), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1203), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(KEYINPUT61), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1202), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1211), .A2(new_n1219), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT63), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1219), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1203), .B(new_n1233), .C1(new_n1204), .C2(new_n1210), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1201), .B1(new_n1234), .B2(KEYINPUT63), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1232), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1192), .B1(new_n1229), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1232), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1220), .A2(new_n1221), .A3(KEYINPUT61), .A4(new_n1227), .ZN(new_n1240));
  OAI211_X1 g1040(.A(KEYINPUT127), .B(new_n1239), .C1(new_n1240), .C2(new_n1202), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(G405));
  NAND2_X1  g1042(.A1(G375), .A2(new_n1183), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1204), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(new_n1202), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(new_n1233), .ZN(G402));
endmodule


