//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G227), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT10), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n195), .A3(G143), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n197), .B(new_n199), .C1(G143), .C2(new_n195), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G128), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n194), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n209), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT79), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT80), .B(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G104), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT81), .B(G101), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n209), .A2(G107), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n216), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n214), .B1(new_n222), .B2(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G101), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n226), .A2(KEYINPUT82), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT82), .B1(new_n226), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n208), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT11), .ZN(new_n232));
  INV_X1    g046(.A(G134), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G137), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(KEYINPUT65), .B(new_n232), .C1(new_n233), .C2(G137), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .A3(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n233), .A2(G137), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n238), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n239), .B1(new_n238), .B2(new_n243), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT83), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n247));
  INV_X1    g061(.A(new_n237), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n240), .A2(G134), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT65), .B1(new_n249), .B2(new_n232), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n243), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G131), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n238), .A2(new_n239), .A3(new_n243), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n216), .A2(new_n225), .ZN(new_n257));
  INV_X1    g071(.A(new_n223), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n256), .B(G101), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n200), .A2(new_n262), .B1(new_n205), .B2(new_n260), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n226), .A2(KEYINPUT4), .ZN(new_n264));
  INV_X1    g078(.A(G101), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n212), .A2(new_n215), .B1(new_n209), .B2(G107), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n223), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n259), .B(new_n263), .C1(new_n264), .C2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n207), .B1(new_n202), .B2(new_n205), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n226), .A2(new_n228), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n194), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n231), .A2(new_n255), .A3(new_n268), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n200), .A2(new_n262), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n205), .A2(new_n260), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n256), .B2(new_n267), .ZN(new_n278));
  OAI21_X1  g092(.A(G101), .B1(new_n257), .B2(new_n258), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n278), .A2(new_n280), .B1(new_n194), .B2(new_n270), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n281), .A2(KEYINPUT84), .A3(new_n231), .A4(new_n255), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n193), .B1(new_n274), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n231), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n252), .A2(new_n253), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n204), .A2(new_n207), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n229), .A2(new_n230), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n270), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT12), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT12), .B(new_n285), .C1(new_n289), .C2(new_n290), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n274), .A2(new_n282), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT85), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n287), .B1(new_n301), .B2(new_n193), .ZN(new_n302));
  OAI21_X1  g116(.A(G469), .B1(new_n302), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT86), .B(G469), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n283), .A2(new_n295), .ZN(new_n307));
  INV_X1    g121(.A(new_n193), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n296), .B2(new_n286), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n304), .B(new_n306), .C1(new_n307), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n283), .A2(new_n295), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n315), .A2(KEYINPUT87), .A3(new_n304), .A4(new_n306), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n189), .B1(new_n303), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G214), .B1(G237), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT91), .B1(new_n288), .B2(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n277), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT91), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n204), .A2(new_n323), .A3(new_n324), .A4(new_n207), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G953), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G224), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT7), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  MUX2_X1   g144(.A(new_n263), .B(new_n288), .S(new_n324), .Z(new_n331));
  INV_X1    g145(.A(new_n328), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(KEYINPUT92), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT7), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n332), .B2(KEYINPUT92), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G116), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G119), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT68), .B(G116), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(G119), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT5), .ZN(new_n342));
  INV_X1    g156(.A(G113), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT88), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT2), .B(G113), .Z(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT88), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n350), .A3(new_n345), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n230), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n226), .A2(KEYINPUT82), .A3(new_n228), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n341), .B(new_n348), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n280), .A2(new_n356), .A3(new_n259), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G110), .B(G122), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT89), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n337), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n361), .B(KEYINPUT8), .Z(new_n364));
  INV_X1    g178(.A(new_n352), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n228), .B2(new_n226), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n353), .A2(new_n354), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n367), .A2(new_n349), .A3(new_n346), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n364), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(G902), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n361), .B1(new_n355), .B2(new_n358), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n367), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n362), .A3(new_n357), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n373), .A3(KEYINPUT6), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n375), .B(new_n361), .C1(new_n355), .C2(new_n358), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n328), .B(KEYINPUT90), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n331), .B(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G210), .B1(G237), .B2(G902), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n370), .A2(new_n379), .A3(new_n381), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n320), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n327), .A3(G214), .ZN(new_n387));
  INV_X1    g201(.A(G143), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G131), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n387), .B(G143), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n239), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT17), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n324), .B2(KEYINPUT73), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT73), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(G125), .A3(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT16), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n324), .B2(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(new_n195), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n394), .B(new_n403), .C1(new_n393), .C2(new_n390), .ZN(new_n404));
  XNOR2_X1  g218(.A(G113), .B(G122), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(new_n209), .ZN(new_n406));
  AND2_X1   g220(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G131), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n195), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n396), .A2(G146), .A3(new_n398), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n391), .A2(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT94), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n389), .A2(G131), .A3(new_n407), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n412), .B2(new_n414), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n404), .B(new_n406), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n417), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n415), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n406), .B1(new_n421), .B2(new_n404), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n304), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G475), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT19), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n409), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n396), .A2(KEYINPUT19), .A3(new_n398), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n195), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT95), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n390), .A2(new_n392), .B1(G146), .B2(new_n402), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n420), .A2(new_n415), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT96), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n406), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n421), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT96), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n419), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(G475), .A2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n437), .A2(KEYINPUT20), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n431), .A2(new_n432), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n434), .B(new_n432), .C1(new_n416), .C2(new_n417), .ZN(new_n443));
  INV_X1    g257(.A(new_n406), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n418), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n441), .B1(new_n446), .B2(new_n438), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n424), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G217), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n187), .A2(new_n449), .A3(G953), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G128), .B(G143), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n452), .A2(KEYINPUT13), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n388), .A2(G128), .ZN(new_n454));
  OAI21_X1  g268(.A(G134), .B1(new_n454), .B2(KEYINPUT13), .ZN(new_n455));
  OR3_X1    g269(.A1(new_n453), .A2(KEYINPUT98), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT98), .B1(new_n453), .B2(new_n455), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n233), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n458), .A2(KEYINPUT99), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(KEYINPUT99), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(new_n457), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT97), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n340), .A2(G122), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n338), .A2(G122), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n462), .A3(new_n464), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n222), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n222), .ZN(new_n469));
  INV_X1    g283(.A(new_n467), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n465), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n461), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n468), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n452), .B(new_n233), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n463), .A2(new_n475), .A3(new_n464), .ZN(new_n476));
  OAI21_X1  g290(.A(G107), .B1(new_n463), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n451), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n471), .A2(new_n468), .ZN(new_n481));
  OAI221_X1 g295(.A(new_n450), .B1(new_n473), .B2(new_n478), .C1(new_n481), .C2(new_n461), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G478), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT100), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n483), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n448), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(G234), .A2(G237), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(G952), .A3(new_n327), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(G902), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(new_n327), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n385), .A2(new_n491), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n318), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n402), .B(G146), .ZN(new_n502));
  XNOR2_X1  g316(.A(G119), .B(G128), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT72), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT24), .B(G110), .Z(new_n506));
  INV_X1    g320(.A(G119), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G128), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n507), .A2(G128), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(KEYINPUT23), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n505), .A2(new_n506), .B1(G110), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n502), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT74), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n402), .A2(G146), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n505), .A2(new_n506), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n511), .A2(G110), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n515), .B(new_n410), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT22), .B(G137), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT75), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT76), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n327), .A2(G221), .A3(G234), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n514), .A2(new_n524), .A3(new_n518), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT77), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT77), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n449), .B1(G234), .B2(new_n304), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G902), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n527), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n524), .B1(new_n514), .B2(new_n518), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n304), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT25), .B1(new_n528), .B2(new_n304), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n533), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n249), .A2(new_n242), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G131), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n288), .A2(new_n545), .A3(new_n253), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n263), .B1(new_n244), .B2(new_n245), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT30), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n356), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n288), .A2(new_n545), .A3(new_n253), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT66), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT66), .B(new_n263), .C1(new_n244), .C2(new_n245), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n556), .A2(KEYINPUT67), .A3(KEYINPUT30), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT67), .ZN(new_n558));
  INV_X1    g372(.A(new_n555), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT66), .B1(new_n285), .B2(new_n263), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n546), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n551), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n356), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n548), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n567));
  INV_X1    g381(.A(G210), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n568), .A2(G237), .A3(G953), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n567), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT26), .B(G101), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n570), .B(new_n571), .Z(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n564), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT67), .B1(new_n556), .B2(KEYINPUT30), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n561), .A2(new_n558), .A3(new_n562), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n550), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT31), .B1(new_n579), .B2(new_n573), .ZN(new_n580));
  INV_X1    g394(.A(new_n572), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n566), .A2(KEYINPUT28), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT28), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n548), .A2(new_n583), .A3(new_n565), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n556), .A2(new_n565), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n581), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n576), .A2(new_n580), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(G472), .A2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT32), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT32), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n566), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n579), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n581), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n572), .B1(new_n586), .B2(new_n587), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT29), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n585), .B1(new_n565), .B2(new_n548), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n572), .A2(KEYINPUT29), .ZN(new_n602));
  OAI211_X1 g416(.A(KEYINPUT71), .B(new_n304), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT71), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n548), .A2(new_n565), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n605), .B(new_n602), .C1(new_n582), .C2(new_n584), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n606), .B2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n543), .B1(new_n595), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n501), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n224), .ZN(G3));
  NAND2_X1  g427(.A1(new_n589), .A2(new_n304), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G472), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n591), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n543), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n318), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT101), .ZN(new_n619));
  INV_X1    g433(.A(new_n384), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n381), .B1(new_n370), .B2(new_n379), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n319), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n480), .A2(new_n482), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT33), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n480), .A2(new_n482), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(G478), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n484), .A2(new_n304), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n483), .B2(new_n484), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n448), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n622), .A2(new_n498), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n619), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(new_n448), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n490), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n637), .A2(new_n622), .A3(new_n498), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n619), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n538), .A2(new_n539), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n528), .A2(KEYINPUT25), .A3(new_n304), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n519), .A2(KEYINPUT36), .A3(new_n524), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n525), .A2(new_n647), .B1(new_n514), .B2(new_n518), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n645), .A2(new_n533), .B1(new_n534), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n642), .B1(new_n616), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n534), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n542), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n615), .A2(new_n653), .A3(KEYINPUT102), .A4(new_n591), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n501), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT37), .B(G110), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(new_n594), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n593), .B1(new_n589), .B2(new_n590), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n609), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n318), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT20), .B1(new_n437), .B2(new_n439), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n446), .A2(new_n441), .A3(new_n438), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G953), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n495), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(KEYINPUT103), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(KEYINPUT103), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n669), .A2(new_n493), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n490), .A2(new_n665), .A3(new_n424), .A4(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n622), .A2(new_n650), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n662), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XOR2_X1   g490(.A(new_n671), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n318), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n597), .A2(new_n581), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n566), .A2(new_n581), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n304), .B1(new_n682), .B2(new_n605), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n595), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n383), .A2(new_n384), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT105), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n687), .B(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n489), .B1(new_n665), .B2(new_n424), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n650), .A2(new_n319), .A3(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n686), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n679), .A2(new_n680), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND3_X1  g509(.A1(new_n448), .A2(new_n630), .A3(new_n672), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n622), .A2(new_n650), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n662), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  INV_X1    g513(.A(new_n315), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n317), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n189), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n610), .A3(new_n632), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n610), .A3(new_n638), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND4_X1  g522(.A1(new_n661), .A2(new_n491), .A3(new_n499), .A4(new_n653), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n317), .A2(new_n188), .A3(new_n701), .A4(new_n385), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  AND2_X1   g526(.A1(new_n535), .A2(new_n542), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n601), .A2(new_n581), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n576), .A2(new_n580), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n590), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT106), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(new_n718), .A3(new_n590), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n713), .A2(new_n720), .A3(new_n615), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n687), .A2(new_n319), .A3(new_n691), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n498), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n703), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  AND3_X1   g540(.A1(new_n715), .A2(new_n718), .A3(new_n590), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n718), .B1(new_n715), .B2(new_n590), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n615), .B(new_n653), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n696), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n188), .A2(new_n317), .A3(new_n385), .A4(new_n701), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n696), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n720), .A2(new_n615), .A3(new_n653), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(new_n735), .B2(new_n710), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(G469), .A2(G902), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT108), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n302), .B2(G469), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n317), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n687), .A2(new_n189), .A3(new_n320), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n610), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n739), .B1(new_n745), .B2(new_n696), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n610), .A3(KEYINPUT42), .A4(new_n734), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  OR2_X1    g564(.A1(new_n745), .A2(new_n673), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NAND2_X1  g566(.A1(new_n636), .A2(new_n630), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT43), .Z(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n616), .A3(new_n653), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(KEYINPUT44), .A3(new_n616), .A4(new_n653), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n687), .A2(new_n320), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(KEYINPUT109), .A3(new_n758), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n302), .A2(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n302), .A2(KEYINPUT45), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(G469), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n741), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n769), .A2(new_n770), .B1(new_n312), .B2(new_n316), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n188), .A3(new_n677), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n764), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  INV_X1    g589(.A(new_n759), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n661), .A2(new_n776), .A3(new_n713), .A4(new_n696), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT47), .B1(new_n772), .B2(new_n188), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n783));
  INV_X1    g597(.A(new_n780), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n317), .A2(new_n189), .A3(new_n701), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n778), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n754), .A2(new_n722), .A3(new_n494), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n776), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n702), .A2(new_n776), .A3(new_n189), .A4(new_n493), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n754), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n729), .ZN(new_n793));
  INV_X1    g607(.A(new_n788), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n703), .A2(new_n690), .A3(new_n320), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT50), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n793), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n686), .A2(new_n713), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n791), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n791), .A3(KEYINPUT115), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n448), .A2(new_n630), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n800), .A2(KEYINPUT116), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n790), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n787), .B1(new_n786), .B2(new_n789), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n783), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n792), .A2(new_n611), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT48), .Z(new_n817));
  INV_X1    g631(.A(G952), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n818), .B(G953), .C1(new_n794), .C2(new_n731), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n805), .A2(new_n806), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n817), .B(new_n819), .C1(new_n631), .C2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n786), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n784), .A2(new_n778), .A3(KEYINPUT117), .A4(new_n785), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n789), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n809), .A2(new_n783), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n821), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n732), .B1(new_n730), .B2(new_n731), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n735), .A2(KEYINPUT107), .A3(new_n710), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n318), .B(new_n661), .C1(new_n674), .C2(new_n697), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n723), .B1(new_n595), .B2(new_n684), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n542), .A2(new_n188), .A3(new_n652), .A4(new_n672), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n742), .B2(new_n317), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(KEYINPUT112), .B(new_n834), .C1(new_n742), .C2(new_n317), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n828), .B1(new_n831), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n742), .A2(new_n317), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT112), .B1(new_n841), .B2(new_n834), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n835), .A2(new_n836), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n833), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n737), .A3(KEYINPUT52), .A4(new_n832), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n840), .A2(KEYINPUT113), .A3(new_n845), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n749), .A2(new_n751), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n491), .A2(new_n759), .A3(new_n653), .A4(new_n672), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n662), .A2(new_n852), .B1(new_n747), .B2(new_n730), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n703), .B(new_n610), .C1(new_n632), .C2(new_n638), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n711), .A3(new_n725), .A4(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n318), .A2(new_n617), .A3(new_n632), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n501), .B2(new_n611), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n318), .A2(new_n617), .A3(new_n638), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n655), .B2(new_n501), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT110), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(KEYINPUT110), .B(new_n859), .C1(new_n655), .C2(new_n501), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n862), .A2(KEYINPUT111), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT111), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT53), .B1(new_n850), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n711), .A2(new_n725), .A3(new_n854), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n749), .A3(new_n751), .A4(new_n853), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n860), .A2(new_n861), .ZN(new_n870));
  INV_X1    g684(.A(new_n858), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n863), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT111), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n862), .A2(KEYINPUT111), .A3(new_n863), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n846), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n867), .A2(new_n878), .A3(KEYINPUT54), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n850), .B2(new_n866), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT54), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n815), .A2(new_n827), .A3(new_n879), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n702), .A2(KEYINPUT49), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n543), .A2(new_n753), .A3(new_n189), .A4(new_n320), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n702), .A2(KEYINPUT49), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n686), .A3(new_n889), .A4(new_n690), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n886), .B1(new_n887), .B2(new_n890), .ZN(G75));
  NAND2_X1  g705(.A1(new_n818), .A2(G953), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT120), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n876), .A2(new_n882), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n304), .B1(new_n880), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n374), .A2(new_n376), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT118), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n378), .B(KEYINPUT55), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n893), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n840), .A2(KEYINPUT113), .A3(new_n845), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT113), .B1(new_n840), .B2(new_n845), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT53), .B1(new_n905), .B2(new_n876), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n866), .A2(new_n881), .ZN(new_n907));
  OAI21_X1  g721(.A(G902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n902), .B(new_n900), .C1(new_n908), .C2(new_n568), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n896), .A2(KEYINPUT119), .A3(new_n900), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n901), .B1(new_n911), .B2(new_n912), .ZN(G51));
  INV_X1    g727(.A(new_n893), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n866), .B2(new_n881), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n906), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n906), .B2(new_n907), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n880), .A2(KEYINPUT121), .A3(new_n883), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n741), .B(KEYINPUT57), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n315), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n908), .A2(new_n767), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n914), .B1(new_n924), .B2(new_n925), .ZN(G54));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  AND2_X1   g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n895), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n929), .B2(new_n437), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n914), .B1(new_n929), .B2(new_n437), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n895), .A2(KEYINPUT122), .A3(new_n446), .A4(new_n928), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G60));
  XNOR2_X1  g747(.A(new_n628), .B(KEYINPUT59), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n879), .B2(new_n884), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n624), .A2(new_n626), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n893), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n934), .B1(new_n624), .B2(new_n626), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n921), .B2(new_n938), .ZN(G63));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n893), .B1(new_n940), .B2(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n880), .B2(new_n894), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n944), .B2(new_n649), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n946));
  INV_X1    g760(.A(new_n532), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n906), .A2(new_n907), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n943), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n946), .B1(new_n945), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  INV_X1    g766(.A(new_n497), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n327), .B1(new_n953), .B2(G224), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n868), .B1(new_n864), .B2(new_n865), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n327), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n898), .B1(G898), .B2(new_n327), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(G69));
  OAI21_X1  g772(.A(new_n549), .B1(new_n557), .B2(new_n563), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n426), .A2(new_n427), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n611), .A2(new_n723), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n772), .A2(new_n188), .A3(new_n677), .A4(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n737), .A2(new_n832), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n967), .A2(new_n749), .A3(new_n751), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n774), .A2(new_n966), .A3(new_n781), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n327), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n962), .B1(new_n970), .B2(new_n667), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n694), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n637), .A2(new_n631), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n759), .A3(new_n976), .ZN(new_n977));
  OR3_X1    g791(.A1(new_n977), .A2(new_n611), .A3(new_n678), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n973), .A2(new_n774), .A3(new_n781), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n961), .B1(new_n979), .B2(new_n327), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n327), .B1(G227), .B2(G900), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OR3_X1    g797(.A1(new_n971), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n971), .B2(new_n980), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n969), .B2(new_n955), .ZN(new_n989));
  INV_X1    g803(.A(new_n598), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n914), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n988), .B1(new_n979), .B2(new_n955), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n681), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n598), .A2(new_n988), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(new_n681), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n867), .A2(new_n878), .A3(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(KEYINPUT127), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n994), .B1(new_n998), .B2(new_n999), .ZN(G57));
endmodule


