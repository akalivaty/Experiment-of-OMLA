//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n206), .B1(new_n203), .B2(KEYINPUT15), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT87), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n204), .A2(new_n207), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT15), .B(new_n203), .C1(new_n213), .C2(new_n206), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT16), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G8gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n222), .A2(G1gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT89), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(G8gat), .B1(new_n222), .B2(new_n224), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT89), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n230), .B(new_n231), .C1(G1gat), .C2(new_n222), .ZN(new_n232));
  XOR2_X1   g031(.A(G15gat), .B(G22gat), .Z(new_n233));
  INV_X1    g032(.A(KEYINPUT88), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n223), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT88), .B1(new_n222), .B2(G1gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n225), .A3(new_n236), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n229), .A2(new_n232), .B1(new_n237), .B2(G8gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n217), .A2(KEYINPUT17), .A3(new_n218), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n229), .A2(new_n232), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(G8gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n219), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n202), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n219), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(KEYINPUT90), .A3(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n246), .B(KEYINPUT13), .Z(new_n252));
  OR3_X1    g051(.A1(new_n238), .A2(new_n249), .A3(KEYINPUT90), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n240), .A2(new_n244), .A3(KEYINPUT18), .A4(new_n246), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n248), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT86), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G197gat), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT11), .B(G169gat), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n256), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n256), .B2(new_n257), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT31), .B(G50gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n267), .B(G22gat), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(G211gat), .ZN(new_n271));
  INV_X1    g070(.A(G218gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n270), .B1(KEYINPUT22), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT74), .B(G141gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(G148gat), .ZN(new_n279));
  INV_X1    g078(.A(G148gat), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n280), .A2(G141gat), .ZN(new_n281));
  INV_X1    g080(.A(G155gat), .ZN(new_n282));
  INV_X1    g081(.A(G162gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n285));
  OAI22_X1  g084(.A1(new_n279), .A2(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G155gat), .B(G162gat), .Z(new_n287));
  XOR2_X1   g086(.A(KEYINPUT73), .B(KEYINPUT2), .Z(new_n288));
  XNOR2_X1  g087(.A(G141gat), .B(G148gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT75), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n286), .A2(new_n290), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT3), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n277), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n292), .B1(new_n276), .B2(KEYINPUT29), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n295), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT81), .ZN(new_n304));
  OAI211_X1 g103(.A(G228gat), .B(G233gat), .C1(new_n301), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n298), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n296), .A2(new_n297), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n276), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n295), .A2(KEYINPUT77), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n302), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT80), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n314), .A2(new_n315), .B1(G228gat), .B2(G233gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(KEYINPUT80), .A3(new_n302), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n309), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G78gat), .B(G106gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n319), .B(KEYINPUT79), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n305), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n321), .B1(new_n305), .B2(new_n318), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n269), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n318), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n320), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n305), .A2(new_n318), .A3(new_n321), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n268), .A3(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G169gat), .ZN(new_n332));
  INV_X1    g131(.A(G176gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT23), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(G169gat), .B2(G176gat), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT64), .B(G169gat), .Z(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT23), .A3(new_n333), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(G190gat), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT24), .ZN(new_n340));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(KEYINPUT24), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n335), .B(new_n337), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT25), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT65), .B(G183gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G190gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT66), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(new_n342), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT23), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n335), .A2(KEYINPUT25), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n346), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(KEYINPUT1), .ZN(new_n356));
  INV_X1    g155(.A(G127gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G134gat), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(KEYINPUT67), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G134gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G127gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n361), .B(new_n358), .C1(new_n356), .C2(KEYINPUT67), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT27), .B(G183gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(KEYINPUT28), .A3(new_n339), .ZN(new_n367));
  NOR2_X1   g166(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n347), .B2(KEYINPUT27), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(G190gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(new_n370), .B2(KEYINPUT28), .ZN(new_n371));
  NOR2_X1   g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(KEYINPUT26), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n332), .B2(new_n333), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(KEYINPUT26), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n371), .A2(new_n341), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n354), .A2(new_n365), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n365), .B1(new_n354), .B2(new_n376), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n331), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT32), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G15gat), .B(G43gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT68), .ZN(new_n384));
  INV_X1    g183(.A(G71gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n386), .B(G99gat), .Z(new_n387));
  NAND3_X1  g186(.A1(new_n380), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n379), .B(KEYINPUT32), .C1(new_n381), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n354), .A2(new_n376), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n363), .A2(new_n364), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n354), .A2(new_n365), .A3(new_n376), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n330), .A3(new_n395), .ZN(new_n396));
  XOR2_X1   g195(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n391), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n397), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n396), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(new_n388), .A3(new_n390), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n329), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT35), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT71), .ZN(new_n408));
  XNOR2_X1  g207(.A(G64gat), .B(G92gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n410), .B(KEYINPUT72), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT29), .B1(new_n354), .B2(new_n376), .ZN(new_n413));
  AND2_X1   g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n392), .A2(new_n414), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n277), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n416), .B(new_n277), .C1(new_n414), .C2(new_n413), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n412), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n413), .A2(new_n414), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n392), .A2(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n276), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(new_n418), .A3(new_n410), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n406), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n406), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT0), .ZN(new_n430));
  XNOR2_X1  g229(.A(G57gat), .B(G85gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT83), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT5), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n365), .A2(new_n291), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n393), .A2(new_n295), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT76), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n435), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n436), .A2(KEYINPUT4), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n311), .A2(new_n365), .A3(new_n312), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT4), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n445), .B2(KEYINPUT78), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT4), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n393), .B1(new_n291), .B2(new_n292), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n294), .B2(new_n298), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n440), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n442), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n436), .A2(KEYINPUT4), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n311), .A2(new_n365), .A3(new_n455), .A4(new_n312), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n435), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n434), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461));
  INV_X1    g260(.A(new_n432), .ZN(new_n462));
  INV_X1    g261(.A(new_n450), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n299), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n440), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n448), .B2(new_n446), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n458), .B(new_n462), .C1(new_n467), .C2(new_n442), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n460), .A2(new_n461), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT6), .B(new_n432), .C1(new_n453), .C2(new_n459), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT85), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n458), .B1(new_n467), .B2(new_n442), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT6), .A4(new_n432), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n404), .A2(new_n405), .A3(new_n428), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n468), .A2(new_n461), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n449), .A2(new_n452), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n441), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n462), .B1(new_n479), .B2(new_n458), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n470), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n402), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n401), .B1(new_n388), .B2(new_n390), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n324), .A2(new_n328), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n481), .A2(new_n484), .A3(new_n428), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n454), .A2(new_n456), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n440), .B(new_n489), .C1(new_n490), .C2(new_n451), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n465), .B1(new_n464), .B2(new_n457), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT39), .B1(new_n438), .B2(new_n440), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n491), .B(new_n433), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n434), .B1(new_n492), .B2(new_n489), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(KEYINPUT40), .C1(new_n492), .C2(new_n493), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n496), .A2(new_n460), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n424), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n411), .B1(new_n423), .B2(new_n418), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT30), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n426), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT37), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n423), .A2(new_n418), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n410), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n505), .B1(new_n423), .B2(new_n418), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT38), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT37), .B1(new_n417), .B2(new_n419), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n411), .A2(KEYINPUT38), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n506), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n424), .A3(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n504), .B(new_n485), .C1(new_n475), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n481), .A2(new_n428), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n324), .A2(new_n328), .A3(KEYINPUT82), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT82), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n485), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522));
  OAI22_X1  g321(.A1(new_n482), .A2(new_n483), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n399), .A2(new_n402), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n515), .A2(new_n520), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n266), .B1(new_n488), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G57gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT92), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G57gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n533), .A3(G64gat), .ZN(new_n534));
  INV_X1    g333(.A(G64gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G57gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT93), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT92), .B(G57gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(KEYINPUT93), .A3(G64gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT9), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT91), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT91), .B1(new_n542), .B2(new_n543), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n530), .A2(G64gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n544), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n548), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G127gat), .ZN(new_n562));
  XOR2_X1   g361(.A(G183gat), .B(G211gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n238), .B1(new_n558), .B2(new_n557), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT94), .Z(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n282), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n566), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n563), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n562), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT97), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT97), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n577), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT7), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(G85gat), .A3(G92gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(KEYINPUT8), .A2(new_n577), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n584), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n580), .A2(new_n583), .A3(new_n589), .A4(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n221), .A2(new_n239), .A3(new_n596), .ZN(new_n597));
  AND4_X1   g396(.A1(new_n580), .A2(new_n583), .A3(new_n589), .A4(new_n592), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n580), .A2(new_n583), .B1(new_n589), .B2(new_n592), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n219), .A2(new_n600), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n339), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n339), .B1(new_n597), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n272), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(G218gat), .A3(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT96), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT95), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G134gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G162gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT96), .A4(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n576), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n541), .A2(new_n550), .B1(new_n555), .B2(new_n548), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(new_n600), .ZN(new_n625));
  XNOR2_X1  g424(.A(G71gat), .B(G78gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n552), .A2(new_n626), .A3(new_n544), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n538), .B2(new_n540), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n555), .A2(new_n548), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n596), .B(KEYINPUT98), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT99), .B1(new_n557), .B2(new_n596), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n624), .A2(new_n600), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n635));
  NAND4_X1  g434(.A1(new_n631), .A2(new_n632), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n624), .A2(new_n600), .A3(KEYINPUT10), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n622), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(KEYINPUT101), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  AOI211_X1 g439(.A(new_n640), .B(new_n622), .C1(new_n636), .C2(new_n637), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n643), .A2(new_n622), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n638), .B2(new_n644), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n620), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n529), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n481), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n223), .ZN(G1324gat));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n226), .B1(new_n657), .B2(new_n503), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n654), .A2(new_n428), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(KEYINPUT42), .B2(new_n660), .ZN(G1325gat));
  NOR3_X1   g461(.A1(new_n654), .A2(G15gat), .A3(new_n403), .ZN(new_n663));
  INV_X1    g462(.A(new_n526), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n399), .A2(new_n402), .B1(KEYINPUT70), .B2(KEYINPUT36), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT102), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n523), .A2(new_n667), .A3(new_n526), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n657), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n663), .B1(G15gat), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT103), .Z(G1326gat));
  AND3_X1   g472(.A1(new_n324), .A2(new_n328), .A3(KEYINPUT82), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT82), .B1(new_n324), .B2(new_n328), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n654), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n652), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n575), .A2(new_n618), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT104), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n529), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G29gat), .A3(new_n481), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT45), .Z(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n619), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n515), .A2(new_n520), .A3(new_n527), .ZN(new_n689));
  AND4_X1   g488(.A1(new_n405), .A2(new_n484), .A3(new_n428), .A4(new_n485), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n690), .A2(new_n475), .B1(new_n486), .B2(KEYINPUT35), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT105), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT105), .B1(new_n570), .B2(new_n574), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(new_n266), .A3(new_n652), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n515), .A2(new_n520), .A3(new_n666), .A4(new_n668), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n619), .B1(new_n697), .B2(new_n488), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n692), .B(new_n696), .C1(new_n698), .C2(KEYINPUT44), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n481), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n686), .A2(new_n700), .ZN(G1328gat));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n209), .B1(new_n702), .B2(KEYINPUT106), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n684), .A2(new_n428), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(KEYINPUT106), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n699), .B2(new_n428), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1329gat));
  OAI21_X1  g507(.A(G43gat), .B1(new_n699), .B2(new_n669), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n403), .A2(G43gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n684), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g511(.A(G50gat), .B1(new_n699), .B2(new_n485), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n677), .A2(G50gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n529), .A2(new_n683), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(KEYINPUT48), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n717), .B(G50gat), .C1(new_n699), .C2(new_n677), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n715), .A2(KEYINPUT108), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n510), .A2(new_n424), .A3(new_n513), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n722), .A2(new_n471), .A3(new_n469), .A4(new_n474), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n329), .B1(new_n503), .B2(new_n499), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n723), .A2(new_n724), .B1(new_n676), .B2(new_n516), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n725), .A2(new_n669), .B1(new_n487), .B2(new_n476), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n687), .B1(new_n726), .B2(new_n619), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n727), .A2(new_n676), .A3(new_n692), .A4(new_n696), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n721), .B1(new_n728), .B2(G50gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n716), .B1(new_n720), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT109), .B(new_n716), .C1(new_n720), .C2(new_n729), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1331gat));
  NAND2_X1  g533(.A1(new_n697), .A2(new_n488), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n620), .A2(new_n265), .A3(new_n681), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n481), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n539), .ZN(G1332gat));
  NOR2_X1   g538(.A1(new_n737), .A2(new_n428), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT110), .ZN(G1333gat));
  NOR3_X1   g544(.A1(new_n737), .A2(G71gat), .A3(new_n403), .ZN(new_n746));
  INV_X1    g545(.A(new_n737), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n670), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n746), .B1(G71gat), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n676), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  INV_X1    g551(.A(new_n698), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n488), .A2(new_n528), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n753), .A2(new_n687), .B1(new_n754), .B2(new_n688), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n576), .A2(new_n265), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n652), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT111), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n481), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n698), .A2(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n698), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n481), .A2(G85gat), .A3(new_n681), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT112), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n760), .A2(new_n768), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n759), .B2(new_n428), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n681), .B1(new_n763), .B2(new_n764), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(new_n591), .A3(new_n503), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n759), .B2(new_n669), .ZN(new_n778));
  INV_X1    g577(.A(G99gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n771), .A2(new_n779), .A3(new_n484), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT113), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n485), .A2(G106gat), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT53), .B1(new_n771), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT114), .B(G106gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n759), .B2(new_n485), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n755), .A2(new_n676), .A3(new_n758), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n791), .A2(new_n788), .B1(new_n771), .B2(new_n786), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(G1339gat));
  NAND4_X1  g593(.A1(new_n576), .A2(new_n266), .A3(new_n619), .A4(new_n681), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n636), .A2(new_n622), .A3(new_n637), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT54), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n639), .A2(new_n641), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n647), .B1(new_n638), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n796), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n246), .B1(new_n240), .B2(new_n244), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n261), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n248), .A2(new_n254), .A3(new_n255), .A4(new_n262), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n616), .B2(new_n617), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n636), .A2(new_n637), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n621), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n640), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n797), .A2(KEYINPUT54), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n638), .A2(KEYINPUT101), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n650), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n810), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n808), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n652), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n265), .A3(new_n650), .ZN(new_n822));
  INV_X1    g621(.A(new_n803), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n819), .B1(new_n824), .B2(new_n619), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n795), .B1(new_n825), .B2(new_n695), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n677), .ZN(new_n827));
  INV_X1    g626(.A(new_n481), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n428), .A4(new_n484), .ZN(new_n829));
  OAI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n266), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n826), .A2(new_n828), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(new_n428), .A3(new_n404), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n266), .A2(G113gat), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT116), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n830), .B1(new_n837), .B2(new_n839), .ZN(G1340gat));
  INV_X1    g639(.A(G120gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n652), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n834), .B2(new_n836), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n681), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n841), .ZN(new_n846));
  OR3_X1    g645(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n843), .B2(new_n846), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1341gat));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n357), .A3(new_n576), .ZN(new_n850));
  INV_X1    g649(.A(new_n695), .ZN(new_n851));
  OAI21_X1  g650(.A(G127gat), .B1(new_n829), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1342gat));
  NOR2_X1   g652(.A1(new_n503), .A2(new_n619), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n831), .A2(new_n360), .A3(new_n404), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT118), .Z(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n829), .B2(new_n619), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n857), .B(new_n858), .C1(KEYINPUT56), .C2(new_n855), .ZN(G1343gat));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n831), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n669), .A2(new_n329), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n831), .B2(new_n860), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n266), .A2(G141gat), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n861), .A2(new_n863), .A3(new_n428), .A4(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n670), .A2(new_n481), .A3(new_n503), .ZN(new_n866));
  INV_X1    g665(.A(new_n795), .ZN(new_n867));
  INV_X1    g666(.A(new_n819), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n817), .A2(new_n265), .A3(new_n650), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT119), .B1(new_n799), .B2(new_n802), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n816), .A2(new_n871), .A3(new_n801), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n796), .A3(new_n872), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n869), .A2(new_n873), .B1(new_n652), .B2(new_n820), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n868), .B1(new_n874), .B2(new_n618), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n867), .B1(new_n875), .B2(new_n575), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n677), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n826), .A2(new_n329), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n866), .B(new_n877), .C1(KEYINPUT57), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n266), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n865), .B1(new_n880), .B2(new_n278), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT58), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n681), .A2(G148gat), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n861), .A2(new_n863), .A3(new_n428), .A4(new_n883), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT121), .Z(new_n885));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n873), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n618), .B1(new_n886), .B2(new_n821), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n887), .B2(new_n819), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(new_n868), .C1(new_n874), .C2(new_n618), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n575), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n795), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n677), .A2(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n866), .A2(new_n652), .ZN(new_n897));
  OAI21_X1  g696(.A(G148gat), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT59), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n280), .A2(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n879), .B2(new_n681), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n885), .B1(new_n903), .B2(new_n904), .ZN(G1345gat));
  NAND2_X1  g704(.A1(new_n861), .A2(new_n863), .ZN(new_n906));
  OR4_X1    g705(.A1(G155gat), .A2(new_n906), .A3(new_n503), .A4(new_n575), .ZN(new_n907));
  OAI21_X1  g706(.A(G155gat), .B1(new_n879), .B2(new_n851), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n879), .B2(new_n619), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n854), .A2(new_n283), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n906), .B2(new_n911), .ZN(G1347gat));
  AND2_X1   g711(.A1(new_n826), .A2(new_n481), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(new_n503), .A3(new_n404), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n336), .A3(new_n265), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n827), .A2(new_n481), .A3(new_n503), .A4(new_n484), .ZN(new_n916));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n266), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1348gat));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n333), .A3(new_n652), .ZN(new_n919));
  OAI21_X1  g718(.A(G176gat), .B1(new_n916), .B2(new_n681), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1349gat));
  NAND3_X1  g720(.A1(new_n914), .A2(new_n366), .A3(new_n576), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n347), .B1(new_n916), .B2(new_n851), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g724(.A1(new_n914), .A2(new_n339), .A3(new_n618), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT124), .Z(new_n927));
  OAI21_X1  g726(.A(G190gat), .B1(new_n916), .B2(new_n619), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1351gat));
  AND4_X1   g729(.A1(new_n481), .A2(new_n666), .A3(new_n503), .A4(new_n668), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n576), .B1(new_n875), .B2(KEYINPUT123), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n867), .B1(new_n932), .B2(new_n890), .ZN(new_n933));
  INV_X1    g732(.A(new_n893), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n895), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(G197gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(new_n266), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n913), .A2(new_n503), .A3(new_n329), .A4(new_n669), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n938), .A2(KEYINPUT125), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(KEYINPUT125), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n265), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n937), .B1(new_n942), .B2(new_n936), .ZN(G1352gat));
  NOR3_X1   g742(.A1(new_n938), .A2(G204gat), .A3(new_n681), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT62), .ZN(new_n945));
  OAI21_X1  g744(.A(G204gat), .B1(new_n935), .B2(new_n681), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1353gat));
  NAND4_X1  g746(.A1(new_n939), .A2(new_n271), .A3(new_n576), .A4(new_n940), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n271), .B1(KEYINPUT126), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n950), .B(new_n951), .C1(new_n935), .C2(new_n575), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n894), .A2(new_n576), .A3(new_n895), .A4(new_n931), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n954), .B2(new_n950), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n948), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g757(.A(KEYINPUT127), .B(new_n948), .C1(new_n953), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1354gat));
  NAND3_X1  g759(.A1(new_n941), .A2(new_n272), .A3(new_n618), .ZN(new_n961));
  OAI21_X1  g760(.A(G218gat), .B1(new_n935), .B2(new_n619), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1355gat));
endmodule


