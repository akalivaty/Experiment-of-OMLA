//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  XNOR2_X1  g000(.A(KEYINPUT78), .B(G125), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G140), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(KEYINPUT77), .A3(G125), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n188), .A2(KEYINPUT16), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  AOI21_X1  g009(.A(G146), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(G237), .A2(G953), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(G143), .A3(G214), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(G143), .B1(new_n200), .B2(G214), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT17), .B(G131), .C1(new_n202), .C2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n202), .A2(new_n203), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n202), .B2(new_n203), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n204), .B1(new_n209), .B2(KEYINPUT17), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n199), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT88), .B1(new_n202), .B2(new_n203), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n200), .A2(G214), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT88), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(new_n201), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT89), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT18), .A2(G131), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n192), .A2(new_n193), .ZN(new_n224));
  INV_X1    g038(.A(G125), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT78), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G125), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n226), .A2(new_n228), .A3(G140), .ZN(new_n229));
  OAI21_X1  g043(.A(G146), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(G140), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n190), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n230), .A2(new_n233), .B1(new_n221), .B2(new_n205), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n220), .B1(new_n219), .B2(new_n222), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n212), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n219), .A2(new_n222), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT89), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(KEYINPUT90), .A3(new_n223), .A4(new_n234), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n211), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G113), .B(G122), .ZN(new_n243));
  INV_X1    g057(.A(G104), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n242), .A2(KEYINPUT94), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(new_n245), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT94), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n241), .B2(new_n245), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n247), .B(new_n248), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G475), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT92), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n237), .A2(new_n240), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT19), .B1(new_n224), .B2(new_n229), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT19), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n190), .A2(new_n231), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n232), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n198), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n261), .A2(KEYINPUT91), .B1(new_n208), .B2(new_n207), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT91), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n198), .A3(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n255), .B(new_n246), .C1(new_n256), .C2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n237), .A2(new_n240), .B1(new_n262), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT92), .B1(new_n267), .B2(new_n245), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n268), .A3(new_n249), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n270));
  NOR2_X1   g084(.A1(G475), .A2(G902), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n271), .B(KEYINPUT93), .Z(new_n272));
  AND3_X1   g086(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n270), .B1(new_n269), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n254), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT98), .ZN(new_n276));
  XNOR2_X1  g090(.A(G128), .B(G143), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n215), .A2(G128), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n279), .B(G134), .C1(new_n280), .C2(new_n278), .ZN(new_n281));
  XNOR2_X1  g095(.A(G116), .B(G122), .ZN(new_n282));
  INV_X1    g096(.A(G107), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT14), .A3(G122), .ZN(new_n289));
  INV_X1    g103(.A(new_n282), .ZN(new_n290));
  OAI211_X1 g104(.A(G107), .B(new_n289), .C1(new_n290), .C2(KEYINPUT14), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n277), .A2(new_n285), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n292), .A2(new_n286), .B1(new_n283), .B2(new_n282), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n287), .A2(KEYINPUT96), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT82), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT75), .B(G217), .ZN(new_n297));
  INV_X1    g111(.A(G953), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT97), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n296), .A2(KEYINPUT97), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT96), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n281), .A2(new_n284), .A3(new_n305), .A4(new_n286), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n294), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n304), .B1(new_n294), .B2(new_n306), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n276), .B(new_n248), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  OR2_X1    g124(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n309), .B(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n275), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(G234), .A2(G237), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n315), .A2(G902), .A3(G953), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT21), .B(G898), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT99), .A2(G952), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT99), .A2(G952), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n298), .B(new_n315), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT100), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G210), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT65), .B1(new_n232), .B2(G143), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n215), .A3(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n232), .A2(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT64), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n215), .A2(KEYINPUT64), .A3(G146), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT0), .ZN(new_n335));
  INV_X1    g149(.A(G128), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n331), .A2(new_n333), .A3(new_n334), .A4(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n337), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n215), .A2(G146), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n332), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n336), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n187), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n336), .A2(KEYINPUT1), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n331), .A2(new_n333), .A3(new_n334), .A4(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n215), .A2(G146), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n352));
  OAI21_X1  g166(.A(G128), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n341), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n354), .A3(new_n187), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n344), .A2(KEYINPUT87), .A3(new_n345), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n348), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G224), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n359), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n348), .A2(new_n361), .A3(new_n355), .A4(new_n356), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(new_n244), .B2(G107), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n283), .A3(G104), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n244), .A2(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G101), .ZN(new_n370));
  INV_X1    g184(.A(G101), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n365), .A2(new_n367), .A3(new_n371), .A4(new_n368), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(KEYINPUT4), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(new_n374), .A3(G101), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT2), .B(G113), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G116), .B(G119), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(G116), .B(G119), .Z(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n376), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT68), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT68), .B1(new_n379), .B2(new_n381), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n373), .B(new_n375), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n378), .A2(KEYINPUT5), .ZN(new_n385));
  OR3_X1    g199(.A1(new_n288), .A2(KEYINPUT5), .A3(G119), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(G113), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT85), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n244), .A2(G107), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n283), .A2(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(G101), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n372), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n385), .A2(new_n394), .A3(G113), .A4(new_n386), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n388), .A2(new_n393), .A3(new_n395), .A4(new_n379), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n384), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n384), .A2(KEYINPUT86), .A3(new_n396), .ZN(new_n400));
  XNOR2_X1  g214(.A(G110), .B(G122), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n384), .A2(new_n396), .A3(new_n401), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT6), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n401), .B1(new_n397), .B2(new_n398), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n364), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n401), .B(KEYINPUT8), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n387), .A2(new_n379), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(new_n393), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n388), .A2(new_n379), .A3(new_n395), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n393), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n346), .A2(new_n355), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n361), .A2(KEYINPUT7), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n404), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n357), .A2(new_n416), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n327), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n407), .A2(new_n400), .B1(KEYINPUT6), .B2(new_n404), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n363), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n326), .A3(new_n420), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G221), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n296), .B2(new_n248), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G140), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n298), .A2(G227), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n434), .B(new_n435), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n350), .A2(new_n354), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT70), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n350), .A2(KEYINPUT70), .A3(new_n354), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n372), .A2(new_n391), .A3(KEYINPUT10), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n373), .A2(new_n338), .A3(new_n343), .A4(new_n375), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n353), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n392), .B1(new_n446), .B2(new_n350), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n444), .B1(new_n447), .B2(KEYINPUT10), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT11), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(KEYINPUT66), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n285), .A2(G137), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(KEYINPUT66), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n455));
  INV_X1    g269(.A(G137), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT11), .A4(G134), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n285), .A2(G137), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n454), .A2(new_n459), .A3(G131), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n456), .A2(G134), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n451), .B2(new_n452), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n455), .A2(KEYINPUT11), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n455), .A2(KEYINPUT11), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n456), .A2(G134), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n206), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n436), .B1(new_n449), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n467), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n462), .A2(new_n206), .A3(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n443), .B2(new_n448), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n437), .A2(new_n393), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n472), .B1(new_n447), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT12), .B1(new_n472), .B2(KEYINPUT84), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI221_X1 g292(.A(new_n472), .B1(KEYINPUT84), .B2(KEYINPUT12), .C1(new_n447), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n447), .A2(KEYINPUT10), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n481), .A2(new_n468), .A3(new_n442), .A4(new_n444), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n436), .B(KEYINPUT83), .Z(new_n484));
  OAI21_X1  g298(.A(new_n474), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n433), .B1(new_n485), .B2(new_n248), .ZN(new_n486));
  INV_X1    g300(.A(new_n436), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n480), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n473), .B2(new_n482), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n433), .B(new_n248), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n432), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n429), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n325), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n452), .B2(new_n461), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n471), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n471), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n497), .A2(new_n439), .A3(new_n440), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n382), .A2(new_n383), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n338), .B(new_n343), .C1(new_n460), .C2(new_n467), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n505), .B(KEYINPUT73), .Z(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n502), .ZN(new_n507));
  INV_X1    g321(.A(new_n501), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n503), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT72), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(KEYINPUT28), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n200), .A2(G210), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT27), .Z(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT29), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n506), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n503), .A2(new_n504), .ZN(new_n522));
  INV_X1    g336(.A(new_n517), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n437), .A2(new_n471), .A3(new_n495), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n502), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n508), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n522), .A2(new_n523), .A3(new_n505), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n518), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n500), .A2(KEYINPUT30), .A3(new_n502), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  AOI211_X1 g346(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n502), .C2(new_n524), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n508), .B(new_n529), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n523), .B1(new_n534), .B2(new_n503), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n248), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G472), .B1(new_n521), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n505), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n526), .B1(new_n503), .B2(new_n504), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n517), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n503), .A2(new_n523), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n534), .A2(KEYINPUT31), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT31), .B1(new_n534), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT71), .B(new_n542), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n539), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n537), .B1(new_n550), .B2(KEYINPUT32), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n549), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n539), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT74), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n556));
  INV_X1    g370(.A(new_n554), .ZN(new_n557));
  AOI211_X1 g371(.A(new_n556), .B(new_n557), .C1(new_n548), .C2(new_n549), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n551), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G234), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n297), .B1(new_n560), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G119), .B(G128), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT76), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT24), .B(G110), .Z(new_n565));
  INV_X1    g379(.A(G119), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G128), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n336), .A2(KEYINPUT23), .A3(G119), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(G128), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(KEYINPUT23), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n564), .A2(new_n565), .B1(G110), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n196), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT79), .B(new_n571), .C1(new_n572), .C2(new_n196), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT80), .B(G110), .ZN(new_n578));
  OAI22_X1  g392(.A1(new_n564), .A2(new_n565), .B1(new_n570), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n198), .A3(new_n233), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT22), .B(G137), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n430), .A2(new_n560), .A3(G953), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n580), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n248), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n562), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n562), .A2(G902), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n586), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT81), .B1(new_n559), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n534), .A2(new_n543), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT31), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n534), .A2(KEYINPUT31), .A3(new_n543), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT71), .B1(new_n601), .B2(new_n542), .ZN(new_n602));
  INV_X1    g416(.A(new_n549), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n538), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n553), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n554), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n556), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n552), .A2(KEYINPUT74), .A3(new_n554), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n605), .A2(new_n607), .A3(new_n537), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT81), .ZN(new_n610));
  INV_X1    g424(.A(new_n595), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n494), .B1(new_n596), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n371), .ZN(G3));
  NOR2_X1   g428(.A1(new_n307), .A2(new_n308), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n304), .B2(KEYINPUT101), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n310), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n310), .B(new_n248), .C1(new_n307), .C2(new_n308), .ZN(new_n619));
  NAND2_X1  g433(.A1(G478), .A2(G902), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n275), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n427), .A2(new_n428), .A3(new_n323), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n492), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n248), .B1(new_n602), .B2(new_n603), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n550), .B1(new_n627), .B2(G472), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n625), .A2(new_n611), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  INV_X1    g445(.A(new_n624), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n628), .A2(new_n611), .A3(new_n626), .A4(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n254), .B(new_n313), .C1(new_n273), .C2(new_n274), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  XNOR2_X1  g451(.A(new_n588), .B(new_n589), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n581), .B(new_n639), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n638), .A2(new_n562), .B1(new_n593), .B2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n641), .A2(new_n429), .A3(new_n492), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n325), .A2(new_n628), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT37), .B(G110), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  XNOR2_X1  g459(.A(new_n321), .B(KEYINPUT102), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n316), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n634), .A2(new_n649), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n609), .A2(new_n642), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n336), .ZN(G30));
  INV_X1    g466(.A(new_n428), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n649), .B(KEYINPUT39), .Z(new_n654));
  NAND2_X1  g468(.A1(new_n626), .A2(new_n654), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n653), .B(new_n312), .C1(new_n655), .C2(KEYINPUT40), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n427), .B(KEYINPUT38), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(G472), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n534), .A2(new_n503), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n523), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n523), .B1(new_n510), .B2(new_n512), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n663), .A2(G902), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n605), .B1(new_n660), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n607), .A2(new_n608), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n659), .A2(new_n275), .A3(new_n641), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  NOR2_X1   g484(.A1(new_n623), .A2(new_n649), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n671), .B(new_n642), .C1(new_n667), .C2(new_n551), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT103), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n609), .A2(new_n674), .A3(new_n642), .A4(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT104), .B(G146), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G48));
  OAI21_X1  g492(.A(new_n248), .B1(new_n488), .B2(new_n489), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n432), .A3(new_n490), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n680), .A2(new_n490), .A3(KEYINPUT105), .A4(new_n432), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n609), .A2(new_n611), .A3(new_n625), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NOR2_X1   g502(.A1(new_n634), .A2(new_n624), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n609), .A2(new_n611), .A3(new_n685), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  INV_X1    g505(.A(new_n314), .ZN(new_n692));
  INV_X1    g506(.A(new_n681), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n428), .A3(new_n427), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n641), .A3(new_n324), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n609), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n627), .A2(new_n698), .A3(G472), .ZN(new_n699));
  AOI21_X1  g513(.A(G902), .B1(new_n548), .B2(new_n549), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT106), .B1(new_n700), .B2(new_n660), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n653), .B(new_n312), .C1(new_n422), .C2(new_n426), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n275), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n683), .A2(new_n323), .A3(new_n684), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n506), .A2(new_n513), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n517), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n539), .B1(new_n708), .B2(new_n601), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n702), .A2(new_n706), .A3(new_n611), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  AOI21_X1  g526(.A(new_n709), .B1(new_n699), .B2(new_n701), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n640), .A2(new_n593), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n592), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n694), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n671), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n492), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(KEYINPUT107), .B(new_n432), .C1(new_n486), .C2(new_n491), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n427), .A2(new_n653), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n609), .A2(new_n611), .A3(new_n671), .A4(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n551), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n595), .B1(new_n728), .B2(new_n606), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(KEYINPUT42), .A3(new_n671), .A4(new_n724), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(G131), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G33));
  NAND4_X1  g547(.A1(new_n609), .A2(new_n611), .A3(new_n650), .A4(new_n724), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  OAI211_X1 g549(.A(new_n622), .B(new_n254), .C1(new_n274), .C2(new_n273), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n736), .B1(KEYINPUT109), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n738), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n628), .A2(new_n641), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n433), .B1(new_n485), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n745), .B2(new_n485), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT46), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n491), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n748), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n431), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n654), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n723), .B(KEYINPUT110), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n743), .A2(new_n744), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n456), .ZN(G39));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n752), .B(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n559), .A2(new_n595), .A3(new_n671), .A4(new_n723), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G140), .ZN(G42));
  NAND2_X1  g576(.A1(new_n680), .A2(new_n490), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT49), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(KEYINPUT49), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n431), .A2(new_n653), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n611), .A2(new_n764), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n668), .A2(new_n658), .A3(new_n736), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT111), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n651), .B1(new_n673), .B2(new_n675), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n704), .A2(new_n492), .A3(new_n649), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n668), .A2(new_n772), .A3(new_n641), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n718), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n686), .A2(new_n690), .A3(new_n711), .A4(new_n696), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n713), .A2(new_n715), .A3(new_n671), .A4(new_n724), .ZN(new_n777));
  INV_X1    g591(.A(new_n649), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n626), .A2(new_n715), .A3(new_n778), .A4(new_n723), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n609), .A2(new_n692), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n777), .A2(new_n734), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n776), .A2(new_n781), .A3(new_n731), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n775), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n771), .A2(new_n785), .A3(new_n718), .A4(new_n773), .ZN(new_n786));
  INV_X1    g600(.A(new_n494), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n275), .A2(new_n622), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT112), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(new_n633), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n792), .A2(new_n633), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT113), .B1(new_n613), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n643), .A2(new_n635), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n786), .A2(new_n795), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n770), .B1(new_n784), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n782), .B1(KEYINPUT52), .B2(new_n774), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n797), .A2(new_n795), .A3(new_n798), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(KEYINPUT53), .A4(new_n786), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT114), .B1(new_n804), .B2(KEYINPUT54), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n800), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n800), .A2(new_n803), .A3(new_n809), .A4(new_n806), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n805), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n804), .A2(KEYINPUT54), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n808), .A2(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n646), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n740), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n817), .A2(new_n611), .A3(new_n713), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n658), .A2(new_n428), .A3(new_n681), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n680), .A2(new_n431), .A3(new_n490), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n754), .B1(new_n759), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n818), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n817), .A2(new_n693), .A3(new_n723), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n723), .A2(new_n693), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n668), .A2(new_n595), .A3(new_n321), .A4(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n275), .A2(new_n622), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n826), .A2(new_n716), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n822), .A2(new_n825), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT117), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n826), .A2(new_n729), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT48), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n818), .A2(new_n717), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n298), .B1(new_n319), .B2(new_n320), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n828), .B2(new_n791), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n833), .B2(new_n832), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n815), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(G952), .A2(G953), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n769), .B1(new_n844), .B2(new_n845), .ZN(G75));
  NOR2_X1   g660(.A1(new_n298), .A2(G952), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n248), .B1(new_n800), .B2(new_n803), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n849), .B2(G210), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n363), .B(KEYINPUT55), .Z(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT119), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n423), .A2(new_n424), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT118), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n852), .B(new_n854), .Z(new_n855));
  OAI21_X1  g669(.A(new_n848), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n850), .B2(new_n855), .ZN(G51));
  NAND2_X1  g671(.A1(new_n807), .A2(KEYINPUT120), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n800), .A2(new_n803), .A3(new_n859), .A4(new_n806), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n812), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n804), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n748), .B(KEYINPUT57), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n489), .B2(new_n488), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n849), .B(new_n746), .C1(new_n745), .C2(new_n485), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n847), .B1(new_n868), .B2(new_n869), .ZN(G54));
  NAND3_X1  g684(.A1(new_n849), .A2(KEYINPUT58), .A3(G475), .ZN(new_n871));
  INV_X1    g685(.A(new_n269), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(new_n847), .ZN(G60));
  XOR2_X1   g689(.A(new_n620), .B(KEYINPUT59), .Z(new_n876));
  NOR3_X1   g690(.A1(new_n811), .A2(new_n814), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n848), .B1(new_n877), .B2(new_n617), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n879));
  INV_X1    g693(.A(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n617), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n804), .B2(KEYINPUT54), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n862), .B(new_n806), .C1(new_n800), .C2(new_n803), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n879), .B(new_n881), .C1(new_n884), .C2(new_n861), .ZN(new_n885));
  INV_X1    g699(.A(new_n881), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT122), .B1(new_n865), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n878), .A2(new_n888), .ZN(G63));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n890));
  NAND2_X1  g704(.A1(G217), .A2(G902), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT60), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n804), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n586), .A2(new_n587), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(KEYINPUT123), .A3(new_n894), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n804), .A2(new_n640), .A3(new_n892), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n900), .A2(KEYINPUT61), .A3(new_n848), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n890), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n890), .A2(new_n901), .A3(new_n897), .A4(new_n898), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n895), .A2(new_n848), .A3(new_n900), .ZN(new_n904));
  OAI22_X1  g718(.A1(new_n902), .A2(new_n903), .B1(KEYINPUT61), .B2(new_n904), .ZN(G66));
  INV_X1    g719(.A(new_n317), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n298), .B1(new_n906), .B2(G224), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n802), .A2(new_n776), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(new_n298), .ZN(new_n909));
  INV_X1    g723(.A(G898), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n854), .B1(new_n910), .B2(G953), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n909), .B(new_n911), .ZN(G69));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n753), .A2(new_n704), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n729), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n761), .A2(new_n734), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n731), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n756), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n718), .A3(new_n771), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n257), .A2(new_n259), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n647), .B2(new_n298), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n669), .A2(new_n718), .A3(new_n771), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n792), .A2(new_n634), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n655), .A2(new_n653), .A3(new_n427), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n927), .B(new_n928), .C1(new_n789), .C2(new_n788), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n761), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n926), .A2(new_n756), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(KEYINPUT62), .B2(new_n925), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n932), .A2(new_n298), .ZN(new_n933));
  OAI221_X1 g747(.A(new_n913), .B1(new_n920), .B2(new_n924), .C1(new_n933), .C2(new_n923), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n298), .B1(G227), .B2(G900), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G72));
  NAND2_X1  g750(.A1(G472), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT63), .Z(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n919), .B2(new_n908), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n941), .B(new_n938), .C1(new_n919), .C2(new_n908), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n523), .B(new_n661), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n932), .B2(new_n908), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n847), .B1(new_n944), .B2(new_n663), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n534), .A2(new_n543), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n804), .B(new_n938), .C1(new_n946), .C2(new_n535), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT127), .B1(new_n943), .B2(new_n948), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G57));
endmodule


