//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT15), .B1(new_n202), .B2(G43gat), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n203), .B1(G43gat), .B2(new_n202), .ZN(new_n204));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT96), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n204), .B1(KEYINPUT100), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(KEYINPUT99), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n207), .A2(KEYINPUT100), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(KEYINPUT99), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n208), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT97), .B(G43gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n202), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT98), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n202), .A2(G43gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(new_n220), .B2(KEYINPUT98), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT15), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n204), .B1(new_n207), .B2(new_n214), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT101), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n232), .B(new_n233), .C1(G1gat), .C2(new_n230), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n234), .B(G8gat), .Z(new_n235));
  NAND3_X1  g034(.A1(new_n225), .A2(KEYINPUT17), .A3(new_n226), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n235), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n227), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n238), .A4(new_n240), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n227), .B(new_n239), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n238), .B(KEYINPUT13), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT94), .B(KEYINPUT11), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G169gat), .B(G197gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT12), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n248), .A2(KEYINPUT95), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n248), .B2(KEYINPUT95), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G169gat), .ZN(new_n260));
  INV_X1    g059(.A(G176gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT23), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(G169gat), .B2(G176gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT25), .A4(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G190gat), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT24), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n274), .A2(KEYINPUT65), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT65), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n266), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(new_n272), .A3(KEYINPUT64), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n274), .A2(new_n275), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT64), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n282), .A2(new_n283), .A3(new_n285), .A4(new_n267), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT25), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n279), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  AND4_X1   g089(.A1(new_n282), .A2(new_n283), .A3(new_n285), .A4(new_n267), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n281), .ZN(new_n295));
  NAND2_X1  g094(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n272), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT65), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n274), .A2(KEYINPUT65), .A3(new_n275), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n267), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n266), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT67), .B1(new_n293), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n289), .A2(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G127gat), .B(G134gat), .Z(new_n306));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(KEYINPUT1), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(G113gat), .B(G120gat), .Z(new_n309));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G134gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT26), .B1(new_n260), .B2(new_n261), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n314), .A2(new_n265), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT26), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n274), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(G183gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(G190gat), .B1(new_n319), .B2(G183gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n295), .A2(KEYINPUT27), .A3(new_n296), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT28), .B1(new_n325), .B2(new_n323), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g127(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n325), .C2(new_n323), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n318), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n305), .A2(KEYINPUT69), .A3(new_n313), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n308), .A2(new_n312), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n288), .B1(new_n279), .B2(new_n287), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n293), .A2(new_n303), .A3(KEYINPUT67), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n318), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n323), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n321), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n338), .A2(KEYINPUT68), .B1(new_n323), .B2(new_n322), .ZN(new_n339));
  INV_X1    g138(.A(new_n329), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n332), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n330), .A2(new_n333), .A3(new_n313), .A4(new_n334), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n331), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G227gat), .A2(G233gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT34), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(KEYINPUT74), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n348), .B(new_n349), .C1(new_n346), .C2(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n350), .A2(KEYINPUT73), .ZN(new_n353));
  INV_X1    g152(.A(new_n349), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT73), .B(new_n350), .C1(new_n346), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n346), .B2(new_n354), .ZN(new_n359));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT72), .ZN(new_n361));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n359), .A2(KEYINPUT71), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n354), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n366), .A2(KEYINPUT32), .A3(new_n358), .A4(new_n363), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n366), .B2(new_n357), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n369), .A2(KEYINPUT71), .B1(KEYINPUT32), .B2(new_n366), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n356), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n373), .B(new_n356), .C1(new_n368), .C2(new_n370), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n366), .A2(KEYINPUT32), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n359), .A2(new_n378), .A3(new_n364), .ZN(new_n379));
  OAI22_X1  g178(.A1(new_n377), .A2(new_n379), .B1(new_n365), .B2(new_n367), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n376), .B1(new_n380), .B2(new_n356), .ZN(new_n381));
  INV_X1    g180(.A(new_n370), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n369), .A2(new_n378), .ZN(new_n383));
  INV_X1    g182(.A(new_n367), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(KEYINPUT75), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n375), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT36), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT92), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT82), .ZN(new_n393));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  XOR2_X1   g194(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n335), .B2(new_n341), .ZN(new_n398));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n330), .A2(new_n333), .A3(KEYINPUT80), .A4(new_n334), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G197gat), .B(G204gat), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT22), .ZN(new_n404));
  INV_X1    g203(.A(G211gat), .ZN(new_n405));
  INV_X1    g204(.A(G218gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT78), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n410), .B(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(KEYINPUT77), .A3(new_n408), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n293), .A2(new_n303), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n330), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT81), .B(new_n399), .C1(new_n421), .C2(KEYINPUT29), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT29), .B1(new_n330), .B2(new_n420), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(new_n400), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n402), .A2(new_n419), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n398), .A2(new_n427), .A3(new_n399), .A4(new_n401), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n417), .B(KEYINPUT79), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n400), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n395), .B(new_n396), .C1(new_n432), .C2(KEYINPUT37), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n402), .A2(new_n425), .A3(new_n422), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n429), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n428), .A2(new_n430), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n435), .A2(KEYINPUT90), .B1(new_n419), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n438), .A3(new_n429), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n433), .B1(new_n440), .B2(KEYINPUT37), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n432), .A2(new_n395), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n444));
  INV_X1    g243(.A(G155gat), .ZN(new_n445));
  INV_X1    g244(.A(G162gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(KEYINPUT84), .A3(new_n448), .ZN(new_n452));
  INV_X1    g251(.A(G141gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G148gat), .ZN(new_n454));
  INV_X1    g253(.A(G148gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G141gat), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n454), .A2(new_n456), .B1(KEYINPUT2), .B2(new_n448), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n451), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G141gat), .B(G148gat), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n448), .A2(KEYINPUT2), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n450), .B(new_n449), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n332), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n313), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n444), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(KEYINPUT4), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT4), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n313), .A2(new_n464), .A3(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n464), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n458), .A2(KEYINPUT3), .A3(new_n461), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n332), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n313), .A2(new_n464), .A3(KEYINPUT85), .A4(new_n472), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n467), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n469), .B1(new_n474), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G1gat), .B(G29gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT0), .ZN(new_n483));
  XNOR2_X1  g282(.A(G57gat), .B(G85gat), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT86), .A3(new_n473), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n313), .B1(new_n475), .B2(new_n464), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n468), .B1(new_n487), .B2(new_n477), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n489), .A3(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n486), .A2(new_n488), .A3(new_n444), .A4(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n481), .A2(KEYINPUT87), .A3(new_n485), .A4(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n481), .A2(new_n491), .ZN(new_n495));
  INV_X1    g294(.A(new_n485), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n485), .A3(new_n491), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT6), .B1(new_n501), .B2(new_n497), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n443), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n391), .B1(new_n441), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT37), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n426), .B2(new_n431), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(KEYINPUT93), .A3(new_n395), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n509));
  INV_X1    g308(.A(new_n395), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n508), .B(new_n511), .C1(KEYINPUT37), .C2(new_n432), .ZN(new_n512));
  INV_X1    g311(.A(new_n396), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n501), .A2(new_n497), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n493), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n497), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n442), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n505), .B1(new_n437), .B2(new_n439), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n518), .B(KEYINPUT92), .C1(new_n519), .C2(new_n433), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(G228gat), .A2(G233gat), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT29), .B1(new_n413), .B2(new_n416), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n462), .B1(new_n523), .B2(KEYINPUT3), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n476), .A2(new_n427), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n522), .B(new_n524), .C1(new_n419), .C2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G22gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n427), .B1(new_n411), .B2(new_n408), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n415), .A2(new_n409), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n475), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n429), .A2(new_n525), .B1(new_n462), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n527), .B(new_n528), .C1(new_n532), .C2(new_n522), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT88), .ZN(new_n534));
  XOR2_X1   g333(.A(G78gat), .B(G106gat), .Z(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G50gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n527), .B1(new_n532), .B2(new_n522), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G22gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n533), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n534), .A2(new_n540), .A3(new_n533), .A4(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n426), .A2(new_n431), .A3(KEYINPUT30), .A4(new_n510), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT83), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n432), .A2(new_n395), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n442), .B2(KEYINPUT30), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n486), .A2(new_n478), .A3(new_n490), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n468), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n551), .B(KEYINPUT39), .C1(new_n468), .C2(new_n466), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT39), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n553), .A3(new_n468), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n554), .A2(new_n555), .A3(new_n485), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n554), .B2(new_n485), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT40), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(KEYINPUT40), .B(new_n552), .C1(new_n556), .C2(new_n557), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n497), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n544), .B1(new_n549), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n521), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n516), .A2(new_n517), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n544), .B1(new_n549), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n368), .A2(new_n370), .A3(new_n356), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n374), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n373), .B1(new_n380), .B2(new_n356), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n568), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n390), .A2(new_n565), .A3(new_n567), .A4(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n544), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n546), .A2(new_n566), .A3(new_n548), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n375), .A2(new_n388), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n578));
  AOI211_X1 g377(.A(new_n569), .B(new_n544), .C1(new_n372), .C2(new_n374), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n549), .A2(KEYINPUT35), .A3(new_n566), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n259), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT107), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT7), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT107), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n589), .A2(new_n591), .A3(G85gat), .A4(G92gat), .ZN(new_n592));
  INV_X1    g391(.A(G85gat), .ZN(new_n593));
  INV_X1    g392(.A(G92gat), .ZN(new_n594));
  OAI211_X1 g393(.A(KEYINPUT107), .B(new_n590), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n593), .B2(new_n594), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT108), .ZN(new_n599));
  XOR2_X1   g398(.A(G99gat), .B(G106gat), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n599), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n229), .A2(new_n236), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n599), .B(new_n600), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n227), .A2(new_n606), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT109), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n605), .B1(new_n603), .B2(new_n607), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n587), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT110), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n613), .B1(new_n610), .B2(new_n611), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT110), .B1(new_n618), .B2(new_n587), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(KEYINPUT111), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n613), .A2(KEYINPUT111), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n612), .A2(new_n620), .A3(new_n587), .A4(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n617), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT105), .A2(G57gat), .ZN(new_n624));
  INV_X1    g423(.A(G64gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(KEYINPUT9), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT104), .B(G57gat), .Z(new_n632));
  OR2_X1    g431(.A1(new_n632), .A2(G64gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT9), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(G64gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n627), .B(KEYINPUT102), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n629), .B(KEYINPUT103), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n631), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT106), .B(KEYINPUT21), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G127gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n239), .B1(KEYINPUT21), .B2(new_n641), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G155gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n649), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n623), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n602), .A2(new_n642), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n606), .A2(new_n641), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n641), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n658), .A2(new_n659), .ZN(new_n666));
  INV_X1    g465(.A(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(G120gat), .B(G148gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT112), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n665), .A2(new_n668), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n657), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n583), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n566), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n549), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(G8gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT42), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(KEYINPUT42), .B2(new_n686), .ZN(G1325gat));
  INV_X1    g487(.A(new_n680), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n390), .A2(new_n573), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n569), .B1(new_n372), .B2(new_n374), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n583), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(G15gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n679), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n544), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  AOI21_X1  g499(.A(new_n623), .B1(new_n574), .B2(new_n582), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n656), .A2(new_n259), .A3(new_n678), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n209), .A3(new_n566), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n617), .A2(new_n619), .A3(new_n622), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n372), .A2(new_n374), .B1(new_n381), .B2(new_n387), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n567), .B(new_n573), .C1(new_n707), .C2(new_n568), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n546), .A2(new_n548), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n575), .B1(new_n709), .B2(new_n562), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n518), .B1(new_n519), .B2(new_n433), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n711), .A2(new_n391), .B1(new_n513), .B2(new_n512), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n712), .B2(new_n520), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  AOI22_X1  g513(.A1(KEYINPUT35), .A2(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n706), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n701), .A2(KEYINPUT44), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n702), .ZN(new_n721));
  INV_X1    g520(.A(new_n566), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n723), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n703), .A2(new_n210), .A3(new_n549), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT46), .Z(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n721), .B2(new_n709), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1329gat));
  OAI21_X1  g527(.A(new_n219), .B1(new_n721), .B2(new_n691), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n656), .A2(new_n219), .A3(new_n678), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n694), .A2(new_n706), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(KEYINPUT47), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1330gat));
  NAND4_X1  g535(.A1(new_n718), .A2(new_n719), .A3(new_n544), .A4(new_n702), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G50gat), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT48), .B1(new_n738), .B2(KEYINPUT113), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n703), .A2(new_n202), .A3(new_n544), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n739), .B(new_n741), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n574), .A2(new_n582), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n657), .A2(new_n258), .A3(new_n677), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n566), .B(KEYINPUT114), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g548(.A(new_n709), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT115), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1333gat));
  INV_X1    g553(.A(G71gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(new_n755), .A3(new_n693), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n745), .A2(new_n690), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(new_n755), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g558(.A1(new_n745), .A2(new_n544), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT116), .B(G78gat), .Z(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1335gat));
  NOR2_X1   g561(.A1(new_n656), .A2(new_n258), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n678), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n718), .A2(new_n719), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n722), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n769), .B(new_n706), .C1(new_n714), .C2(new_n715), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n763), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n743), .B2(new_n706), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n716), .A2(KEYINPUT117), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n774), .A2(new_n775), .A3(new_n763), .A4(new_n770), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n678), .A2(new_n593), .A3(new_n566), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n768), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  AOI21_X1  g578(.A(new_n594), .B1(new_n766), .B2(new_n549), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n549), .A2(new_n678), .A3(new_n594), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n781), .B(new_n782), .C1(new_n777), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT119), .B1(KEYINPUT120), .B2(KEYINPUT51), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n770), .A2(new_n763), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n774), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n774), .A2(new_n788), .A3(new_n763), .A4(new_n770), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT120), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n787), .B1(new_n790), .B2(new_n775), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n783), .B(KEYINPUT118), .Z(new_n792));
  AOI21_X1  g591(.A(new_n780), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n784), .B1(new_n793), .B2(new_n782), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n767), .B2(new_n691), .ZN(new_n795));
  INV_X1    g594(.A(G99gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n693), .A2(new_n796), .A3(new_n678), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n777), .B2(new_n797), .ZN(G1338gat));
  AOI21_X1  g597(.A(KEYINPUT51), .B1(new_n789), .B2(KEYINPUT120), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n575), .A2(G106gat), .A3(new_n677), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n799), .A2(new_n787), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n766), .B2(new_n544), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT53), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n773), .A2(new_n776), .A3(new_n800), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT121), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n773), .A2(new_n776), .A3(new_n808), .A4(new_n800), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n804), .A2(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n805), .A2(new_n812), .ZN(G1339gat));
  NOR3_X1   g612(.A1(new_n657), .A2(new_n258), .A3(new_n678), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n661), .A2(new_n662), .A3(new_n667), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n667), .B1(new_n661), .B2(new_n662), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n675), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n676), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT55), .B1(new_n816), .B2(new_n819), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n258), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n245), .A2(new_n246), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n238), .B1(new_n237), .B2(new_n240), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n253), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n248), .A2(new_n254), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n678), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n623), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n828), .A2(new_n832), .A3(new_n827), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n828), .A2(new_n827), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT122), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n706), .A2(new_n823), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n656), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n814), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR4_X1   g638(.A1(new_n839), .A2(new_n544), .A3(new_n389), .A4(new_n746), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n709), .ZN(new_n841));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n258), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n679), .A2(new_n259), .ZN(new_n843));
  INV_X1    g642(.A(new_n837), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n656), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n579), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n566), .A3(new_n709), .ZN(new_n847));
  INV_X1    g646(.A(G113gat), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n847), .A2(new_n848), .A3(new_n259), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n842), .A2(new_n849), .ZN(G1340gat));
  NOR2_X1   g649(.A1(new_n677), .A2(G120gat), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT123), .Z(new_n852));
  NAND2_X1  g651(.A1(new_n841), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n847), .B2(new_n677), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1341gat));
  INV_X1    g654(.A(G127gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n856), .A3(new_n656), .ZN(new_n857));
  OAI21_X1  g656(.A(G127gat), .B1(new_n847), .B2(new_n838), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n623), .A2(new_n549), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n847), .B2(new_n623), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n709), .A2(new_n566), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n690), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n834), .A2(new_n677), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n822), .A2(KEYINPUT124), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n822), .A2(KEYINPUT124), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n821), .A2(new_n256), .A3(new_n257), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n836), .B1(new_n875), .B2(new_n706), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n814), .B1(new_n876), .B2(new_n838), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n877), .A2(new_n878), .A3(new_n575), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n839), .B2(new_n575), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n869), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n453), .B1(new_n881), .B2(new_n258), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n690), .A2(new_n575), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n845), .A2(new_n747), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n549), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n258), .A2(new_n453), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT125), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT58), .B1(new_n882), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n259), .B(new_n869), .C1(new_n879), .C2(new_n880), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n888), .B(new_n891), .C1(new_n892), .C2(new_n453), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(G1344gat));
  NOR3_X1   g693(.A1(new_n884), .A2(new_n549), .A3(new_n677), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n455), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n880), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n869), .A2(new_n677), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n874), .B1(new_n872), .B2(new_n871), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n706), .B1(new_n902), .B2(new_n829), .ZN(new_n903));
  AND4_X1   g702(.A1(new_n706), .A2(new_n823), .A3(new_n833), .A4(new_n835), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n838), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n575), .B1(new_n905), .B2(new_n843), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n901), .B1(new_n906), .B2(KEYINPUT57), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT126), .B(new_n878), .C1(new_n877), .C2(new_n575), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n845), .A2(KEYINPUT57), .A3(new_n544), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n899), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n897), .B(new_n900), .C1(new_n911), .C2(new_n912), .ZN(G1345gat));
  INV_X1    g712(.A(new_n881), .ZN(new_n914));
  OAI21_X1  g713(.A(G155gat), .B1(new_n914), .B2(new_n838), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n885), .A2(new_n445), .A3(new_n656), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n914), .B2(new_n623), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n861), .A2(new_n446), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n884), .B2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n747), .A2(new_n709), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n846), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(new_n260), .A3(new_n259), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n709), .A2(new_n566), .ZN(new_n924));
  AND4_X1   g723(.A1(new_n575), .A2(new_n845), .A3(new_n707), .A4(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n258), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n923), .A2(new_n926), .ZN(G1348gat));
  OAI21_X1  g726(.A(G176gat), .B1(new_n922), .B2(new_n677), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n261), .A3(new_n678), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  OAI22_X1  g729(.A1(new_n922), .A2(new_n838), .B1(new_n270), .B2(new_n269), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n281), .A2(KEYINPUT27), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n838), .A2(new_n932), .A3(new_n320), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT60), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n925), .A2(new_n272), .A3(new_n706), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n846), .A2(new_n706), .A3(new_n921), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(G190gat), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n941), .B2(G190gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  NAND3_X1  g745(.A1(new_n845), .A2(new_n883), .A3(new_n924), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n947), .A2(G197gat), .A3(new_n259), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT127), .Z(new_n949));
  INV_X1    g748(.A(G197gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n691), .A2(new_n921), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n910), .A2(new_n258), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n949), .B1(new_n950), .B2(new_n953), .ZN(G1352gat));
  NOR3_X1   g753(.A1(new_n947), .A2(G204gat), .A3(new_n677), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n910), .A2(new_n678), .A3(new_n952), .ZN(new_n959));
  INV_X1    g758(.A(G204gat), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n957), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(G1353gat));
  OR3_X1    g760(.A1(new_n947), .A2(G211gat), .A3(new_n838), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n910), .A2(new_n656), .A3(new_n952), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  AND3_X1   g765(.A1(new_n910), .A2(new_n706), .A3(new_n952), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n706), .A2(new_n406), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n967), .A2(new_n406), .B1(new_n947), .B2(new_n968), .ZN(G1355gat));
endmodule


