//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G101), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT4), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(G101), .B1(new_n188), .B2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n189), .A2(new_n198), .A3(new_n192), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n189), .A2(new_n198), .A3(new_n192), .A4(KEYINPUT80), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n197), .B1(new_n204), .B2(new_n195), .ZN(new_n205));
  AND2_X1   g019(.A1(G116), .A2(G119), .ZN(new_n206));
  NOR2_X1   g020(.A1(G116), .A2(G119), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT2), .B(G113), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT68), .B1(new_n210), .B2(KEYINPUT67), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n209), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT2), .A2(G113), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT2), .A2(G113), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n214), .B(new_n215), .C1(new_n206), .C2(new_n207), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n213), .A3(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n218), .B1(new_n216), .B2(new_n217), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n212), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n191), .A2(G104), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n193), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n201), .B2(new_n202), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n229), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n207), .A2(new_n206), .B1(new_n230), .B2(new_n231), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n210), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n228), .A2(new_n237), .A3(KEYINPUT85), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT85), .B1(new_n228), .B2(new_n237), .ZN(new_n239));
  OAI22_X1  g053(.A1(new_n205), .A2(new_n224), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT86), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n240), .A2(KEYINPUT86), .A3(new_n242), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n187), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT87), .B1(new_n240), .B2(new_n242), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n220), .A2(new_n223), .ZN(new_n249));
  INV_X1    g063(.A(new_n195), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT4), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n196), .B1(new_n201), .B2(new_n202), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT87), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n256));
  INV_X1    g070(.A(new_n227), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n203), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n235), .A2(new_n236), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n216), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n256), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n228), .A2(new_n237), .A3(KEYINPUT85), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n254), .A2(new_n255), .A3(new_n241), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n248), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n243), .B2(KEYINPUT6), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n240), .A2(KEYINPUT88), .A3(new_n187), .A4(new_n242), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n247), .A2(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G146), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT64), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G146), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n273), .A3(G143), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n270), .A2(G143), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n270), .A2(G143), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n271), .A2(new_n273), .ZN(new_n281));
  INV_X1    g095(.A(G143), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n278), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G125), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT89), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n291));
  INV_X1    g105(.A(G128), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n274), .B2(KEYINPUT1), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n293), .B2(new_n283), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT64), .B(G146), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n279), .B1(new_n295), .B2(G143), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT1), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n295), .B2(G143), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT65), .B(new_n296), .C1(new_n298), .C2(new_n292), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n292), .A2(KEYINPUT1), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n274), .A2(new_n276), .A3(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n294), .A2(new_n299), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(KEYINPUT89), .A3(G125), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n290), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G953), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G224), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n305), .B(new_n307), .Z(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n288), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(KEYINPUT7), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n310), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n290), .A2(new_n303), .A3(new_n304), .A4(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT5), .B1(new_n206), .B2(new_n207), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n235), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n228), .B1(new_n315), .B2(new_n210), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n241), .B(KEYINPUT8), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n316), .B(new_n317), .C1(new_n228), .C2(new_n260), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n249), .A2(new_n253), .B1(new_n261), .B2(new_n262), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n255), .B1(new_n321), .B2(new_n241), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n240), .A2(KEYINPUT87), .A3(new_n242), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n325));
  INV_X1    g139(.A(G902), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n319), .B1(new_n248), .B2(new_n264), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT90), .B1(new_n328), .B2(G902), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n269), .A2(new_n308), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G210), .B1(G237), .B2(G902), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT91), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n331), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n329), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n267), .A2(new_n268), .ZN(new_n335));
  INV_X1    g149(.A(new_n246), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT86), .B1(new_n240), .B2(new_n242), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT6), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n265), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n308), .B(new_n335), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT91), .ZN(new_n342));
  INV_X1    g156(.A(new_n331), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n332), .A2(new_n333), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G125), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n300), .A2(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT16), .ZN(new_n349));
  OR3_X1    g163(.A1(new_n300), .A2(KEYINPUT16), .A3(G140), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(G146), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT73), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT73), .A4(G146), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n349), .A2(new_n350), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n353), .B(new_n354), .C1(G146), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(G237), .A2(G953), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n358), .A2(G143), .A3(G214), .ZN(new_n359));
  AOI21_X1  g173(.A(G143), .B1(new_n358), .B2(G214), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT17), .B(G131), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT93), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n357), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n361), .B(KEYINPUT92), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT93), .B1(new_n366), .B2(new_n356), .ZN(new_n367));
  INV_X1    g181(.A(new_n360), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n358), .A2(G143), .A3(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G131), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT17), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n365), .A2(new_n367), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(new_n188), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n370), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n380), .A2(new_n270), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n295), .A2(new_n380), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n375), .A2(new_n377), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n377), .B1(new_n375), .B2(new_n384), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n326), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G475), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT20), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n380), .B(KEYINPUT19), .Z(new_n391));
  OAI21_X1  g205(.A(new_n351), .B1(new_n391), .B2(new_n281), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n384), .B1(new_n372), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n377), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(G475), .A2(G902), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n390), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n397), .ZN(new_n399));
  AOI211_X1 g213(.A(KEYINPUT20), .B(new_n399), .C1(new_n385), .C2(new_n395), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n389), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G116), .B(G122), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G122), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(G116), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n191), .B1(new_n406), .B2(KEYINPUT14), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n404), .A2(new_n407), .B1(new_n191), .B2(new_n402), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n292), .A2(G143), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT96), .Z(new_n410));
  INV_X1    g224(.A(G134), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n282), .A2(G128), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT94), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n410), .B2(new_n413), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n408), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n409), .B(KEYINPUT96), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n413), .A2(new_n419), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n411), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n402), .B(new_n191), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n417), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT9), .B(G234), .ZN(new_n426));
  INV_X1    g240(.A(G217), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n426), .A2(new_n427), .A3(G953), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n417), .B(new_n428), .C1(new_n422), .C2(new_n424), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n326), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n433), .A2(new_n435), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(G234), .A2(G237), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n440), .A2(G952), .A3(new_n306), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n440), .A2(G902), .A3(G953), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(G898), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n401), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  OAI21_X1  g260(.A(G221), .B1(new_n426), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G469), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(new_n326), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT11), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n411), .B2(G137), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n411), .A2(G137), .ZN(new_n453));
  INV_X1    g267(.A(G137), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT11), .A3(G134), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G131), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n452), .A2(new_n455), .A3(new_n371), .A4(new_n453), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(KEYINPUT69), .A3(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n275), .B1(new_n295), .B2(G143), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n296), .A2(new_n285), .B1(new_n464), .B2(new_n277), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT10), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n292), .B1(new_n279), .B2(KEYINPUT1), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n302), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n203), .A3(new_n257), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n253), .A2(new_n465), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n294), .A2(new_n299), .A3(new_n302), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT81), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n466), .B(new_n227), .C1(new_n201), .C2(new_n202), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n471), .B2(new_n473), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n463), .B(new_n470), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT82), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n471), .B2(new_n228), .ZN(new_n478));
  INV_X1    g292(.A(new_n302), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n296), .B1(new_n298), .B2(new_n292), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n291), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n481), .A2(KEYINPUT82), .A3(new_n299), .A4(new_n258), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n469), .ZN(new_n484));
  INV_X1    g298(.A(new_n463), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT12), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n469), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n478), .B2(new_n482), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n489));
  INV_X1    g303(.A(new_n459), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n476), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n306), .A2(G227), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(G140), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT78), .B(G110), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT79), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n471), .A2(new_n473), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT81), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT83), .B1(new_n502), .B2(new_n470), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT83), .B(new_n470), .C1(new_n474), .C2(new_n475), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n485), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n496), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n476), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n492), .A2(new_n498), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n450), .B1(new_n510), .B2(G469), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n507), .B1(new_n506), .B2(new_n476), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n484), .A2(KEYINPUT12), .A3(new_n459), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n489), .B1(new_n488), .B2(new_n463), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n449), .B(new_n326), .C1(new_n512), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n448), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n345), .A2(new_n445), .A3(new_n446), .A4(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT32), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n358), .A2(G210), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT27), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT26), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n225), .ZN(new_n524));
  INV_X1    g338(.A(new_n453), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n411), .A2(G137), .ZN(new_n526));
  OAI21_X1  g340(.A(G131), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n458), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n471), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n461), .A2(new_n465), .A3(new_n462), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n224), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n528), .B1(new_n481), .B2(new_n299), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(KEYINPUT30), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT70), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n530), .A2(new_n537), .A3(KEYINPUT30), .A4(new_n531), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n224), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT66), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n490), .A2(new_n287), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n471), .B2(new_n529), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n542), .B2(KEYINPUT30), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  OAI211_X1 g358(.A(KEYINPUT66), .B(new_n544), .C1(new_n534), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n533), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT31), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI211_X1 g363(.A(KEYINPUT31), .B(new_n533), .C1(new_n539), .C2(new_n546), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n532), .A2(KEYINPUT71), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT71), .B1(new_n532), .B2(new_n551), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n532), .B1(new_n224), .B2(new_n542), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT28), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n524), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n549), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(G472), .A2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n519), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n532), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n539), .B2(new_n546), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n524), .A2(KEYINPUT29), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n530), .A2(new_n531), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n249), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n551), .B1(new_n567), .B2(new_n532), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n568), .A2(new_n552), .A3(new_n553), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT29), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n524), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n554), .A2(new_n556), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT29), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n565), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n539), .A2(new_n546), .ZN(new_n576));
  INV_X1    g390(.A(new_n533), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT31), .ZN(new_n579));
  INV_X1    g393(.A(new_n524), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n547), .A2(new_n548), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT32), .A3(new_n559), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n561), .A2(new_n575), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n427), .B1(G234), .B2(new_n326), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT23), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n233), .B2(G128), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n292), .A2(KEYINPUT23), .A3(G119), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n589), .B(new_n590), .C1(G119), .C2(new_n292), .ZN(new_n591));
  XNOR2_X1  g405(.A(G119), .B(G128), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT24), .B(G110), .Z(new_n593));
  OAI22_X1  g407(.A1(new_n591), .A2(G110), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n351), .A3(new_n382), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(G110), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT72), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT72), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n591), .A2(new_n598), .A3(G110), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n597), .A2(new_n599), .B1(new_n592), .B2(new_n593), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n600), .A2(new_n356), .A3(KEYINPUT74), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT74), .B1(new_n600), .B2(new_n356), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n356), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT74), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n600), .A2(KEYINPUT74), .A3(new_n356), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(KEYINPUT75), .A3(new_n595), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n306), .A2(G221), .A3(G234), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT22), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G137), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n595), .B(new_n614), .C1(new_n601), .C2(new_n602), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT76), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n610), .A2(KEYINPUT76), .A3(new_n595), .A4(new_n614), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n616), .A2(new_n621), .A3(new_n326), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT25), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(KEYINPUT77), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n587), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT77), .B(KEYINPUT25), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n616), .A2(new_n621), .A3(new_n326), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n616), .A2(new_n621), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n586), .A2(G902), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n625), .A2(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n585), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n518), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n225), .ZN(G3));
  AND3_X1   g448(.A1(new_n334), .A2(new_n331), .A3(new_n340), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n331), .B1(new_n334), .B2(new_n340), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n446), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT97), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n639), .B(new_n446), .C1(new_n635), .C2(new_n636), .ZN(new_n640));
  INV_X1    g454(.A(new_n444), .ZN(new_n641));
  INV_X1    g455(.A(new_n401), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n429), .A2(KEYINPUT99), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n425), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n425), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(KEYINPUT33), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n434), .A2(G902), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT98), .B1(new_n432), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  AOI211_X1 g464(.A(new_n650), .B(KEYINPUT33), .C1(new_n430), .C2(new_n431), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n646), .B(new_n647), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n433), .A2(new_n434), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n642), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n638), .A2(new_n640), .A3(new_n641), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n511), .A2(new_n516), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n447), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n583), .A2(new_n559), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n558), .A2(G902), .ZN(new_n661));
  INV_X1    g475(.A(G472), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n631), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n657), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT34), .B(G104), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NOR2_X1   g480(.A1(new_n401), .A2(new_n438), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n638), .A2(new_n640), .A3(new_n641), .A4(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n668), .A2(new_n659), .A3(new_n663), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT35), .B(G107), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  AND2_X1   g485(.A1(new_n345), .A2(new_n446), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n605), .A2(new_n611), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n615), .A2(KEYINPUT36), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n605), .B(new_n611), .C1(KEYINPUT36), .C2(new_n615), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n676), .A2(new_n630), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n625), .B2(new_n627), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(KEYINPUT100), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  AOI211_X1 g495(.A(new_n681), .B(new_n678), .C1(new_n625), .C2(new_n627), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n673), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n517), .A2(new_n445), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n672), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G12));
  NOR2_X1   g501(.A1(new_n680), .A2(new_n682), .ZN(new_n688));
  AND4_X1   g502(.A1(new_n517), .A2(new_n688), .A3(new_n638), .A4(new_n640), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n442), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n441), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n401), .A2(new_n438), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n585), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  AND2_X1   g512(.A1(new_n561), .A2(new_n584), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n524), .B1(new_n567), .B2(new_n532), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT101), .Z(new_n701));
  OAI21_X1  g515(.A(new_n326), .B1(new_n701), .B2(new_n547), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G472), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n642), .A2(new_n438), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n446), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n625), .A2(new_n627), .ZN(new_n708));
  INV_X1    g522(.A(new_n678), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n345), .B(KEYINPUT38), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT102), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT102), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n693), .B(KEYINPUT39), .Z(new_n716));
  NOR2_X1   g530(.A1(new_n659), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT40), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n714), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  NAND3_X1  g534(.A1(new_n401), .A2(new_n654), .A3(new_n693), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n699), .B2(new_n575), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n689), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  OAI21_X1  g538(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT83), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n463), .B1(new_n727), .B2(new_n504), .ZN(new_n728));
  INV_X1    g542(.A(new_n476), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n496), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n515), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n326), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G469), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n734), .A2(new_n447), .A3(new_n516), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n585), .A3(new_n631), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n657), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT41), .B(G113), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G15));
  NOR2_X1   g553(.A1(new_n668), .A2(new_n736), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(G116), .Z(G18));
  NAND3_X1  g555(.A1(new_n688), .A2(new_n585), .A3(new_n445), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n638), .A2(new_n640), .A3(new_n735), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT103), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n638), .A2(new_n640), .A3(new_n735), .A4(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n742), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n233), .ZN(G21));
  OAI211_X1 g562(.A(new_n579), .B(new_n582), .C1(new_n524), .C2(new_n569), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n559), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n631), .B(new_n750), .C1(new_n661), .C2(new_n662), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n734), .A2(new_n447), .A3(new_n516), .A4(new_n641), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n640), .A3(new_n638), .A4(new_n705), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  NAND2_X1  g569(.A1(new_n744), .A2(new_n746), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n710), .B(new_n750), .C1(new_n662), .C2(new_n661), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n721), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n401), .A2(new_n654), .A3(KEYINPUT104), .A4(new_n693), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n707), .B1(new_n330), .B2(new_n331), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n517), .A2(new_n332), .A3(new_n344), .A4(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n632), .A2(new_n767), .A3(new_n761), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n769), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n332), .A2(new_n766), .A3(new_n344), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n585), .A3(new_n631), .A4(new_n517), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT106), .B(new_n771), .C1(new_n773), .C2(new_n761), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n632), .B(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n761), .ZN(new_n778));
  INV_X1    g592(.A(new_n767), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(KEYINPUT42), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NAND4_X1  g596(.A1(new_n779), .A2(new_n585), .A3(new_n631), .A4(new_n695), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n642), .A2(new_n654), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT108), .Z(new_n788));
  NOR2_X1   g602(.A1(new_n785), .A2(new_n786), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT109), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n583), .A2(new_n326), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n792), .A2(G472), .B1(new_n559), .B2(new_n583), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n679), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n798), .B(new_n772), .C1(new_n797), .C2(new_n795), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n729), .B1(new_n513), .B2(new_n514), .ZN(new_n800));
  OAI22_X1  g614(.A1(new_n800), .A2(new_n497), .B1(new_n728), .B2(new_n508), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n449), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  INV_X1    g618(.A(new_n450), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(KEYINPUT46), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n516), .B1(new_n806), .B2(KEYINPUT46), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n447), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n809), .A2(new_n716), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n799), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n454), .ZN(G39));
  XNOR2_X1  g627(.A(new_n809), .B(KEYINPUT111), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT47), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n585), .A2(new_n631), .A3(new_n721), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n772), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  AND2_X1   g632(.A1(new_n734), .A2(new_n516), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n447), .A2(new_n446), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n821), .A2(new_n822), .A3(new_n785), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n712), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n699), .A2(new_n631), .A3(new_n703), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n401), .A2(new_n439), .A3(new_n694), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n779), .A2(new_n585), .A3(new_n688), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT113), .B1(new_n762), .B2(new_n779), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n792), .A2(G472), .B1(new_n559), .B2(new_n749), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n759), .A3(new_n710), .A4(new_n760), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n832), .A2(new_n767), .A3(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n783), .B(new_n829), .C1(new_n830), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n775), .B2(new_n780), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n345), .A2(new_n446), .A3(new_n656), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n793), .A2(new_n631), .A3(new_n517), .A4(new_n641), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n518), .A2(new_n632), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(KEYINPUT112), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(KEYINPUT112), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n840), .A2(new_n841), .A3(new_n747), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n663), .A2(new_n659), .A3(new_n444), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n672), .A3(new_n667), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n685), .A3(new_n754), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n736), .B1(new_n657), .B2(new_n668), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n836), .A2(new_n842), .A3(KEYINPUT114), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n689), .B1(new_n696), .B2(new_n722), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n638), .A2(new_n640), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n706), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n517), .A2(new_n679), .A3(new_n693), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n763), .A2(new_n849), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n763), .A2(new_n849), .A3(KEYINPUT52), .A4(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n848), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n742), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n756), .A2(new_n862), .B1(new_n839), .B2(KEYINPUT112), .ZN(new_n863));
  INV_X1    g677(.A(new_n841), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n847), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT114), .B1(new_n865), .B2(new_n836), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n861), .B2(new_n866), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n865), .A4(new_n836), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n869), .B1(KEYINPUT54), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n692), .B1(new_n788), .B2(new_n790), .ZN(new_n875));
  INV_X1    g689(.A(new_n751), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n756), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT119), .ZN(new_n880));
  INV_X1    g694(.A(G952), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n772), .A2(new_n735), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT117), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n883), .A2(new_n441), .A3(new_n826), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n881), .B(G953), .C1(new_n884), .C2(new_n656), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n886), .A2(KEYINPUT120), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n825), .A2(new_n707), .A3(new_n735), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n877), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT50), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n820), .A2(new_n447), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n772), .B(new_n878), .C1(new_n815), .C2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n401), .A2(new_n654), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n875), .A2(new_n883), .ZN(new_n897));
  INV_X1    g711(.A(new_n757), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n884), .A2(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n893), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT51), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n777), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT48), .Z(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n886), .B2(KEYINPUT120), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n899), .A2(KEYINPUT118), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(new_n901), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n899), .A2(KEYINPUT118), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n893), .A2(new_n895), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n887), .A2(new_n902), .A3(new_n905), .A4(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n874), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(G952), .A2(G953), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n827), .B1(new_n911), .B2(new_n912), .ZN(G75));
  NOR2_X1   g727(.A1(new_n306), .A2(G952), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n871), .A2(new_n872), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n326), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n269), .B(KEYINPUT121), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(new_n308), .Z(new_n921));
  OAI21_X1  g735(.A(new_n915), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n918), .B2(new_n921), .ZN(G51));
  XNOR2_X1  g737(.A(new_n873), .B(KEYINPUT54), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n450), .B(KEYINPUT57), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n732), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n916), .A2(new_n326), .A3(new_n804), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n914), .B1(new_n927), .B2(new_n928), .ZN(G54));
  AND2_X1   g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n917), .A2(new_n396), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n396), .B1(new_n917), .B2(new_n930), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n914), .ZN(G60));
  OR2_X1    g747(.A1(new_n649), .A2(new_n651), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n646), .ZN(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n874), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n924), .A2(new_n935), .A3(new_n937), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n914), .A3(new_n939), .ZN(G63));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n427), .A2(new_n326), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n871), .B2(new_n872), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n941), .B(new_n915), .C1(new_n946), .C2(new_n629), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n915), .B1(new_n946), .B2(new_n629), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n676), .A2(new_n677), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n873), .A2(new_n951), .A3(new_n944), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT124), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n628), .B1(new_n916), .B2(new_n945), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n946), .A2(new_n951), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n954), .A2(new_n955), .A3(new_n915), .A4(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n949), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  AOI22_X1  g772(.A1(new_n957), .A2(new_n953), .B1(new_n948), .B2(new_n947), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(G66));
  NAND2_X1  g774(.A1(new_n842), .A2(new_n847), .ZN(new_n961));
  NAND2_X1  g775(.A1(G224), .A2(G953), .ZN(new_n962));
  OAI22_X1  g776(.A1(new_n961), .A2(G953), .B1(new_n443), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(G898), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n919), .B1(new_n964), .B2(G953), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G69));
  NAND2_X1  g780(.A1(new_n536), .A2(new_n538), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n546), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(new_n391), .ZN(new_n969));
  INV_X1    g783(.A(new_n812), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n763), .A2(new_n849), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n777), .A2(new_n640), .A3(new_n638), .A4(new_n705), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n971), .B(new_n783), .C1(new_n810), .C2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n775), .B2(new_n780), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n970), .A2(new_n817), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n306), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n306), .A2(G900), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n977), .B1(new_n976), .B2(new_n979), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n969), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(G227), .A2(G900), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(G953), .ZN(new_n985));
  INV_X1    g799(.A(new_n969), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n970), .A2(new_n817), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n719), .A2(new_n971), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n772), .B1(new_n656), .B2(new_n667), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(new_n632), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n717), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n988), .B2(KEYINPUT62), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n987), .A2(new_n989), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n986), .B1(new_n994), .B2(G953), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n983), .A2(new_n985), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n976), .A2(new_n979), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n980), .ZN(new_n999));
  OAI211_X1 g813(.A(G953), .B(new_n984), .C1(new_n999), .C2(new_n986), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(G72));
  XNOR2_X1  g815(.A(new_n563), .B(KEYINPUT127), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n994), .A2(new_n865), .ZN(new_n1003));
  XNOR2_X1  g817(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n662), .A2(new_n326), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n524), .B(new_n1002), .C1(new_n1003), .C2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n578), .B1(new_n524), .B2(new_n563), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n868), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1006), .B1(new_n975), .B2(new_n961), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1002), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n580), .A3(new_n1012), .ZN(new_n1013));
  AND4_X1   g827(.A1(new_n915), .A2(new_n1008), .A3(new_n1010), .A4(new_n1013), .ZN(G57));
endmodule


