//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n202));
  AND2_X1   g001(.A1(G15gat), .A2(G22gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G15gat), .A2(G22gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(new_n203), .B2(new_n204), .ZN(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT91), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G8gat), .ZN(new_n211));
  OAI221_X1 g010(.A(new_n206), .B1(new_n202), .B2(G1gat), .C1(new_n203), .C2(new_n204), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n210), .A2(G8gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n214), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n209), .A2(new_n216), .A3(new_n211), .A4(new_n212), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219));
  INV_X1    g018(.A(G43gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G50gat), .ZN(new_n221));
  INV_X1    g020(.A(G50gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G43gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(G43gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(G50gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT86), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(KEYINPUT15), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT14), .ZN(new_n229));
  INV_X1    g028(.A(G29gat), .ZN(new_n230));
  INV_X1    g029(.A(G36gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n221), .A2(KEYINPUT88), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT15), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(new_n226), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n235), .B(new_n236), .C1(new_n237), .C2(KEYINPUT88), .ZN(new_n238));
  NAND2_X1  g037(.A1(G29gat), .A2(G36gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT89), .Z(new_n240));
  NAND4_X1  g039(.A1(new_n228), .A2(new_n234), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(KEYINPUT87), .A3(new_n233), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT87), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n239), .A3(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n246), .A2(KEYINPUT15), .A3(new_n227), .A4(new_n224), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n241), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n242), .B1(new_n241), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n218), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n241), .A2(new_n247), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(new_n215), .A3(new_n217), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n252), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n218), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(KEYINPUT92), .A3(new_n253), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n251), .B(KEYINPUT13), .Z(new_n260));
  INV_X1    g059(.A(KEYINPUT92), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n261), .A3(new_n218), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n251), .A4(new_n253), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n256), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT11), .B(G169gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(G197gat), .ZN(new_n267));
  XOR2_X1   g066(.A(G113gat), .B(G141gat), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT12), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n256), .A2(new_n263), .A3(new_n270), .A4(new_n264), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G230gat), .A2(G233gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(G99gat), .A2(G106gat), .ZN(new_n277));
  INV_X1    g076(.A(G85gat), .ZN(new_n278));
  INV_X1    g077(.A(G92gat), .ZN(new_n279));
  AOI22_X1  g078(.A1(KEYINPUT8), .A2(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT7), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n278), .B2(new_n279), .ZN(new_n282));
  NAND3_X1  g081(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(G99gat), .A2(G106gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n277), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n277), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n280), .A2(new_n287), .A3(new_n282), .A4(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G71gat), .ZN(new_n290));
  INV_X1    g089(.A(G78gat), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT93), .ZN(new_n292));
  NAND2_X1  g091(.A1(G71gat), .A2(G78gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G71gat), .A2(G78gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(KEYINPUT93), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G64gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT94), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G64gat), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n298), .A2(new_n300), .A3(G57gat), .ZN(new_n301));
  AOI21_X1  g100(.A(G57gat), .B1(new_n298), .B2(new_n300), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n293), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n296), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(KEYINPUT96), .A2(G64gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(KEYINPUT96), .A2(G64gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT95), .ZN(new_n310));
  INV_X1    g109(.A(G57gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n290), .A2(new_n291), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n293), .B1(new_n313), .B2(new_n304), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n307), .A2(KEYINPUT95), .A3(G57gat), .A4(new_n308), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n289), .B1(new_n306), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT99), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n300), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n311), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n298), .A2(new_n300), .A3(G57gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n305), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n296), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n288), .A4(new_n286), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n317), .A2(new_n318), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n325), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(KEYINPUT99), .A3(new_n289), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT10), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n276), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n329), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n334), .A2(new_n276), .ZN(new_n335));
  XNOR2_X1  g134(.A(G120gat), .B(G148gat), .ZN(new_n336));
  INV_X1    g135(.A(G176gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G204gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n333), .A2(new_n335), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n276), .B(KEYINPUT100), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n330), .B2(new_n332), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n344), .A2(new_n335), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(new_n345), .B2(new_n341), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n275), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT75), .B(KEYINPUT6), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(G141gat), .B(G148gat), .Z(new_n353));
  INV_X1    g152(.A(G155gat), .ZN(new_n354));
  INV_X1    g153(.A(G162gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT2), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G155gat), .B(G162gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n353), .A2(new_n358), .A3(new_n356), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT1), .ZN(new_n363));
  XNOR2_X1  g162(.A(G127gat), .B(G134gat), .ZN(new_n364));
  INV_X1    g163(.A(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G113gat), .ZN(new_n366));
  INV_X1    g165(.A(G113gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G120gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT67), .B1(new_n367), .B2(G120gat), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n363), .B(new_n364), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n364), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n366), .A2(new_n368), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(KEYINPUT1), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n362), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n361), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n372), .A2(new_n375), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n352), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n376), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n360), .A2(new_n361), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n386), .B(new_n379), .C1(new_n362), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n383), .B1(new_n382), .B2(new_n351), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT5), .B(new_n381), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n382), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n392), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n380), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n352), .A2(KEYINPUT5), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n393), .A2(new_n388), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G85gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n350), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT76), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n398), .A2(new_n403), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n407), .B(new_n350), .C1(new_n398), .C2(new_n403), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI211_X1 g208(.A(new_n402), .B(new_n350), .C1(new_n391), .C2(new_n397), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G197gat), .B(G204gat), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n412), .B1(KEYINPUT70), .B2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n413), .A2(KEYINPUT70), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G211gat), .B(G218gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT71), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n418), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G183gat), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT27), .B1(new_n427), .B2(KEYINPUT66), .ZN(new_n428));
  INV_X1    g227(.A(G190gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G183gat), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n428), .B(new_n429), .C1(KEYINPUT66), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT28), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT27), .B(G183gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(G190gat), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G169gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n337), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT26), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(G169gat), .B2(G176gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n427), .A2(new_n429), .ZN(new_n443));
  NOR4_X1   g242(.A1(new_n436), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(KEYINPUT23), .ZN(new_n446));
  OR3_X1    g245(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n446), .A2(new_n447), .B1(G169gat), .B2(G176gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI22_X1  g249(.A1(new_n450), .A2(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT24), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n427), .B2(new_n429), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT65), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n449), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n448), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT25), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT64), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n453), .B1(new_n450), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n453), .A2(new_n459), .B1(G183gat), .B2(G190gat), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n448), .B(new_n458), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT29), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n426), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n425), .B1(new_n445), .B2(new_n464), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n424), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n426), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n445), .B2(new_n464), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n470), .B(new_n423), .C1(new_n426), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G64gat), .B(G92gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT72), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(G8gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G36gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n469), .A2(new_n477), .A3(new_n472), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n473), .A2(new_n482), .A3(new_n478), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n409), .A2(new_n411), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT68), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n445), .A2(new_n464), .A3(new_n379), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n457), .A2(new_n463), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n376), .B1(new_n487), .B2(new_n444), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G227gat), .ZN(new_n490));
  INV_X1    g289(.A(G233gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n485), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n492), .A4(new_n488), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(new_n493), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT34), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n489), .A2(new_n501), .A3(new_n493), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G43gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n504), .B(new_n505), .Z(new_n506));
  NAND3_X1  g305(.A1(new_n498), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT33), .B1(new_n494), .B2(new_n495), .ZN(new_n508));
  INV_X1    g307(.A(new_n506), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n500), .B(new_n502), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT32), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G78gat), .B(G106gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT31), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(new_n222), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT77), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n419), .A2(new_n466), .A3(new_n422), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n362), .B1(new_n519), .B2(new_n387), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n386), .A2(new_n466), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n423), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(G228gat), .B(G233gat), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n466), .B1(new_n417), .B2(new_n418), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n416), .A2(new_n420), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n385), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n526), .A2(new_n378), .B1(G228gat), .B2(G233gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n522), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G22gat), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n530), .B1(new_n523), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n518), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n517), .A2(KEYINPUT77), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(KEYINPUT78), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n535), .B(new_n518), .C1(new_n531), .C2(new_n532), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n512), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n507), .A2(new_n510), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n484), .A2(new_n513), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT35), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n507), .A2(new_n510), .A3(new_n540), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n507), .B2(new_n510), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n397), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n389), .A2(new_n390), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n381), .A2(KEYINPUT5), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n349), .B1(new_n550), .B2(new_n402), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n402), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n398), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n410), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n481), .A2(new_n483), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n559));
  AND3_X1   g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n546), .A2(new_n560), .A3(new_n539), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n393), .A2(new_n388), .A3(new_n395), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n352), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n380), .A2(new_n352), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n564), .B(KEYINPUT39), .C1(new_n566), .C2(new_n377), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT80), .B(KEYINPUT39), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n352), .A3(new_n568), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n569), .A2(KEYINPUT81), .A3(new_n553), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT81), .B1(new_n569), .B2(new_n553), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT82), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(KEYINPUT40), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI221_X1 g374(.A(new_n567), .B1(new_n573), .B2(KEYINPUT40), .C1(new_n570), .C2(new_n571), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(new_n555), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n577), .A2(new_n558), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT83), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n473), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n469), .A2(KEYINPUT37), .A3(new_n472), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n477), .A4(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n581), .A2(new_n477), .A3(new_n583), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT38), .B1(new_n473), .B2(new_n478), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n556), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n578), .A2(new_n579), .A3(new_n539), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n556), .A2(new_n584), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n583), .A2(new_n477), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n586), .B1(new_n590), .B2(new_n581), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n539), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n558), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT83), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT69), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n598), .B(new_n599), .C1(new_n544), .C2(new_n545), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n513), .A2(new_n596), .A3(new_n597), .A4(new_n541), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n600), .B(new_n601), .C1(new_n539), .C2(new_n484), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n562), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT85), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n562), .B(KEYINPUT85), .C1(new_n595), .C2(new_n602), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n348), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  INV_X1    g407(.A(G211gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n328), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n218), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(G183gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n427), .A3(new_n218), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n614), .A2(new_n620), .A3(new_n615), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n619), .B1(new_n617), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n610), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n617), .A2(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n618), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n627));
  INV_X1    g426(.A(new_n610), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n624), .A2(new_n629), .A3(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n289), .B1(new_n248), .B2(new_n249), .ZN(new_n638));
  NAND3_X1  g437(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n289), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n252), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT98), .ZN(new_n643));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n638), .A2(new_n646), .A3(new_n639), .A4(new_n641), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n643), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n645), .B1(new_n643), .B2(new_n647), .ZN(new_n649));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n639), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n252), .A2(KEYINPUT17), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n241), .A2(new_n242), .A3(new_n247), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n655), .B1(new_n658), .B2(new_n289), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n646), .B1(new_n659), .B2(new_n641), .ZN(new_n660));
  INV_X1    g459(.A(new_n647), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n644), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n643), .A2(new_n645), .A3(new_n647), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n652), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n637), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n607), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n409), .A2(new_n411), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT101), .B(G1gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1324gat));
  OAI21_X1  g471(.A(G8gat), .B1(new_n667), .B2(new_n558), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n667), .ZN(new_n676));
  INV_X1    g475(.A(new_n558), .ZN(new_n677));
  INV_X1    g476(.A(G8gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n202), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n202), .A2(new_n678), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n676), .A2(new_n677), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n675), .B1(new_n683), .B2(new_n684), .ZN(G1325gat));
  NAND2_X1  g484(.A1(new_n600), .A2(new_n601), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n676), .A2(G15gat), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(G15gat), .B1(new_n676), .B2(new_n546), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(G1326gat));
  NOR2_X1   g488(.A1(new_n667), .A2(new_n539), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(new_n665), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n605), .B2(new_n606), .ZN(new_n695));
  INV_X1    g494(.A(new_n637), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n348), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n669), .A2(G29gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n693), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n703), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(KEYINPUT45), .A3(new_n701), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n654), .B2(new_n664), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n653), .B1(new_n648), .B2(new_n649), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n662), .A2(new_n652), .A3(new_n663), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT106), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n603), .A2(new_n707), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n695), .B2(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n333), .A2(new_n335), .A3(new_n341), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n341), .B1(new_n344), .B2(new_n335), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT104), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n696), .A2(new_n275), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n716), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n722), .B2(new_n669), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n704), .A2(new_n706), .A3(new_n723), .ZN(G1328gat));
  OAI21_X1  g523(.A(G36gat), .B1(new_n722), .B2(new_n558), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n558), .A2(G36gat), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n695), .A2(new_n726), .A3(new_n697), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT107), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n698), .A2(new_n727), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n725), .B(new_n729), .C1(new_n726), .C2(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n686), .A3(new_n720), .A4(new_n721), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G43gat), .ZN(new_n734));
  AND4_X1   g533(.A1(new_n220), .A2(new_n695), .A3(new_n546), .A4(new_n697), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n732), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g536(.A(KEYINPUT47), .B(new_n735), .C1(new_n733), .C2(G43gat), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(G1330gat));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740));
  INV_X1    g539(.A(new_n539), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n716), .A2(new_n741), .A3(new_n720), .A4(new_n721), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G50gat), .ZN(new_n743));
  AND4_X1   g542(.A1(new_n222), .A2(new_n695), .A3(new_n741), .A4(new_n697), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n740), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  AOI211_X1 g545(.A(KEYINPUT48), .B(new_n744), .C1(new_n742), .C2(G50gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(G1331gat));
  AND3_X1   g547(.A1(new_n603), .A2(new_n666), .A3(new_n275), .ZN(new_n749));
  INV_X1    g548(.A(new_n720), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n669), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n311), .ZN(G1332gat));
  XNOR2_X1  g552(.A(new_n558), .B(KEYINPUT108), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  XOR2_X1   g558(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n751), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n290), .B1(new_n762), .B2(new_n686), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n546), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766));
  INV_X1    g565(.A(new_n546), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n751), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n761), .B(new_n764), .C1(new_n769), .C2(G71gat), .ZN(new_n770));
  AOI21_X1  g569(.A(G71gat), .B1(new_n765), .B2(new_n768), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n760), .B1(new_n771), .B2(new_n763), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1334gat));
  NOR2_X1   g572(.A1(new_n751), .A2(new_n539), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(new_n291), .ZN(G1335gat));
  NAND2_X1  g574(.A1(new_n637), .A2(new_n275), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT111), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(new_n346), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n716), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n669), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n603), .A3(new_n665), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT112), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  OR3_X1    g583(.A1(new_n781), .A2(KEYINPUT112), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n346), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n668), .A2(new_n278), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n780), .B1(new_n786), .B2(new_n787), .ZN(G1336gat));
  OAI21_X1  g587(.A(G92gat), .B1(new_n779), .B2(new_n754), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n754), .A2(G92gat), .A3(new_n720), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n783), .A2(new_n785), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n716), .A2(new_n677), .A3(new_n778), .ZN(new_n794));
  INV_X1    g593(.A(new_n782), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n794), .A2(G92gat), .B1(new_n795), .B2(new_n792), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n791), .A2(new_n793), .B1(new_n790), .B2(new_n796), .ZN(G1337gat));
  INV_X1    g596(.A(new_n686), .ZN(new_n798));
  OAI21_X1  g597(.A(G99gat), .B1(new_n779), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n767), .A2(G99gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n786), .B2(new_n800), .ZN(G1338gat));
  NOR3_X1   g600(.A1(new_n720), .A2(G106gat), .A3(new_n539), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n783), .A2(new_n785), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n716), .A2(new_n741), .A3(new_n778), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(G106gat), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n806), .A2(G106gat), .B1(new_n795), .B2(new_n802), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n805), .A2(new_n807), .B1(new_n808), .B2(new_n804), .ZN(G1339gat));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n810), .B(new_n343), .C1(new_n330), .C2(new_n332), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n340), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n334), .A2(new_n331), .ZN(new_n813));
  INV_X1    g612(.A(new_n343), .ZN(new_n814));
  INV_X1    g613(.A(new_n332), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(KEYINPUT54), .A3(new_n333), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT114), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n821), .B(KEYINPUT55), .C1(new_n812), .C2(new_n817), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n340), .A4(new_n811), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n812), .A2(KEYINPUT113), .A3(new_n817), .A4(KEYINPUT55), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n717), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n828), .A3(new_n274), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n260), .B1(new_n259), .B2(new_n262), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n251), .B1(new_n250), .B2(new_n253), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n269), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n273), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n346), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n713), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  AND4_X1   g634(.A1(new_n713), .A2(new_n828), .A3(new_n823), .A4(new_n833), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n637), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n635), .A2(new_n636), .A3(new_n694), .A4(new_n275), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(new_n346), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n544), .A2(new_n741), .A3(new_n545), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n668), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n754), .ZN(new_n844));
  OAI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n275), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n274), .A2(new_n367), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT115), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n844), .B2(new_n847), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n844), .B2(new_n720), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n843), .A2(new_n365), .A3(new_n754), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n719), .B2(new_n850), .ZN(G1341gat));
  NOR2_X1   g650(.A1(new_n844), .A2(new_n637), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(G127gat), .Z(G1342gat));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n694), .A2(new_n677), .A3(G134gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n843), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n665), .A3(new_n754), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n857), .A2(new_n858), .B1(G134gat), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n854), .B1(new_n843), .B2(new_n855), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1343gat));
  NAND2_X1  g662(.A1(new_n840), .A2(new_n668), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT120), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n686), .A2(new_n539), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT121), .Z(new_n867));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n840), .A2(new_n868), .A3(new_n668), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n865), .A2(new_n754), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(G141gat), .A3(new_n275), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(G141gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n798), .A2(new_n668), .A3(new_n754), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n826), .A2(new_n827), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n818), .A2(new_n819), .B1(new_n272), .B2(new_n273), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n342), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n273), .A2(new_n832), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT118), .B1(new_n719), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n346), .A2(new_n833), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n665), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n637), .B1(new_n836), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n539), .B1(new_n885), .B2(new_n839), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n875), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT57), .B(new_n539), .C1(new_n837), .C2(new_n839), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(new_n275), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n872), .B1(new_n873), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT119), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n539), .B1(new_n837), .B2(new_n839), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n887), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n838), .A2(new_n346), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n713), .A2(new_n828), .A3(new_n823), .A4(new_n833), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n882), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n828), .B2(new_n877), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(new_n665), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n895), .B1(new_n899), .B2(new_n637), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n539), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n894), .A2(new_n901), .A3(new_n902), .A4(new_n875), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n873), .B1(new_n904), .B2(new_n274), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT58), .B1(new_n905), .B2(new_n871), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n906), .ZN(G1344gat));
  OR2_X1    g706(.A1(new_n893), .A2(new_n887), .ZN(new_n908));
  AND4_X1   g707(.A1(new_n665), .A2(new_n823), .A3(new_n828), .A4(new_n833), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n637), .B1(new_n909), .B2(new_n884), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n910), .A2(new_n839), .A3(KEYINPUT123), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT123), .B1(new_n910), .B2(new_n839), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n887), .B(new_n741), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  AND4_X1   g712(.A1(new_n346), .A2(new_n908), .A3(new_n913), .A4(new_n875), .ZN(new_n914));
  INV_X1    g713(.A(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT59), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT119), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n878), .A2(new_n883), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n694), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n696), .B1(new_n919), .B2(new_n896), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n741), .B1(new_n920), .B2(new_n895), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n874), .B1(new_n921), .B2(KEYINPUT57), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n902), .B1(new_n922), .B2(new_n894), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n346), .B1(new_n917), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n915), .A2(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT122), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n719), .B1(new_n892), .B2(new_n903), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  INV_X1    g727(.A(new_n925), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n916), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  OR3_X1    g730(.A1(new_n870), .A2(G148gat), .A3(new_n719), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1345gat));
  AOI21_X1  g732(.A(new_n637), .B1(new_n892), .B2(new_n903), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(new_n354), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n696), .A2(new_n354), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n870), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT124), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  OAI221_X1 g738(.A(new_n939), .B1(new_n870), .B2(new_n936), .C1(new_n934), .C2(new_n354), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n938), .A2(new_n940), .ZN(G1346gat));
  NOR3_X1   g740(.A1(new_n694), .A2(new_n677), .A3(G162gat), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n865), .A2(new_n867), .A3(new_n869), .A4(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n904), .A2(new_n713), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n355), .ZN(G1347gat));
  AOI211_X1 g744(.A(new_n668), .B(new_n754), .C1(new_n837), .C2(new_n839), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(new_n841), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n437), .A3(new_n274), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n669), .A2(new_n677), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT125), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n842), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G169gat), .B1(new_n951), .B2(new_n275), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n948), .A2(new_n952), .ZN(G1348gat));
  AOI21_X1  g752(.A(G176gat), .B1(new_n947), .B2(new_n346), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n951), .A2(new_n337), .A3(new_n720), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(new_n955), .ZN(G1349gat));
  NAND3_X1  g755(.A1(new_n947), .A2(new_n696), .A3(new_n434), .ZN(new_n957));
  OAI21_X1  g756(.A(G183gat), .B1(new_n951), .B2(new_n637), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n947), .A2(new_n429), .A3(new_n713), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n842), .A2(new_n665), .A3(new_n950), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n963), .A2(new_n964), .A3(G190gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n963), .B2(G190gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1351gat));
  NAND4_X1  g766(.A1(new_n908), .A2(new_n913), .A3(new_n798), .A4(new_n950), .ZN(new_n968));
  OAI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n275), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n946), .A2(new_n866), .ZN(new_n970));
  INV_X1    g769(.A(G197gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n275), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n969), .B(new_n975), .C1(new_n972), .C2(new_n275), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(G1352gat));
  NAND3_X1  g776(.A1(new_n970), .A2(new_n339), .A3(new_n346), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  OAI21_X1  g778(.A(G204gat), .B1(new_n968), .B2(new_n720), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(G1353gat));
  NAND3_X1  g781(.A1(new_n970), .A2(new_n609), .A3(new_n696), .ZN(new_n983));
  OR2_X1    g782(.A1(new_n968), .A2(new_n637), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n985));
  OAI211_X1 g784(.A(KEYINPUT63), .B(G211gat), .C1(new_n968), .C2(new_n637), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n983), .B1(new_n985), .B2(new_n987), .ZN(G1354gat));
  OAI21_X1  g787(.A(G218gat), .B1(new_n968), .B2(new_n694), .ZN(new_n989));
  INV_X1    g788(.A(G218gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n970), .A2(new_n990), .A3(new_n713), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(G1355gat));
endmodule


