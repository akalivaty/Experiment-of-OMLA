//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(G36gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT17), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  INV_X1    g015(.A(G1gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(KEYINPUT16), .A3(new_n217), .ZN(new_n218));
  OAI221_X1 g017(.A(new_n218), .B1(KEYINPUT92), .B2(G8gat), .C1(new_n217), .C2(new_n216), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n220));
  XOR2_X1   g019(.A(new_n219), .B(new_n220), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n219), .B(new_n220), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n214), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT93), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(KEYINPUT18), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(KEYINPUT94), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n224), .A2(new_n214), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n223), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(KEYINPUT18), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n228), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT11), .B(G169gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n228), .A2(new_n242), .A3(new_n233), .A4(new_n234), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT102), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT9), .ZN(new_n246));
  INV_X1    g045(.A(G71gat), .ZN(new_n247));
  INV_X1    g046(.A(G78gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT96), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(G57gat), .B(G64gat), .Z(new_n252));
  XNOR2_X1  g051(.A(G71gat), .B(G78gat), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT96), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT97), .ZN(new_n256));
  INV_X1    g055(.A(new_n253), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n257), .A2(KEYINPUT95), .B1(new_n252), .B2(new_n249), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(KEYINPUT95), .B2(new_n257), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT98), .B(KEYINPUT21), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G231gat), .A2(G233gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G127gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G183gat), .B(G211gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n221), .B1(new_n268), .B2(new_n260), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n269), .B(KEYINPUT99), .Z(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n271));
  INV_X1    g070(.A(G155gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n270), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n266), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n265), .B(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n270), .B(new_n273), .Z(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G85gat), .A2(G92gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT7), .ZN(new_n282));
  NAND2_X1  g081(.A1(G99gat), .A2(G106gat), .ZN(new_n283));
  INV_X1    g082(.A(G85gat), .ZN(new_n284));
  INV_X1    g083(.A(G92gat), .ZN(new_n285));
  AOI22_X1  g084(.A1(KEYINPUT8), .A2(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G99gat), .B(G106gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n215), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(G232gat), .A2(G233gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n214), .A2(new_n289), .B1(KEYINPUT41), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G190gat), .B(G218gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n292), .A2(KEYINPUT41), .ZN(new_n297));
  XNOR2_X1  g096(.A(G134gat), .B(G162gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n299), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n280), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n260), .B(new_n290), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n256), .A2(new_n289), .A3(KEYINPUT10), .A4(new_n259), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n306), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT100), .ZN(new_n313));
  XOR2_X1   g112(.A(G120gat), .B(G148gat), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT101), .ZN(new_n315));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(KEYINPUT100), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n310), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n317), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n310), .B2(new_n312), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n245), .B1(new_n304), .B2(new_n325), .ZN(new_n326));
  NOR4_X1   g125(.A1(new_n280), .A2(new_n303), .A3(KEYINPUT102), .A4(new_n324), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n244), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(KEYINPUT74), .B(G71gat), .Z(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(G99gat), .ZN(new_n330));
  XOR2_X1   g129(.A(G15gat), .B(G43gat), .Z(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n336));
  NOR3_X1   g135(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(KEYINPUT70), .ZN(new_n338));
  INV_X1    g137(.A(G169gat), .ZN(new_n339));
  INV_X1    g138(.A(G176gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT26), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n334), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT71), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT69), .ZN(new_n347));
  AND2_X1   g146(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n352));
  AND4_X1   g151(.A1(new_n347), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n350), .A2(new_n351), .B1(new_n347), .B2(new_n352), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(KEYINPUT71), .B(new_n334), .C1(new_n338), .C2(new_n343), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n346), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359));
  INV_X1    g158(.A(G113gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G113gat), .B(G120gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G113gat), .B(G120gat), .Z(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n359), .ZN(new_n367));
  INV_X1    g166(.A(new_n358), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n362), .A2(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n334), .A2(KEYINPUT24), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT24), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(G183gat), .A3(G190gat), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n341), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(G176gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT64), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n339), .ZN(new_n380));
  NAND2_X1  g179(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n374), .B1(new_n383), .B2(KEYINPUT65), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT65), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n377), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT25), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n388), .A2(KEYINPUT23), .B1(new_n335), .B2(KEYINPUT66), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n341), .A2(new_n376), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n335), .A2(KEYINPUT66), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .A4(KEYINPUT25), .ZN(new_n392));
  OR2_X1    g191(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n393));
  INV_X1    g192(.A(G183gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT68), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n350), .A2(KEYINPUT68), .A3(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n371), .A2(new_n373), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n392), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n357), .B(new_n369), .C1(new_n387), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT73), .ZN(new_n404));
  INV_X1    g203(.A(new_n402), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n340), .A2(KEYINPUT23), .ZN(new_n406));
  AND2_X1   g205(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n335), .B1(new_n388), .B2(KEYINPUT23), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT65), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n374), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n386), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT25), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n405), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT73), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n369), .A4(new_n357), .ZN(new_n418));
  INV_X1    g217(.A(new_n354), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n350), .A2(new_n351), .A3(new_n347), .A4(new_n352), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n356), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n342), .B1(new_n341), .B2(KEYINPUT26), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n337), .A2(KEYINPUT70), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n335), .A4(new_n336), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT71), .B1(new_n424), .B2(new_n334), .ZN(new_n425));
  OAI22_X1  g224(.A1(new_n387), .A2(new_n402), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n362), .A2(new_n365), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n367), .A2(new_n368), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n404), .A2(new_n418), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n333), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n431), .B2(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  AOI221_X4 g239(.A(new_n437), .B1(KEYINPUT33), .B2(new_n332), .C1(new_n431), .C2(new_n433), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n404), .A2(new_n432), .A3(new_n418), .A4(new_n430), .ZN(new_n443));
  XOR2_X1   g242(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(KEYINPUT75), .A2(KEYINPUT34), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n443), .A2(new_n446), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n443), .B2(new_n444), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT33), .B1(new_n431), .B2(new_n433), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n438), .A2(new_n451), .A3(new_n333), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n452), .B2(new_n441), .ZN(new_n453));
  INV_X1    g252(.A(G148gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT83), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G148gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n457), .A3(G141gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n454), .A2(G141gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461));
  INV_X1    g260(.A(G162gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n272), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n458), .A2(new_n460), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT84), .B(G155gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G162gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT2), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT2), .ZN(new_n469));
  INV_X1    g268(.A(G141gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(G148gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n459), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n461), .A2(KEYINPUT82), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(G155gat), .A3(G162gat), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n473), .A2(new_n474), .A3(new_n463), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n464), .A2(new_n467), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT78), .ZN(new_n477));
  OR2_X1    g276(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT22), .B1(new_n480), .B2(G211gat), .ZN(new_n481));
  XOR2_X1   g280(.A(G197gat), .B(G204gat), .Z(new_n482));
  OAI21_X1  g281(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  INV_X1    g283(.A(G211gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n478), .B2(new_n479), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n484), .B(KEYINPUT78), .C1(KEYINPUT22), .C2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G211gat), .B(G218gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n481), .A2(new_n482), .ZN(new_n491));
  INV_X1    g290(.A(new_n488), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT78), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n489), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT3), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n476), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n464), .A2(new_n467), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n475), .A2(new_n472), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n490), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(KEYINPUT89), .A3(new_n490), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n493), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n502), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n502), .B2(new_n506), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n510), .A2(new_n496), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n497), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(G22gat), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n508), .B(new_n516), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT31), .B(G50gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n515), .A2(KEYINPUT90), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n524), .A2(new_n520), .B1(new_n515), .B2(new_n517), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n448), .B(new_n453), .C1(new_n522), .C2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT4), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n476), .A2(new_n527), .A3(new_n369), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT87), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n476), .A2(new_n369), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(KEYINPUT87), .A3(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n499), .A2(new_n500), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n369), .B1(new_n535), .B2(KEYINPUT3), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT85), .A3(new_n501), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT85), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n429), .B1(new_n476), .B2(new_n495), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n499), .A2(new_n495), .A3(new_n500), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G225gat), .A2(G233gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT5), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n534), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n528), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n527), .B1(new_n476), .B2(new_n369), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n541), .B2(new_n537), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n429), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT86), .A3(new_n530), .ZN(new_n552));
  OR3_X1    g351(.A1(new_n476), .A2(new_n369), .A3(KEYINPUT86), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n544), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT5), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n546), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G1gat), .B(G29gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT0), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G85gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n544), .B1(new_n531), .B2(new_n528), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT85), .B1(new_n536), .B2(new_n501), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n539), .A2(new_n540), .A3(new_n538), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(KEYINPUT5), .A3(new_n554), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n546), .A3(new_n560), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n556), .A2(KEYINPUT6), .A3(new_n561), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G226gat), .ZN(new_n573));
  INV_X1    g372(.A(G233gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n426), .B2(new_n490), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(new_n416), .B2(new_n357), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT79), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n506), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT79), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT29), .B1(new_n416), .B2(new_n357), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(new_n575), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n426), .A2(new_n575), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n582), .B2(new_n575), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n506), .ZN(new_n587));
  XNOR2_X1  g386(.A(G8gat), .B(G36gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G64gat), .B(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  AND3_X1   g391(.A1(new_n584), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n592), .B1(new_n584), .B2(new_n587), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n584), .A2(new_n587), .ZN(new_n597));
  INV_X1    g396(.A(new_n592), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n597), .A2(KEYINPUT30), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n572), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT35), .B1(new_n526), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n598), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n587), .A3(new_n592), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(KEYINPUT30), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n576), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n580), .B1(new_n605), .B2(new_n585), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n421), .A2(new_n425), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n396), .A2(new_n397), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT68), .B1(new_n350), .B2(new_n394), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n401), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n392), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n413), .A2(new_n414), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n490), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT79), .B1(new_n613), .B2(new_n577), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n586), .B2(KEYINPUT79), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n606), .B1(new_n615), .B2(new_n580), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n595), .A3(new_n592), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n604), .A2(new_n617), .B1(new_n571), .B2(new_n570), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n452), .A2(new_n450), .A3(new_n441), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n447), .B1(new_n440), .B2(new_n442), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT35), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n524), .A2(new_n520), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n515), .A2(new_n517), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n521), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n618), .A2(new_n621), .A3(new_n622), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n601), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n552), .A2(new_n553), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(new_n543), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n532), .A2(new_n533), .B1(new_n537), .B2(new_n541), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(new_n543), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n534), .A2(new_n542), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n629), .A3(new_n544), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n633), .A2(new_n635), .A3(KEYINPUT40), .A4(new_n560), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n560), .B1(new_n568), .B2(new_n546), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n635), .A3(new_n560), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n604), .A2(new_n617), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n579), .A2(new_n506), .A3(new_n583), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n586), .B2(new_n580), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n647), .B(new_n598), .C1(KEYINPUT37), .C2(new_n597), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n648), .A2(new_n571), .A3(new_n570), .A4(new_n603), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n592), .B1(new_n616), .B2(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n597), .A2(KEYINPUT37), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n642), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n641), .B(new_n626), .C1(new_n649), .C2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n522), .A2(new_n525), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n600), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT76), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n619), .B2(new_n620), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n453), .A2(new_n448), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n653), .A2(new_n655), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n328), .B1(new_n628), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n572), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT103), .B(G1gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1324gat));
  NOR2_X1   g468(.A1(new_n596), .A2(new_n599), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n671), .A2(G8gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT16), .B(G8gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT42), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(KEYINPUT42), .B2(new_n674), .ZN(G1325gat));
  INV_X1    g475(.A(G15gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n665), .A2(new_n677), .A3(new_n621), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT104), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n663), .A2(KEYINPUT104), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n665), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n678), .B1(new_n683), .B2(new_n677), .ZN(G1326gat));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n654), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT105), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n601), .A2(new_n689), .A3(new_n627), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n601), .B2(new_n627), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n664), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n302), .A2(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n628), .A2(new_n664), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n303), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n692), .A2(new_n693), .B1(new_n695), .B2(KEYINPUT44), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n280), .ZN(new_n698));
  INV_X1    g497(.A(new_n244), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n698), .A2(new_n699), .A3(new_n324), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n572), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n302), .B1(new_n628), .B2(new_n664), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(new_n700), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n206), .A3(new_n666), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n202), .A3(new_n670), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT46), .Z(new_n709));
  INV_X1    g508(.A(new_n670), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n701), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  INV_X1    g512(.A(G43gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n701), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n682), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n704), .A2(new_n714), .A3(new_n621), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n663), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT107), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n701), .A2(new_n721), .A3(new_n663), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n720), .A2(new_n714), .A3(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n717), .A2(new_n713), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n718), .B1(new_n723), .B2(new_n724), .ZN(G1330gat));
  OAI21_X1  g524(.A(G50gat), .B1(new_n701), .B2(new_n626), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT48), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n626), .A2(G50gat), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT108), .Z(new_n730));
  NAND2_X1  g529(.A1(new_n704), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n728), .B(new_n732), .ZN(G1331gat));
  NAND2_X1  g532(.A1(new_n304), .A2(new_n699), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n325), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n692), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n572), .B(KEYINPUT110), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g540(.A1(new_n736), .A2(new_n710), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  NOR4_X1   g545(.A1(new_n736), .A2(new_n247), .A3(new_n680), .A4(new_n681), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT111), .B1(new_n737), .B2(new_n621), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(G71gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n737), .A2(KEYINPUT111), .A3(new_n621), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n736), .A2(new_n626), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n248), .ZN(G1335gat));
  NAND2_X1  g554(.A1(new_n699), .A2(new_n280), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n325), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT113), .B1(new_n696), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  INV_X1    g559(.A(new_n693), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n628), .A2(KEYINPUT106), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n601), .A2(new_n627), .A3(new_n689), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n761), .B1(new_n764), .B2(new_n664), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n703), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n760), .B(new_n757), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n759), .A2(new_n666), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n284), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n302), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n692), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n692), .A2(KEYINPUT51), .A3(new_n773), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n324), .A2(new_n666), .A3(new_n284), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n772), .B1(new_n778), .B2(new_n779), .ZN(G1336gat));
  NOR4_X1   g579(.A1(new_n778), .A2(G92gat), .A3(new_n710), .A4(new_n325), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(KEYINPUT52), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n697), .A2(new_n757), .ZN(new_n783));
  OAI21_X1  g582(.A(G92gat), .B1(new_n783), .B2(new_n710), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n759), .A2(new_n670), .A3(new_n768), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n786), .A2(new_n787), .A3(G92gat), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n786), .B2(G92gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n788), .A2(new_n789), .A3(new_n781), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(G1337gat));
  NAND3_X1  g591(.A1(new_n759), .A2(new_n682), .A3(new_n768), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G99gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n621), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n795), .A2(new_n325), .A3(G99gat), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n778), .B2(new_n796), .ZN(G1338gat));
  OAI21_X1  g596(.A(G106gat), .B1(new_n783), .B2(new_n626), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n325), .A2(new_n626), .A3(G106gat), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n776), .B2(new_n777), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n759), .A2(new_n654), .A3(new_n768), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n802), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT116), .B1(new_n807), .B2(KEYINPUT53), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n801), .B1(new_n805), .B2(G106gat), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n809), .A2(new_n810), .A3(new_n803), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n804), .B1(new_n808), .B2(new_n811), .ZN(G1339gat));
  NOR2_X1   g611(.A1(new_n734), .A2(new_n324), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n310), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n322), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n308), .A2(new_n306), .A3(new_n309), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT117), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n310), .A2(new_n814), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(KEYINPUT55), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n231), .A2(new_n232), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n223), .B1(new_n222), .B2(new_n225), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n239), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT118), .B(new_n239), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n243), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n821), .A2(new_n828), .A3(new_n302), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n320), .B1(new_n820), .B2(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n324), .A2(new_n243), .A3(new_n827), .A4(new_n826), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n819), .ZN(new_n834));
  INV_X1    g633(.A(new_n816), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n836), .A2(new_n837), .B1(new_n241), .B2(new_n243), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n838), .B2(new_n830), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n831), .B1(new_n839), .B2(new_n303), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n813), .B1(new_n840), .B2(new_n280), .ZN(new_n841));
  NOR4_X1   g640(.A1(new_n841), .A2(new_n670), .A3(new_n526), .A4(new_n738), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n360), .A3(new_n244), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n841), .A2(new_n654), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n710), .A2(new_n666), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n795), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n244), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n844), .B1(new_n850), .B2(G113gat), .ZN(new_n851));
  AOI211_X1 g650(.A(KEYINPUT119), .B(new_n360), .C1(new_n849), .C2(new_n244), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n843), .B1(new_n851), .B2(new_n852), .ZN(G1340gat));
  AND3_X1   g652(.A1(new_n849), .A2(G120gat), .A3(new_n324), .ZN(new_n854));
  AOI21_X1  g653(.A(G120gat), .B1(new_n842), .B2(new_n324), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n848), .B2(new_n280), .ZN(new_n857));
  INV_X1    g656(.A(G127gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n858), .A3(new_n698), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1342gat));
  NOR2_X1   g659(.A1(new_n841), .A2(new_n738), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n302), .A2(new_n670), .A3(G134gat), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n626), .A3(new_n621), .A4(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n848), .B2(new_n302), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n719), .A2(new_n846), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n841), .A2(new_n869), .A3(new_n626), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n244), .B1(KEYINPUT55), .B2(new_n820), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n321), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n832), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AOI22_X1  g673(.A1(new_n874), .A2(new_n302), .B1(new_n830), .B2(new_n829), .ZN(new_n875));
  OAI22_X1  g674(.A1(new_n875), .A2(new_n698), .B1(new_n324), .B2(new_n734), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n654), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n244), .B(new_n868), .C1(new_n870), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G141gat), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT120), .B1(new_n682), .B2(new_n626), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n682), .A2(new_n626), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n861), .A2(new_n880), .A3(new_n710), .A4(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n699), .A2(G141gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n879), .A2(new_n887), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n868), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n869), .B1(new_n841), .B2(new_n626), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n876), .A2(KEYINPUT57), .A3(new_n654), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n470), .B1(new_n896), .B2(new_n244), .ZN(new_n897));
  INV_X1    g696(.A(new_n886), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n891), .B1(new_n884), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n889), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n892), .A2(new_n900), .ZN(G1344gat));
  OAI21_X1  g700(.A(new_n699), .B1(new_n326), .B2(new_n327), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n875), .B2(new_n698), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n903), .B2(new_n654), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n324), .B(new_n868), .C1(new_n870), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G148gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT59), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n455), .A2(new_n457), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(KEYINPUT59), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI211_X1 g711(.A(new_n908), .B(new_n912), .C1(new_n896), .C2(new_n324), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n324), .B(new_n868), .C1(new_n870), .C2(new_n877), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT122), .B1(new_n914), .B2(new_n911), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n907), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n885), .A2(new_n910), .A3(new_n324), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1345gat));
  AOI21_X1  g717(.A(new_n465), .B1(new_n885), .B2(new_n698), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n698), .A2(new_n465), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT123), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n896), .B2(new_n921), .ZN(G1346gat));
  AOI21_X1  g721(.A(new_n462), .B1(new_n896), .B2(new_n303), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n302), .A2(new_n670), .A3(G162gat), .ZN(new_n924));
  AND4_X1   g723(.A1(new_n861), .A2(new_n880), .A3(new_n883), .A4(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n923), .A2(new_n925), .ZN(G1347gat));
  NAND2_X1  g725(.A1(new_n738), .A2(new_n670), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n795), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n845), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n699), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n841), .A2(new_n666), .A3(new_n710), .A4(new_n526), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n931), .A2(new_n380), .A3(new_n381), .A4(new_n244), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1348gat));
  OAI21_X1  g732(.A(G176gat), .B1(new_n929), .B2(new_n325), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n340), .A3(new_n324), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  NAND2_X1  g735(.A1(new_n698), .A2(new_n351), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G183gat), .B1(new_n929), .B2(new_n280), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT124), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n931), .A2(new_n350), .A3(new_n303), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n845), .A2(new_n303), .A3(new_n928), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(G190gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n944), .B2(G190gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  NOR2_X1   g747(.A1(new_n841), .A2(new_n666), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n950), .B1(new_n881), .B2(new_n670), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n881), .A2(new_n950), .A3(new_n670), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n244), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n870), .A2(new_n904), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n682), .A2(new_n927), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n244), .A2(G197gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n324), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G204gat), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n325), .A2(G204gat), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n954), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT126), .A3(new_n964), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT126), .B1(new_n967), .B2(new_n964), .ZN(new_n969));
  OAI221_X1 g768(.A(new_n963), .B1(new_n964), .B2(new_n967), .C1(new_n968), .C2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n485), .A3(new_n698), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n958), .B(new_n698), .C1(new_n870), .C2(new_n904), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  AOI21_X1  g774(.A(G218gat), .B1(new_n955), .B2(new_n303), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n303), .A2(new_n480), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT127), .Z(new_n978));
  AOI21_X1  g777(.A(new_n976), .B1(new_n959), .B2(new_n978), .ZN(G1355gat));
endmodule


