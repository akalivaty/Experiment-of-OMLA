//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT66), .B1(new_n459), .B2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(new_n458), .A3(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n466), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AND4_X1   g045(.A1(G137), .A2(new_n460), .A3(new_n462), .A4(new_n458), .ZN(new_n471));
  NOR3_X1   g046(.A1(new_n465), .A2(new_n470), .A3(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n460), .A2(new_n462), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n458), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n458), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT67), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND4_X1  g057(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n458), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G138), .A4(new_n458), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n460), .A2(new_n462), .A3(G126), .A4(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT68), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n489), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n488), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n504), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XOR2_X1   g091(.A(new_n516), .B(KEYINPUT69), .Z(new_n517));
  AOI21_X1  g092(.A(new_n505), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n514), .A2(new_n518), .ZN(G166));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n510), .A2(new_n520), .B1(new_n512), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n522), .A2(new_n528), .ZN(G168));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT70), .B(G52), .Z(new_n531));
  OAI22_X1  g106(.A1(new_n510), .A2(new_n530), .B1(new_n512), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n505), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n532), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(new_n501), .A2(new_n503), .ZN(new_n537));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  INV_X1    g113(.A(G68), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n500), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT71), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  OAI221_X1 g117(.A(new_n542), .B1(new_n539), .B2(new_n500), .C1(new_n537), .C2(new_n538), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(G651), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n541), .A2(KEYINPUT72), .A3(new_n543), .A4(G651), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n506), .A2(new_n508), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n537), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n500), .ZN(new_n550));
  AOI22_X1  g125(.A1(G81), .A2(new_n549), .B1(new_n550), .B2(G43), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G860), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT73), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n501), .A2(new_n503), .A3(G65), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n563), .A2(KEYINPUT75), .A3(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n549), .A2(G91), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n509), .A2(new_n571), .A3(G53), .A4(G543), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n506), .A2(new_n508), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n572), .A2(new_n570), .A3(new_n574), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n568), .B(new_n569), .C1(new_n575), .C2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  INV_X1    g154(.A(G74), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n505), .B1(new_n537), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  AOI22_X1  g157(.A1(G87), .A2(new_n549), .B1(new_n550), .B2(G49), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n537), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  AOI22_X1  g164(.A1(G86), .A2(new_n549), .B1(new_n550), .B2(G48), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n510), .A2(new_n594), .B1(new_n512), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n537), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G651), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n596), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n605));
  OR4_X1    g180(.A1(new_n604), .A2(new_n537), .A3(new_n548), .A4(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n510), .B2(new_n604), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n550), .A2(G54), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n505), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(G168), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT79), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(KEYINPUT79), .B2(new_n617), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(KEYINPUT79), .B2(new_n617), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n613), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n613), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(new_n552), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(G868), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g204(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n630));
  XNOR2_X1  g205(.A(G323), .B(new_n630), .ZN(G282));
  NAND2_X1  g206(.A1(new_n467), .A2(new_n469), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n485), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n474), .A2(G123), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n476), .A2(G135), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n458), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n636), .A2(new_n637), .A3(new_n644), .ZN(G156));
  INV_X1    g220(.A(G14), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT83), .B(G2438), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  OR3_X1    g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n651), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n661), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1341), .B(G1348), .Z(new_n665));
  AOI21_X1  g240(.A(new_n646), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n664), .ZN(new_n667));
  INV_X1    g242(.A(new_n665), .ZN(new_n668));
  AOI21_X1  g243(.A(KEYINPUT84), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g244(.A(KEYINPUT84), .B(new_n668), .C1(new_n662), .C2(new_n663), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT87), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n677), .A2(new_n680), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2072), .B(G2078), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2100), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G2096), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(G2096), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n684), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n683), .A3(new_n691), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(G227));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1956), .B(G2474), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1961), .B(G1966), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1971), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT19), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n705), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n701), .A2(new_n702), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n706), .A2(KEYINPUT20), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n707), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(new_n703), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n709), .B(new_n711), .C1(KEYINPUT20), .C2(new_n706), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1991), .ZN(new_n713));
  INV_X1    g288(.A(G1996), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G1991), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n712), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G1996), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n698), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(G1996), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n713), .A2(new_n714), .ZN(new_n722));
  INV_X1    g297(.A(new_n698), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g299(.A1(new_n719), .A2(new_n720), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(new_n719), .B2(new_n724), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(G229));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G6), .ZN(new_n729));
  INV_X1    g304(.A(G305), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n728), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT32), .B(G1981), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G16), .A2(G23), .ZN(new_n734));
  INV_X1    g309(.A(G288), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G16), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT33), .B(G1976), .Z(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G22), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G166), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT91), .B(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n736), .A2(new_n737), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n733), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT34), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G24), .ZN(new_n747));
  XNOR2_X1  g322(.A(G290), .B(KEYINPUT90), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1986), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n474), .A2(G119), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n476), .A2(G131), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n458), .A2(G107), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  MUX2_X1   g330(.A(G25), .B(new_n755), .S(G29), .Z(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT35), .B(G1991), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n756), .B(new_n757), .Z(new_n758));
  NAND3_X1  g333(.A1(new_n746), .A2(new_n750), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT36), .ZN(new_n760));
  NAND2_X1  g335(.A1(G168), .A2(G16), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G16), .B2(G21), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT98), .Z(new_n765));
  NOR2_X1   g340(.A1(G29), .A2(G33), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n485), .A2(G127), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n458), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n769), .B(new_n772), .C1(G139), .C2(new_n476), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(G29), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(G2072), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT94), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n498), .A2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G29), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G27), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n778), .A2(G32), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT26), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G141), .B2(new_n476), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n474), .A2(G129), .B1(G105), .B2(new_n632), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(new_n778), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT97), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT27), .B(G1996), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n765), .A2(new_n776), .A3(new_n782), .A4(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n763), .A2(new_n762), .B1(new_n774), .B2(G2072), .ZN(new_n795));
  NAND2_X1  g370(.A1(G160), .A2(G29), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n797));
  INV_X1    g372(.A(G34), .ZN(new_n798));
  AOI21_X1  g373(.A(G29), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(KEYINPUT96), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n799), .A2(new_n802), .B1(new_n798), .B2(new_n797), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n796), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2084), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n795), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT30), .B(G28), .ZN(new_n807));
  OR2_X1    g382(.A1(KEYINPUT31), .A2(G11), .ZN(new_n808));
  NAND2_X1  g383(.A1(KEYINPUT31), .A2(G11), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n807), .A2(new_n778), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n642), .B2(new_n778), .ZN(new_n811));
  NAND2_X1  g386(.A1(G171), .A2(G16), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G5), .B2(G16), .ZN(new_n813));
  INV_X1    g388(.A(G1961), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G1348), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n613), .A2(G16), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G4), .B2(G16), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n806), .B(new_n815), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n813), .A2(new_n820), .A3(new_n814), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n818), .A2(new_n816), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n820), .B1(new_n813), .B2(new_n814), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n794), .A2(new_n819), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n728), .A2(G19), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n628), .B2(new_n728), .ZN(new_n827));
  MUX2_X1   g402(.A(new_n826), .B(new_n827), .S(KEYINPUT92), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G1341), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(G1341), .ZN(new_n830));
  INV_X1    g405(.A(G2067), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n778), .A2(G26), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n474), .A2(G128), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n476), .A2(G140), .ZN(new_n834));
  OR2_X1    g409(.A1(G104), .A2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n832), .B1(new_n837), .B2(G29), .ZN(new_n838));
  MUX2_X1   g413(.A(new_n832), .B(new_n838), .S(KEYINPUT28), .Z(new_n839));
  INV_X1    g414(.A(new_n780), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n831), .A2(new_n839), .B1(new_n840), .B2(G2078), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n841), .B1(new_n831), .B2(new_n839), .C1(new_n792), .C2(new_n791), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n778), .A2(G35), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G162), .B2(new_n778), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT29), .Z(new_n845));
  INV_X1    g420(.A(G2090), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n825), .A2(new_n829), .A3(new_n830), .A4(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n728), .A2(G20), .ZN(new_n850));
  NAND2_X1  g425(.A1(G299), .A2(G16), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(KEYINPUT23), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(KEYINPUT23), .B2(new_n850), .ZN(new_n853));
  INV_X1    g428(.A(G1956), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n849), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(KEYINPUT100), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(KEYINPUT100), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n848), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n760), .A2(new_n860), .ZN(G311));
  NAND2_X1  g436(.A1(new_n760), .A2(new_n860), .ZN(G150));
  INV_X1    g437(.A(G67), .ZN(new_n863));
  INV_X1    g438(.A(G80), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n537), .A2(new_n863), .B1(new_n864), .B2(new_n500), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT102), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  OAI221_X1 g442(.A(new_n867), .B1(new_n864), .B2(new_n500), .C1(new_n537), .C2(new_n863), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(G651), .A3(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(G93), .A2(new_n549), .B1(new_n550), .B2(G55), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(KEYINPUT103), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n869), .B2(new_n870), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G860), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT37), .Z(new_n877));
  OAI21_X1  g452(.A(new_n552), .B1(new_n872), .B2(new_n874), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n878), .A2(KEYINPUT104), .B1(new_n628), .B2(new_n871), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(new_n552), .C1(new_n872), .C2(new_n874), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT101), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT38), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n612), .A2(new_n624), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT39), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n553), .B1(new_n884), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n877), .B1(new_n888), .B2(new_n889), .ZN(G145));
  NAND2_X1  g465(.A1(new_n476), .A2(G142), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT106), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n458), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n474), .A2(G130), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n755), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT107), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n634), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n898), .B(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n634), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n494), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n488), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n837), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n789), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n773), .B(KEYINPUT105), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n908), .B(new_n788), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n773), .A2(KEYINPUT105), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n642), .B(G160), .Z(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(new_n481), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n911), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n918), .A2(new_n900), .A3(new_n904), .A4(new_n920), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n922), .A2(KEYINPUT108), .A3(new_n923), .A4(new_n924), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g505(.A(new_n882), .B(new_n626), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n612), .B(G299), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(KEYINPUT41), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n931), .ZN(new_n935));
  INV_X1    g510(.A(G290), .ZN(new_n936));
  NAND2_X1  g511(.A1(G305), .A2(G288), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(G305), .A2(G288), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n939), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(G290), .A3(new_n937), .ZN(new_n942));
  XNOR2_X1  g517(.A(G166), .B(KEYINPUT109), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n940), .B2(new_n942), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT42), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n935), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n935), .A2(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n875), .A2(new_n616), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(G295));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n951), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  XNOR2_X1  g529(.A(G286), .B(G301), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n879), .A2(new_n881), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n879), .B2(new_n881), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n934), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n882), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n932), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n956), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n946), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT110), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n959), .A2(new_n963), .A3(new_n946), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n946), .B1(new_n959), .B2(new_n963), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(G37), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n954), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(G397));
  AOI21_X1  g554(.A(G1384), .B1(new_n488), .B2(new_n906), .ZN(new_n980));
  INV_X1    g555(.A(new_n465), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n471), .A2(new_n470), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n982), .A3(G40), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n980), .A2(new_n983), .A3(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n714), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT112), .Z(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT46), .Z(new_n987));
  XNOR2_X1  g562(.A(new_n837), .B(G2067), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n988), .B2(new_n788), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n789), .A2(new_n714), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n986), .A2(new_n789), .B1(new_n984), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n755), .A2(new_n757), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n984), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n984), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n1000), .A2(G1986), .A3(G290), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT48), .Z(new_n1002));
  NAND2_X1  g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n837), .A2(G2067), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n995), .B2(new_n997), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n992), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT63), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G305), .A2(G1981), .ZN(new_n1009));
  INV_X1    g584(.A(G1981), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n591), .A2(new_n1010), .A3(new_n592), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT114), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1009), .A2(new_n1015), .A3(KEYINPUT49), .A4(new_n1011), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  INV_X1    g593(.A(G40), .ZN(new_n1019));
  NOR4_X1   g594(.A1(new_n465), .A2(new_n471), .A3(new_n470), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1018), .B1(new_n980), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n735), .A2(G1976), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(new_n1024), .B2(new_n1021), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT113), .B1(new_n735), .B2(G1976), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1021), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1026), .B(new_n1021), .C1(new_n1024), .C2(KEYINPUT52), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1017), .A2(new_n1023), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n907), .A2(KEYINPUT45), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1020), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n498), .B2(new_n1031), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(G1971), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n494), .B1(new_n484), .B2(new_n487), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT50), .B1(new_n1037), .B2(G1384), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n498), .A2(new_n1031), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1020), .B(new_n1038), .C1(new_n1039), .C2(KEYINPUT50), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(G2090), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G303), .A2(G8), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT55), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n983), .B1(new_n980), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1036), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n1044), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1030), .A2(new_n1045), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n1031), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n907), .A2(new_n1031), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n983), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n498), .A2(KEYINPUT115), .A3(KEYINPUT45), .A4(new_n1031), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1020), .B1(new_n1058), .B2(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1047), .B1(new_n498), .B2(new_n1031), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2084), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n763), .A2(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1067), .A2(new_n1018), .A3(G286), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1008), .B1(new_n1054), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1008), .B1(new_n1051), .B2(new_n1044), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1030), .A2(new_n1053), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1017), .A2(new_n1023), .ZN(new_n1074));
  OR2_X1    g649(.A1(G288), .A2(G1976), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1011), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1076), .A2(new_n1021), .B1(new_n1052), .B2(new_n1030), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(G2078), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1020), .B(new_n1081), .C1(new_n980), .C2(KEYINPUT45), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1032), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1039), .A2(new_n1059), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n983), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n781), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1084), .B1(new_n1087), .B2(new_n1080), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n1049), .B2(new_n814), .ZN(new_n1090));
  AOI211_X1 g665(.A(KEYINPUT121), .B(G1961), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1088), .B(G301), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT122), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n814), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT121), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1049), .A2(new_n1089), .A3(new_n814), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(G301), .A4(new_n1088), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .A4(new_n1081), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1094), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT120), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1094), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1087), .A2(new_n1080), .ZN(new_n1107));
  AOI21_X1  g682(.A(G301), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1079), .B1(new_n1100), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G168), .A2(new_n1018), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT51), .B1(new_n1112), .B2(KEYINPUT119), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1062), .A2(new_n763), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(G8), .B(new_n1114), .C1(new_n1117), .C2(G286), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1112), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1119), .B(new_n1113), .C1(new_n1067), .C2(new_n1018), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1118), .A2(new_n1120), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n612), .A2(KEYINPUT60), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT117), .B1(new_n1058), .B2(new_n983), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n980), .A2(new_n1020), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n831), .A3(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1122), .B(new_n1126), .C1(new_n1065), .C2(G1348), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT58), .B(G1341), .Z(new_n1128));
  AND3_X1   g703(.A1(new_n980), .A2(new_n1020), .A3(new_n1124), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1124), .B1(new_n980), .B2(new_n1020), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1085), .A2(new_n714), .A3(new_n1086), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n552), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1127), .B1(new_n1133), .B2(KEYINPUT59), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  AOI211_X1 g710(.A(new_n1135), .B(new_n552), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT56), .B(G2072), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT116), .B(G1956), .Z(new_n1140));
  AOI22_X1  g715(.A1(new_n1035), .A2(new_n1139), .B1(new_n1040), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n566), .A2(new_n567), .B1(G91), .B2(new_n549), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT57), .B1(new_n572), .B2(new_n574), .ZN(new_n1143));
  AOI22_X1  g718(.A1(G299), .A2(KEYINPUT57), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1138), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n576), .A2(new_n575), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT75), .B1(new_n563), .B2(G651), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n565), .B(new_n505), .C1(new_n561), .C2(new_n562), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n569), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT57), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n498), .A2(new_n1047), .A3(new_n1031), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1020), .B1(new_n980), .B2(new_n1047), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1140), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1085), .A2(new_n1086), .A3(new_n1139), .ZN(new_n1155));
  AOI221_X4 g730(.A(KEYINPUT118), .B1(new_n1150), .B2(new_n1151), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1145), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1144), .B1(new_n1155), .B2(new_n1154), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1138), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1049), .A2(new_n816), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1165), .A2(new_n612), .A3(new_n1126), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n612), .B1(new_n1165), .B2(new_n1126), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT60), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1137), .A2(new_n1161), .A3(new_n1164), .A4(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1170), .A2(new_n1167), .B1(new_n1159), .B2(new_n1158), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1121), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1106), .A2(G301), .A3(new_n1107), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT124), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1097), .A2(new_n1088), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1097), .A2(KEYINPUT125), .A3(new_n1088), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(G171), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1106), .A2(new_n1180), .A3(G301), .A4(new_n1107), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1174), .A2(new_n1179), .A3(KEYINPUT54), .A4(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(KEYINPUT123), .B(new_n1079), .C1(new_n1100), .C2(new_n1108), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1111), .A2(new_n1172), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1121), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1121), .A2(new_n1185), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1186), .A2(new_n1187), .A3(new_n1108), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1054), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1078), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AND2_X1   g766(.A1(G290), .A2(G1986), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1001), .B1(new_n984), .B2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT111), .Z(new_n1194));
  NAND2_X1  g769(.A1(new_n999), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1007), .B1(new_n1191), .B2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g771(.A1(new_n694), .A2(new_n696), .A3(new_n456), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1198), .A2(KEYINPUT127), .ZN(new_n1199));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n1200));
  NAND4_X1  g774(.A1(new_n694), .A2(new_n696), .A3(new_n1200), .A4(new_n456), .ZN(new_n1201));
  NAND3_X1  g775(.A1(new_n672), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  NOR3_X1   g776(.A1(new_n1202), .A2(new_n725), .A3(new_n726), .ZN(new_n1203));
  OAI211_X1 g777(.A(new_n929), .B(new_n1203), .C1(new_n972), .C2(new_n973), .ZN(G225));
  INV_X1    g778(.A(G225), .ZN(G308));
endmodule


