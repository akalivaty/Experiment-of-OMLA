

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U324 ( .A(n397), .B(n396), .ZN(n541) );
  NOR2_X1 U325 ( .A1(n482), .A2(n581), .ZN(n483) );
  XNOR2_X1 U326 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U327 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n292) );
  XOR2_X1 U328 ( .A(n440), .B(KEYINPUT20), .Z(n293) );
  XOR2_X1 U329 ( .A(KEYINPUT40), .B(n493), .Z(n294) );
  XOR2_X1 U330 ( .A(G71GAT), .B(G120GAT), .Z(n295) );
  XOR2_X1 U331 ( .A(n342), .B(n341), .Z(n296) );
  XOR2_X1 U332 ( .A(n465), .B(KEYINPUT25), .Z(n297) );
  NOR2_X1 U333 ( .A1(n539), .A2(n466), .ZN(n467) );
  INV_X1 U334 ( .A(KEYINPUT55), .ZN(n438) );
  XNOR2_X1 U335 ( .A(n442), .B(n292), .ZN(n443) );
  XNOR2_X1 U336 ( .A(n343), .B(n296), .ZN(n344) );
  XNOR2_X1 U337 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U338 ( .A(n345), .B(n344), .ZN(n350) );
  INV_X1 U339 ( .A(G183GAT), .ZN(n453) );
  XNOR2_X1 U340 ( .A(n450), .B(n449), .ZN(n513) );
  XNOR2_X1 U341 ( .A(n453), .B(KEYINPUT124), .ZN(n454) );
  XNOR2_X1 U342 ( .A(n455), .B(n454), .ZN(G1350GAT) );
  XNOR2_X1 U343 ( .A(G183GAT), .B(G71GAT), .ZN(n298) );
  XNOR2_X1 U344 ( .A(G8GAT), .B(G1GAT), .ZN(n354) );
  XNOR2_X1 U345 ( .A(n298), .B(n354), .ZN(n311) );
  XOR2_X1 U346 ( .A(G57GAT), .B(KEYINPUT13), .Z(n372) );
  XOR2_X1 U347 ( .A(G22GAT), .B(G155GAT), .Z(n314) );
  XOR2_X1 U348 ( .A(n372), .B(n314), .Z(n300) );
  NAND2_X1 U349 ( .A1(G231GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U351 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n302) );
  XNOR2_X1 U352 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U354 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U355 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XOR2_X1 U356 ( .A(KEYINPUT82), .B(G64GAT), .Z(n306) );
  XNOR2_X1 U357 ( .A(G78GAT), .B(G211GAT), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n442), .B(n307), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n529) );
  XOR2_X1 U362 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n313) );
  XNOR2_X1 U363 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n318) );
  XOR2_X1 U365 ( .A(KEYINPUT22), .B(G218GAT), .Z(n316) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G162GAT), .Z(n332) );
  XNOR2_X1 U367 ( .A(n332), .B(n314), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U369 ( .A(n318), .B(n317), .Z(n320) );
  NAND2_X1 U370 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n322) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n321), .B(KEYINPUT2), .ZN(n419) );
  XOR2_X1 U374 ( .A(n322), .B(n419), .Z(n330) );
  XNOR2_X1 U375 ( .A(G148GAT), .B(KEYINPUT73), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n323), .B(KEYINPUT74), .ZN(n324) );
  XOR2_X1 U377 ( .A(n324), .B(G204GAT), .Z(n326) );
  XNOR2_X1 U378 ( .A(G78GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n376) );
  XOR2_X1 U380 ( .A(G211GAT), .B(KEYINPUT21), .Z(n328) );
  XNOR2_X1 U381 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n405) );
  XNOR2_X1 U383 ( .A(n376), .B(n405), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n464) );
  XOR2_X1 U385 ( .A(G43GAT), .B(G134GAT), .Z(n447) );
  XOR2_X1 U386 ( .A(G36GAT), .B(G218GAT), .Z(n402) );
  AND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n402), .B(n331), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n447), .B(n334), .ZN(n345) );
  XOR2_X1 U391 ( .A(G92GAT), .B(KEYINPUT80), .Z(n336) );
  XNOR2_X1 U392 ( .A(KEYINPUT79), .B(KEYINPUT11), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U394 ( .A(KEYINPUT81), .B(G106GAT), .Z(n338) );
  XNOR2_X1 U395 ( .A(G190GAT), .B(G99GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U397 ( .A(n340), .B(n339), .Z(n343) );
  XOR2_X1 U398 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n342) );
  XNOR2_X1 U399 ( .A(KEYINPUT9), .B(KEYINPUT66), .ZN(n341) );
  XOR2_X1 U400 ( .A(G29GAT), .B(KEYINPUT7), .Z(n347) );
  XNOR2_X1 U401 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n358) );
  XNOR2_X1 U403 ( .A(G85GAT), .B(KEYINPUT75), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n348), .B(KEYINPUT76), .ZN(n381) );
  XNOR2_X1 U405 ( .A(n358), .B(n381), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n551) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G113GAT), .Z(n352) );
  XNOR2_X1 U408 ( .A(G50GAT), .B(G36GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U410 ( .A(n353), .B(G43GAT), .Z(n357) );
  INV_X1 U411 ( .A(n354), .ZN(n355) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(n355), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U414 ( .A(n358), .B(KEYINPUT67), .Z(n360) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U417 ( .A(n362), .B(n361), .Z(n370) );
  XOR2_X1 U418 ( .A(KEYINPUT71), .B(G22GAT), .Z(n364) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(G141GAT), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U421 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n366) );
  XNOR2_X1 U422 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n571) );
  XNOR2_X1 U426 ( .A(G92GAT), .B(G64GAT), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n371), .B(KEYINPUT77), .ZN(n403) );
  XOR2_X1 U428 ( .A(n403), .B(KEYINPUT78), .Z(n374) );
  XNOR2_X1 U429 ( .A(n372), .B(KEYINPUT33), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n385) );
  XOR2_X1 U432 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n378) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U435 ( .A(n379), .B(KEYINPUT32), .Z(n383) );
  XNOR2_X1 U436 ( .A(G99GAT), .B(G176GAT), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n295), .B(n380), .ZN(n440) );
  XNOR2_X1 U438 ( .A(n440), .B(n381), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n577) );
  XNOR2_X1 U441 ( .A(KEYINPUT41), .B(n577), .ZN(n547) );
  NAND2_X1 U442 ( .A1(n571), .A2(n547), .ZN(n386) );
  XNOR2_X1 U443 ( .A(KEYINPUT46), .B(n386), .ZN(n387) );
  NAND2_X1 U444 ( .A1(n387), .A2(n529), .ZN(n388) );
  NOR2_X1 U445 ( .A1(n551), .A2(n388), .ZN(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT109), .B(KEYINPUT47), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n395) );
  INV_X1 U448 ( .A(n529), .ZN(n581) );
  XNOR2_X1 U449 ( .A(n551), .B(KEYINPUT36), .ZN(n584) );
  NAND2_X1 U450 ( .A1(n581), .A2(n584), .ZN(n391) );
  XOR2_X1 U451 ( .A(KEYINPUT45), .B(n391), .Z(n392) );
  NAND2_X1 U452 ( .A1(n577), .A2(n392), .ZN(n393) );
  NOR2_X1 U453 ( .A1(n571), .A2(n393), .ZN(n394) );
  NOR2_X1 U454 ( .A1(n395), .A2(n394), .ZN(n397) );
  XNOR2_X1 U455 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n398), .B(KEYINPUT19), .ZN(n399) );
  XOR2_X1 U457 ( .A(n399), .B(KEYINPUT17), .Z(n401) );
  XNOR2_X1 U458 ( .A(G169GAT), .B(G190GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n448) );
  XNOR2_X1 U460 ( .A(G204GAT), .B(n402), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n409) );
  XOR2_X1 U462 ( .A(KEYINPUT94), .B(n405), .Z(n407) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U465 ( .A(n409), .B(n408), .Z(n414) );
  XOR2_X1 U466 ( .A(KEYINPUT96), .B(KEYINPUT93), .Z(n411) );
  XNOR2_X1 U467 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(G176GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n448), .B(n415), .ZN(n490) );
  NOR2_X1 U472 ( .A1(n541), .A2(n490), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n416), .B(KEYINPUT54), .ZN(n437) );
  XOR2_X1 U474 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n418) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n423) );
  XOR2_X1 U477 ( .A(G162GAT), .B(n419), .Z(n421) );
  XOR2_X1 U478 ( .A(G113GAT), .B(KEYINPUT0), .Z(n445) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(n445), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n436) );
  XOR2_X1 U482 ( .A(G85GAT), .B(KEYINPUT81), .Z(n425) );
  XNOR2_X1 U483 ( .A(G134GAT), .B(G120GAT), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U485 ( .A(G57GAT), .B(G155GAT), .Z(n427) );
  XNOR2_X1 U486 ( .A(G127GAT), .B(G148GAT), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U488 ( .A(n429), .B(n428), .Z(n434) );
  XOR2_X1 U489 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n431) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U492 ( .A(KEYINPUT92), .B(n432), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n487) );
  NAND2_X1 U495 ( .A1(n437), .A2(n487), .ZN(n569) );
  NOR2_X1 U496 ( .A1(n464), .A2(n569), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n451) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n293), .B(n441), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U501 ( .A(n448), .B(n447), .Z(n449) );
  NAND2_X1 U502 ( .A1(n451), .A2(n513), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n452), .B(KEYINPUT120), .ZN(n565) );
  NOR2_X1 U504 ( .A1(n529), .A2(n565), .ZN(n455) );
  XOR2_X1 U505 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n473) );
  NAND2_X1 U506 ( .A1(n571), .A2(n577), .ZN(n484) );
  XOR2_X1 U507 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n457) );
  INV_X1 U508 ( .A(n551), .ZN(n564) );
  NAND2_X1 U509 ( .A1(n581), .A2(n564), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(n471) );
  XNOR2_X1 U511 ( .A(KEYINPUT87), .B(n513), .ZN(n459) );
  XNOR2_X1 U512 ( .A(KEYINPUT27), .B(n490), .ZN(n462) );
  OR2_X1 U513 ( .A1(n487), .A2(n462), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n464), .B(KEYINPUT28), .ZN(n515) );
  NOR2_X1 U515 ( .A1(n458), .A2(n515), .ZN(n522) );
  NAND2_X1 U516 ( .A1(n459), .A2(n522), .ZN(n470) );
  XOR2_X1 U517 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n461) );
  INV_X1 U518 ( .A(n513), .ZN(n520) );
  NAND2_X1 U519 ( .A1(n464), .A2(n520), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(n570) );
  NOR2_X1 U521 ( .A1(n570), .A2(n462), .ZN(n539) );
  NOR2_X1 U522 ( .A1(n520), .A2(n490), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U524 ( .A(KEYINPUT98), .B(n297), .ZN(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT99), .B(n467), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n468), .A2(n487), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n481) );
  NAND2_X1 U528 ( .A1(n471), .A2(n481), .ZN(n497) );
  NOR2_X1 U529 ( .A1(n484), .A2(n497), .ZN(n479) );
  INV_X1 U530 ( .A(n487), .ZN(n538) );
  NAND2_X1 U531 ( .A1(n479), .A2(n538), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n474), .Z(G1324GAT) );
  INV_X1 U534 ( .A(n490), .ZN(n511) );
  NAND2_X1 U535 ( .A1(n479), .A2(n511), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n475), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U538 ( .A1(n479), .A2(n513), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U540 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NAND2_X1 U541 ( .A1(n515), .A2(n479), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n480), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U543 ( .A1(n584), .A2(n481), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(KEYINPUT37), .ZN(n509) );
  NOR2_X1 U545 ( .A1(n509), .A2(n484), .ZN(n486) );
  XOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n494) );
  NOR2_X1 U548 ( .A1(n487), .A2(n494), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n490), .A2(n494), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1329GAT) );
  NOR2_X1 U554 ( .A1(n520), .A2(n494), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n294), .ZN(G1330GAT) );
  INV_X1 U556 ( .A(n515), .ZN(n495) );
  NOR2_X1 U557 ( .A1(n495), .A2(n494), .ZN(n496) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n499) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(n547), .Z(n558) );
  OR2_X1 U561 ( .A1(n558), .A2(n571), .ZN(n508) );
  NOR2_X1 U562 ( .A1(n508), .A2(n497), .ZN(n504) );
  NAND2_X1 U563 ( .A1(n504), .A2(n538), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(G1332GAT) );
  XOR2_X1 U565 ( .A(G64GAT), .B(KEYINPUT105), .Z(n501) );
  NAND2_X1 U566 ( .A1(n504), .A2(n511), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n504), .A2(n513), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n502), .B(KEYINPUT106), .ZN(n503) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n503), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n515), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n507), .Z(G1335GAT) );
  NOR2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n538), .A2(n516), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n511), .A2(n516), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(n512), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n518) );
  NAND2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U585 ( .A(G106GAT), .B(n519), .Z(G1339GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n541), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT110), .B(n523), .ZN(n533) );
  INV_X1 U589 ( .A(n571), .ZN(n555) );
  NOR2_X1 U590 ( .A1(n533), .A2(n555), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1340GAT) );
  NOR2_X1 U593 ( .A1(n533), .A2(n558), .ZN(n527) );
  XNOR2_X1 U594 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(n528), .ZN(G1341GAT) );
  XNOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT113), .ZN(n531) );
  NOR2_X1 U598 ( .A1(n529), .A2(n533), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  NOR2_X1 U601 ( .A1(n564), .A2(n533), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n535) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n552), .A2(n571), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(KEYINPUT116), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n545) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U614 ( .A(KEYINPUT52), .B(n546), .Z(n549) );
  NAND2_X1 U615 ( .A1(n552), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n581), .A2(n552), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT119), .Z(n554) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1347GAT) );
  NOR2_X1 U622 ( .A1(n565), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  NOR2_X1 U625 ( .A1(n565), .A2(n558), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n560) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(KEYINPUT56), .B(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n568), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n583) );
  NAND2_X1 U637 ( .A1(n583), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(n574), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U643 ( .A(n577), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n583), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

