//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n438, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(new_n438));
  INV_X1    g013(.A(new_n438), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(new_n438), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n458));
  AND3_X1   g033(.A1(new_n454), .A2(new_n458), .A3(G2106), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n458), .B1(new_n454), .B2(G2106), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n455), .A2(G567), .ZN(new_n461));
  NOR3_X1   g036(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n467), .A2(new_n473), .A3(new_n470), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n464), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n463), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n478), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n472), .A2(new_n480), .A3(KEYINPUT70), .A4(new_n474), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(KEYINPUT71), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g060(.A1(KEYINPUT71), .A2(G100), .A3(G2105), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G112), .B2(new_n464), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n487), .B(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n464), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n493));
  AOI22_X1  g068(.A1(G124), .A2(new_n492), .B1(new_n493), .B2(G136), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT73), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n489), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n496), .A2(new_n498), .ZN(G162));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(new_n503), .A3(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(G138), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n490), .A2(new_n491), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G138), .A4(new_n464), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n505), .B1(new_n507), .B2(new_n510), .ZN(G164));
  NAND2_X1  g086(.A1(KEYINPUT74), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(KEYINPUT74), .A2(KEYINPUT6), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(G88), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n514), .B2(new_n515), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  OAI21_X1  g099(.A(G62), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n518), .B(new_n521), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n532));
  AND3_X1   g107(.A1(KEYINPUT74), .A2(KEYINPUT6), .A3(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT6), .B1(KEYINPUT74), .B2(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(G543), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT76), .B(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n532), .B(KEYINPUT77), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n533), .A2(new_n534), .B1(new_n523), .B2(new_n524), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n542), .A2(G89), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n539), .A2(new_n540), .A3(new_n546), .ZN(G168));
  NAND2_X1  g122(.A1(new_n520), .A2(G52), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n516), .A2(G90), .A3(new_n517), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n522), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n523), .A2(new_n524), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n542), .A2(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n520), .A2(G43), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n567));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n541), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT80), .A4(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n554), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n569), .A2(new_n570), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n535), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n520), .A2(G53), .A3(new_n575), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n580), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n574), .B1(new_n581), .B2(new_n582), .ZN(G299));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n551), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G77), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G64), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n554), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n589), .A2(KEYINPUT81), .A3(new_n548), .A4(new_n549), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G301));
  NAND3_X1  g167(.A1(new_n539), .A2(new_n540), .A3(new_n546), .ZN(G286));
  INV_X1    g168(.A(G166), .ZN(G303));
  NAND2_X1  g169(.A1(new_n520), .A2(G49), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n596));
  INV_X1    g171(.A(G87), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n541), .ZN(G288));
  NAND3_X1  g173(.A1(new_n516), .A2(G86), .A3(new_n517), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT82), .A4(G86), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G61), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n554), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G48), .B2(new_n520), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(G72), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G60), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n554), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G651), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT83), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n611), .A2(new_n614), .A3(G651), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT84), .B(G47), .Z(new_n616));
  AOI22_X1  g191(.A1(new_n542), .A2(G85), .B1(new_n520), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n613), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT85), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n613), .A2(new_n620), .A3(new_n617), .A4(new_n615), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(G290));
  NAND2_X1  g197(.A1(new_n520), .A2(G54), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n522), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n541), .B2(new_n627), .ZN(new_n628));
  NOR3_X1   g203(.A1(new_n541), .A2(new_n626), .A3(new_n627), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  MUX2_X1   g207(.A(new_n632), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g208(.A(new_n632), .B(G301), .S(G868), .Z(G321));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(G299), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(G168), .ZN(G297));
  OAI21_X1  g212(.A(new_n636), .B1(new_n635), .B2(G168), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n631), .B1(new_n639), .B2(G860), .ZN(G148));
  OR3_X1    g215(.A1(new_n632), .A2(KEYINPUT86), .A3(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(KEYINPUT86), .B1(new_n632), .B2(G559), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  MUX2_X1   g218(.A(new_n560), .B(new_n643), .S(G868), .Z(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n493), .A2(G135), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT89), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n492), .A2(G123), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n464), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT90), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n653), .A2(G2096), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(G2096), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n508), .A2(new_n469), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT13), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT88), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(new_n655), .A3(new_n661), .ZN(G156));
  INV_X1    g237(.A(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2427), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2430), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT15), .B(G2435), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  XOR2_X1   g245(.A(G1341), .B(G1348), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n668), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2443), .B(G2446), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(G14), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(G401));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n679));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(KEYINPUT17), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n682), .B2(KEYINPUT18), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT91), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n685), .B(new_n686), .ZN(new_n692));
  INV_X1    g267(.A(new_n690), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(G227));
  XOR2_X1   g270(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1956), .B(G2474), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1961), .B(G1966), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(KEYINPUT93), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n699), .A2(new_n700), .A3(KEYINPUT93), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n698), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT20), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(new_n707), .B(new_n706), .S(new_n698), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT94), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n714));
  XOR2_X1   g289(.A(new_n713), .B(new_n714), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n710), .A2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(G229));
  MUX2_X1   g294(.A(G23), .B(G288), .S(G16), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT33), .ZN(new_n721));
  INV_X1    g296(.A(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G6), .ZN(new_n725));
  INV_X1    g300(.A(G305), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT32), .B(G1981), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n724), .A2(G22), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G166), .B2(new_n724), .ZN(new_n731));
  INV_X1    g306(.A(G1971), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  OR3_X1    g309(.A1(new_n723), .A2(KEYINPUT34), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT34), .B1(new_n723), .B2(new_n734), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n724), .A2(G24), .ZN(new_n737));
  INV_X1    g312(.A(G290), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n724), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n739), .A2(G1986), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G25), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n493), .A2(G131), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n745));
  INV_X1    g320(.A(G107), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G2105), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G119), .B2(new_n492), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n742), .B1(new_n750), .B2(new_n741), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT35), .B(G1991), .Z(new_n752));
  XOR2_X1   g327(.A(new_n751), .B(new_n752), .Z(new_n753));
  NOR2_X1   g328(.A1(new_n739), .A2(G1986), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n740), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n735), .A2(new_n736), .A3(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT36), .Z(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G35), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G162), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT29), .ZN(new_n760));
  INV_X1    g335(.A(G2090), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n493), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n492), .A2(G128), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n464), .A2(G116), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n741), .A2(G26), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT28), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2067), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  NOR2_X1   g348(.A1(G171), .A2(new_n724), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G5), .B2(new_n724), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2078), .ZN(new_n777));
  NAND2_X1  g352(.A1(G164), .A2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G27), .B2(G29), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n776), .B1(new_n777), .B2(new_n779), .C1(new_n653), .C2(new_n741), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n724), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n561), .B2(new_n724), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1341), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n631), .A2(G16), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G4), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n783), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n775), .A2(new_n773), .ZN(new_n790));
  NOR2_X1   g365(.A1(G29), .A2(G33), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT96), .Z(new_n792));
  AND2_X1   g367(.A1(new_n508), .A2(G127), .ZN(new_n793));
  AND2_X1   g368(.A1(G115), .A2(G2104), .ZN(new_n794));
  OAI21_X1  g369(.A(G2105), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n796));
  NAND2_X1  g371(.A1(G103), .A2(G2104), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n493), .A2(G139), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(new_n741), .ZN(new_n802));
  INV_X1    g377(.A(G2072), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT99), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n806), .A2(new_n805), .A3(G28), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n805), .B2(G28), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n741), .B1(new_n805), .B2(G28), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G11), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n802), .B2(new_n803), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n779), .A2(new_n777), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n790), .A2(new_n804), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n780), .A2(new_n789), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G34), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(KEYINPUT24), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(KEYINPUT24), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n741), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G160), .B2(new_n741), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G2084), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n741), .A2(G32), .ZN(new_n822));
  NAND3_X1  g397(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT26), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n492), .A2(G129), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n493), .A2(G141), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n469), .A2(G105), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT97), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n822), .B1(new_n835), .B2(new_n741), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT27), .B(G1996), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT98), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n724), .A2(G20), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT23), .Z(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G299), .B2(G16), .ZN(new_n842));
  INV_X1    g417(.A(G1956), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n724), .A2(G21), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G168), .B2(new_n724), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G1966), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n839), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n762), .A2(new_n815), .A3(new_n821), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n757), .A2(new_n849), .ZN(G311));
  OR2_X1    g425(.A1(new_n757), .A2(new_n849), .ZN(G150));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  INV_X1    g427(.A(G67), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n554), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G651), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n542), .A2(G93), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n520), .A2(G55), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n631), .A2(G559), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(G651), .A2(new_n556), .B1(new_n542), .B2(G81), .ZN(new_n864));
  AOI22_X1  g439(.A1(G651), .A2(new_n854), .B1(new_n542), .B2(G93), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n559), .A4(new_n857), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n560), .A2(new_n858), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n863), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT101), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(G860), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n860), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT102), .Z(G145));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n878), .A2(new_n464), .A3(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n464), .B2(G118), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n879), .A2(G2104), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n492), .A2(G130), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n493), .A2(G142), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n744), .B2(new_n748), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n744), .A2(new_n748), .A3(new_n885), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n658), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(new_n658), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n890), .A2(new_n891), .A3(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n877), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n890), .B2(new_n886), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(new_n658), .A3(new_n888), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT105), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n801), .B1(new_n832), .B2(new_n834), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n500), .A2(new_n504), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n509), .B1(new_n493), .B2(G138), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n767), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n801), .A2(new_n830), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n898), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n903), .B1(new_n898), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n893), .A2(new_n906), .A3(new_n907), .A4(new_n896), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n482), .A2(KEYINPUT103), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n482), .A2(KEYINPUT103), .ZN(new_n914));
  OAI21_X1  g489(.A(G162), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n482), .A2(KEYINPUT103), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n496), .A2(new_n498), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n912), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n652), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n652), .B1(new_n915), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n911), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n889), .A2(new_n892), .ZN(new_n923));
  OAI221_X1 g498(.A(new_n909), .B1(new_n908), .B2(new_n923), .C1(new_n919), .C2(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g501(.A(new_n643), .B(new_n868), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n632), .A2(G299), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n578), .A2(new_n579), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT79), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n631), .A3(new_n574), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n928), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n928), .B2(new_n934), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n927), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n928), .A2(new_n934), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n927), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(G290), .A2(new_n726), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n619), .A2(G305), .A3(new_n621), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(G166), .B(G288), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n949), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n946), .A3(new_n947), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n943), .B2(KEYINPUT42), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n939), .B(new_n941), .C1(new_n943), .C2(KEYINPUT42), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n945), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n945), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g532(.A(G868), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n858), .A2(new_n635), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(G295));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n959), .ZN(G331));
  INV_X1    g536(.A(new_n868), .ZN(new_n962));
  NAND2_X1  g537(.A1(G286), .A2(new_n551), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G286), .B1(new_n585), .B2(new_n590), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n591), .A2(G168), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n868), .A3(new_n963), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n966), .B(new_n968), .C1(new_n935), .C2(new_n937), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n967), .A2(new_n868), .A3(new_n963), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n868), .B1(new_n967), .B2(new_n963), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n940), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n972), .A3(KEYINPUT108), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n970), .A2(new_n971), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n974), .B(new_n975), .C1(new_n937), .C2(new_n935), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n953), .ZN(new_n978));
  INV_X1    g553(.A(G37), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n950), .A2(new_n952), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n973), .A2(new_n980), .A3(new_n976), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n973), .B2(new_n976), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n928), .A2(new_n934), .A3(KEYINPUT109), .A4(new_n936), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n966), .A2(new_n985), .A3(new_n968), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n928), .A2(new_n934), .A3(new_n936), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n987), .B(new_n988), .C1(new_n940), .C2(new_n929), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n953), .B1(new_n990), .B2(new_n972), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  NOR4_X1   g567(.A1(new_n984), .A2(new_n991), .A3(new_n992), .A4(G37), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT44), .B1(new_n983), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n977), .B2(new_n953), .ZN(new_n995));
  INV_X1    g570(.A(new_n991), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n992), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n982), .B2(new_n992), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n994), .B1(KEYINPUT44), .B2(new_n999), .ZN(G397));
  XNOR2_X1  g575(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(G164), .B2(G1384), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n472), .A2(new_n480), .A3(G40), .A4(new_n474), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n835), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G2067), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n767), .B(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1006), .B(new_n1008), .C1(new_n1005), .C2(new_n830), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n749), .B(new_n752), .Z(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1986), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n738), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n738), .A2(new_n1012), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1004), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(G166), .B2(new_n1017), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT55), .B(G8), .C1(new_n529), .C2(new_n530), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n902), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n467), .A2(new_n473), .A3(new_n470), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n473), .B1(new_n467), .B2(new_n470), .ZN(new_n1024));
  INV_X1    g599(.A(G40), .ZN(new_n1025));
  NOR4_X1   g600(.A1(new_n1023), .A2(new_n1024), .A3(new_n478), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1002), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n732), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n902), .A2(new_n1029), .A3(new_n1021), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1026), .A4(new_n761), .ZN(new_n1032));
  AOI221_X4 g607(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .C1(new_n1028), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n722), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(KEYINPUT111), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n1037), .B(KEYINPUT52), .C1(G288), .C2(new_n722), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n542), .A2(G87), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1040), .A2(G1976), .A3(new_n595), .A4(new_n596), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n902), .A2(new_n1021), .ZN(new_n1042));
  OAI211_X1 g617(.A(G8), .B(new_n1041), .C1(new_n1042), .C2(new_n1003), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1981), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n603), .A2(new_n607), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n520), .A2(G48), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1051), .B(new_n599), .C1(new_n1052), .C2(new_n522), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G1981), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1048), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G164), .A2(G1384), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1017), .B1(new_n1026), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(new_n1054), .A3(new_n1048), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1045), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G288), .A2(G1976), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1060), .A2(new_n1063), .B1(new_n1049), .B2(new_n726), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1058), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1034), .A2(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n1067));
  INV_X1    g642(.A(G1966), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT45), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(G164), .B2(G1384), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1026), .A3(new_n1071), .ZN(new_n1072));
  OR3_X1    g647(.A1(G164), .A2(G1384), .A3(new_n1001), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1070), .B2(new_n1026), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1068), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1031), .A2(new_n1030), .A3(new_n1026), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT116), .B(G2084), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1017), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT117), .B1(new_n1081), .B2(G168), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT45), .B1(new_n902), .B2(new_n1021), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT115), .B1(new_n1083), .B2(new_n1003), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n1073), .A3(new_n1072), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1085), .A2(new_n1068), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  NOR4_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1017), .A4(G286), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1082), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1061), .B1(new_n1090), .B2(new_n1055), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1043), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT114), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1045), .A2(new_n1060), .A3(new_n1094), .A4(new_n1061), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1033), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1078), .A2(new_n761), .B1(new_n1027), .B2(new_n732), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT113), .B(new_n1098), .C1(new_n1099), .C2(new_n1017), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1017), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1097), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1067), .B1(new_n1089), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1102), .A2(new_n1097), .ZN(new_n1107));
  NOR4_X1   g682(.A1(new_n1107), .A2(new_n1033), .A3(new_n1062), .A4(new_n1067), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1088), .B2(new_n1082), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1066), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1077), .A2(new_n843), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n578), .B2(new_n579), .ZN(new_n1112));
  AOI22_X1  g687(.A1(G299), .A2(KEYINPUT57), .B1(new_n574), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1002), .A2(new_n1022), .A3(new_n1026), .A4(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1042), .A2(new_n1003), .A3(G2067), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n786), .B2(new_n1077), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(new_n632), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1113), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(new_n1120), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1003), .B1(new_n1042), .B2(KEYINPUT50), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n1126), .B2(new_n1030), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1127), .B2(new_n1117), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1118), .A2(KEYINPUT60), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n631), .ZN(new_n1130));
  NAND2_X1  g705(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n574), .A2(new_n1112), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1956), .B1(new_n1126), .B2(new_n1030), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1115), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n1116), .A3(KEYINPUT61), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1124), .A2(new_n1130), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1042), .A2(new_n1003), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT58), .B(G1341), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1027), .A2(G1996), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n561), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(KEYINPUT59), .A3(new_n561), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1144), .B(new_n1145), .C1(new_n631), .C2(new_n1129), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1121), .B1(new_n1138), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G168), .A2(new_n1017), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT119), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1150), .B1(new_n1081), .B2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(KEYINPUT120), .B(new_n1152), .C1(new_n1086), .C2(new_n1017), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(KEYINPUT51), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1086), .A2(new_n1152), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT51), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1150), .B(new_n1158), .C1(new_n1081), .C2(new_n1153), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1002), .A2(new_n1022), .A3(new_n1026), .A4(new_n777), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1162), .A2(new_n1163), .B1(new_n1077), .B2(new_n773), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(G2078), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n480), .A2(G40), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n475), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n472), .A2(KEYINPUT121), .A3(new_n474), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1168), .A2(new_n1002), .A3(new_n1022), .A4(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1164), .A2(KEYINPUT122), .A3(G301), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1077), .A2(new_n773), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(G301), .A3(new_n1173), .A4(new_n1170), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1084), .A2(new_n1073), .A3(new_n1072), .A4(new_n1165), .ZN(new_n1177));
  AOI21_X1  g752(.A(G301), .B1(new_n1164), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1161), .B(new_n1171), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1164), .A2(G301), .A3(new_n1177), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1181));
  OAI211_X1 g756(.A(KEYINPUT54), .B(new_n1180), .C1(new_n1181), .C2(new_n551), .ZN(new_n1182));
  AND4_X1   g757(.A1(new_n1104), .A2(new_n1179), .A3(new_n1096), .A4(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(KEYINPUT118), .B(new_n1121), .C1(new_n1138), .C2(new_n1146), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1149), .A2(new_n1160), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1110), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1096), .A2(new_n1104), .A3(new_n1178), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1160), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1156), .A2(KEYINPUT62), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1016), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1008), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1004), .B1(new_n1193), .B2(new_n831), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1004), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1195), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT46), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1194), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT47), .Z(new_n1200));
  XNOR2_X1  g775(.A(KEYINPUT124), .B(KEYINPUT48), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(new_n1013), .B2(new_n1195), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(new_n1011), .B2(new_n1195), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1013), .A2(new_n1195), .A3(new_n1201), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n750), .A2(new_n752), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT123), .Z(new_n1207));
  OAI22_X1  g782(.A1(new_n1207), .A2(new_n1009), .B1(G2067), .B2(new_n767), .ZN(new_n1208));
  AOI211_X1 g783(.A(new_n1200), .B(new_n1205), .C1(new_n1004), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1192), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n1212));
  AND3_X1   g786(.A1(G319), .A2(new_n691), .A3(new_n694), .ZN(new_n1213));
  OAI21_X1  g787(.A(new_n1213), .B1(new_n676), .B2(new_n677), .ZN(new_n1214));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g790(.A(new_n1213), .B(KEYINPUT125), .C1(new_n676), .C2(new_n677), .ZN(new_n1217));
  NAND4_X1  g791(.A1(new_n1216), .A2(new_n717), .A3(new_n718), .A4(new_n1217), .ZN(new_n1218));
  AOI21_X1  g792(.A(new_n1218), .B1(new_n922), .B2(new_n924), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1212), .B1(new_n998), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n992), .B1(new_n995), .B2(new_n981), .ZN(new_n1221));
  NOR4_X1   g795(.A1(new_n984), .A2(new_n991), .A3(KEYINPUT43), .A4(G37), .ZN(new_n1222));
  OAI211_X1 g796(.A(new_n1219), .B(new_n1212), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  INV_X1    g797(.A(new_n1223), .ZN(new_n1224));
  NOR2_X1   g798(.A1(new_n1220), .A2(new_n1224), .ZN(G308));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1219), .ZN(G225));
endmodule


