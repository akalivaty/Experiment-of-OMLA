

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744;

  OR2_X1 U374 ( .A1(n743), .A2(n744), .ZN(n359) );
  INV_X1 U375 ( .A(n599), .ZN(n494) );
  XNOR2_X1 U376 ( .A(n577), .B(KEYINPUT6), .ZN(n570) );
  INV_X1 U377 ( .A(n577), .ZN(n606) );
  NAND2_X2 U378 ( .A1(n603), .A2(n602), .ZN(n599) );
  INV_X4 U379 ( .A(G953), .ZN(n735) );
  XNOR2_X1 U380 ( .A(n529), .B(n528), .ZN(n594) );
  NOR2_X1 U381 ( .A1(G953), .A2(G237), .ZN(n464) );
  AND2_X1 U382 ( .A1(n594), .A2(n593), .ZN(n640) );
  AND2_X4 U383 ( .A1(n646), .A2(n645), .ZN(n713) );
  XNOR2_X2 U384 ( .A(n432), .B(n397), .ZN(n673) );
  OR2_X1 U385 ( .A1(n644), .A2(n643), .ZN(n646) );
  BUF_X1 U386 ( .A(n640), .Z(n733) );
  AND2_X1 U387 ( .A1(n512), .A2(n361), .ZN(n360) );
  XNOR2_X1 U388 ( .A(n582), .B(n581), .ZN(n585) );
  NOR2_X1 U389 ( .A1(n382), .A2(n563), .ZN(n548) );
  AND2_X1 U390 ( .A1(n520), .A2(n494), .ZN(n495) );
  XNOR2_X1 U391 ( .A(n547), .B(KEYINPUT0), .ZN(n563) );
  INV_X2 U392 ( .A(n576), .ZN(n603) );
  XNOR2_X1 U393 ( .A(n368), .B(G146), .ZN(n444) );
  OR2_X2 U394 ( .A1(n742), .A2(KEYINPUT44), .ZN(n586) );
  XNOR2_X2 U395 ( .A(n731), .B(G146), .ZN(n432) );
  XNOR2_X2 U396 ( .A(n445), .B(n388), .ZN(n731) );
  XNOR2_X1 U397 ( .A(n444), .B(n367), .ZN(n461) );
  INV_X1 U398 ( .A(KEYINPUT10), .ZN(n367) );
  OR2_X1 U399 ( .A1(n649), .A2(n378), .ZN(n377) );
  NAND2_X1 U400 ( .A1(G234), .A2(G237), .ZN(n402) );
  XNOR2_X1 U401 ( .A(G119), .B(G128), .ZN(n414) );
  INV_X1 U402 ( .A(n429), .ZN(n418) );
  NAND2_X1 U403 ( .A1(n457), .A2(n381), .ZN(n379) );
  XNOR2_X1 U404 ( .A(n410), .B(n409), .ZN(n514) );
  INV_X1 U405 ( .A(KEYINPUT67), .ZN(n409) );
  XNOR2_X1 U406 ( .A(n473), .B(n472), .ZN(n706) );
  XNOR2_X1 U407 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U408 ( .A(n539), .B(n521), .ZN(n572) );
  INV_X1 U409 ( .A(n379), .ZN(n376) );
  XNOR2_X1 U410 ( .A(n439), .B(n438), .ZN(n520) );
  XNOR2_X1 U411 ( .A(n372), .B(KEYINPUT84), .ZN(n371) );
  XOR2_X1 U412 ( .A(G131), .B(G140), .Z(n466) );
  XNOR2_X1 U413 ( .A(n359), .B(n357), .ZN(n358) );
  AND2_X1 U414 ( .A1(n363), .A2(n362), .ZN(n361) );
  AND2_X1 U415 ( .A1(n526), .A2(n354), .ZN(n362) );
  INV_X1 U416 ( .A(G237), .ZN(n453) );
  INV_X1 U417 ( .A(KEYINPUT87), .ZN(n404) );
  INV_X1 U418 ( .A(G125), .ZN(n368) );
  XNOR2_X1 U419 ( .A(G116), .B(G101), .ZN(n393) );
  XNOR2_X1 U420 ( .A(KEYINPUT3), .B(G119), .ZN(n392) );
  INV_X1 U421 ( .A(KEYINPUT33), .ZN(n383) );
  XNOR2_X1 U422 ( .A(n419), .B(n732), .ZN(n663) );
  XNOR2_X1 U423 ( .A(n432), .B(n384), .ZN(n655) );
  XNOR2_X1 U424 ( .A(n431), .B(n437), .ZN(n384) );
  XNOR2_X1 U425 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U426 ( .A1(n735), .A2(G224), .ZN(n372) );
  NOR2_X1 U427 ( .A1(n515), .A2(n366), .ZN(n365) );
  NAND2_X1 U428 ( .A1(n351), .A2(n514), .ZN(n366) );
  AND2_X1 U429 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U430 ( .A1(n380), .A2(n355), .ZN(n534) );
  XNOR2_X1 U431 ( .A(n364), .B(n353), .ZN(n501) );
  OR2_X1 U432 ( .A1(n706), .A2(G902), .ZN(n364) );
  AND2_X1 U433 ( .A1(n501), .A2(n490), .ZN(n513) );
  XNOR2_X1 U434 ( .A(n370), .B(n564), .ZN(n579) );
  NOR2_X1 U435 ( .A1(n563), .A2(n562), .ZN(n370) );
  AND2_X1 U436 ( .A1(n377), .A2(n375), .ZN(n374) );
  NOR2_X1 U437 ( .A1(n376), .A2(n459), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n442), .B(n441), .ZN(n692) );
  AND2_X1 U439 ( .A1(n614), .A2(n576), .ZN(n351) );
  AND2_X1 U440 ( .A1(n365), .A2(n695), .ZN(n352) );
  XOR2_X1 U441 ( .A(KEYINPUT13), .B(G475), .Z(n353) );
  OR2_X1 U442 ( .A1(n619), .A2(KEYINPUT74), .ZN(n354) );
  AND2_X1 U443 ( .A1(n377), .A2(n379), .ZN(n355) );
  NOR2_X1 U444 ( .A1(n623), .A2(n382), .ZN(n356) );
  XNOR2_X1 U445 ( .A(KEYINPUT46), .B(KEYINPUT77), .ZN(n357) );
  NAND2_X1 U446 ( .A1(n360), .A2(n358), .ZN(n529) );
  XNOR2_X1 U447 ( .A(n703), .B(KEYINPUT78), .ZN(n363) );
  NAND2_X1 U448 ( .A1(n369), .A2(n574), .ZN(n575) );
  INV_X1 U449 ( .A(n579), .ZN(n369) );
  XNOR2_X1 U450 ( .A(n373), .B(n371), .ZN(n446) );
  XNOR2_X1 U451 ( .A(n444), .B(n443), .ZN(n373) );
  NAND2_X1 U452 ( .A1(n380), .A2(n374), .ZN(n460) );
  OR2_X1 U453 ( .A1(n457), .A2(n381), .ZN(n378) );
  NAND2_X1 U454 ( .A1(n649), .A2(n457), .ZN(n380) );
  INV_X1 U455 ( .A(n639), .ZN(n381) );
  NOR2_X1 U456 ( .A1(n382), .A2(n628), .ZN(n629) );
  XNOR2_X2 U457 ( .A(n541), .B(n383), .ZN(n382) );
  BUF_X1 U458 ( .A(n553), .Z(n598) );
  XNOR2_X1 U459 ( .A(n520), .B(n519), .ZN(n553) );
  NAND2_X1 U460 ( .A1(n440), .A2(n520), .ZN(n442) );
  XNOR2_X2 U461 ( .A(n477), .B(KEYINPUT4), .ZN(n445) );
  XOR2_X1 U462 ( .A(KEYINPUT75), .B(n689), .Z(n385) );
  AND2_X1 U463 ( .A1(n558), .A2(n557), .ZN(n386) );
  INV_X1 U464 ( .A(KEYINPUT71), .ZN(n433) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n542) );
  XNOR2_X1 U466 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U467 ( .A(n430), .B(G104), .ZN(n431) );
  XNOR2_X1 U468 ( .A(n527), .B(KEYINPUT66), .ZN(n528) );
  XNOR2_X1 U469 ( .A(n461), .B(n418), .ZN(n732) );
  INV_X1 U470 ( .A(KEYINPUT117), .ZN(n634) );
  INV_X1 U471 ( .A(KEYINPUT83), .ZN(n521) );
  INV_X1 U472 ( .A(KEYINPUT103), .ZN(n441) );
  XNOR2_X1 U473 ( .A(n635), .B(n634), .ZN(n636) );
  INV_X1 U474 ( .A(KEYINPUT125), .ZN(n667) );
  XNOR2_X1 U475 ( .A(n506), .B(n505), .ZN(n743) );
  XNOR2_X1 U476 ( .A(n638), .B(n637), .ZN(G75) );
  INV_X1 U477 ( .A(KEYINPUT74), .ZN(n488) );
  XNOR2_X2 U478 ( .A(G128), .B(KEYINPUT64), .ZN(n387) );
  XNOR2_X2 U479 ( .A(n387), .B(G143), .ZN(n477) );
  XNOR2_X1 U480 ( .A(G131), .B(G134), .ZN(n388) );
  XOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n390) );
  NAND2_X1 U482 ( .A1(n464), .A2(G210), .ZN(n389) );
  XNOR2_X1 U483 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U484 ( .A(n391), .B(KEYINPUT92), .Z(n396) );
  XNOR2_X1 U485 ( .A(n393), .B(n392), .ZN(n448) );
  XNOR2_X1 U486 ( .A(G113), .B(G137), .ZN(n394) );
  XNOR2_X1 U487 ( .A(n448), .B(n394), .ZN(n395) );
  XNOR2_X1 U488 ( .A(n396), .B(n395), .ZN(n397) );
  INV_X1 U489 ( .A(G902), .ZN(n454) );
  NAND2_X1 U490 ( .A1(n673), .A2(n454), .ZN(n399) );
  INV_X1 U491 ( .A(G472), .ZN(n398) );
  XNOR2_X2 U492 ( .A(n399), .B(n398), .ZN(n577) );
  XNOR2_X1 U493 ( .A(KEYINPUT15), .B(G902), .ZN(n639) );
  NAND2_X1 U494 ( .A1(G234), .A2(n639), .ZN(n400) );
  XNOR2_X1 U495 ( .A(KEYINPUT20), .B(n400), .ZN(n420) );
  AND2_X1 U496 ( .A1(n420), .A2(G221), .ZN(n401) );
  XNOR2_X1 U497 ( .A(n401), .B(KEYINPUT21), .ZN(n602) );
  INV_X1 U498 ( .A(n602), .ZN(n561) );
  XNOR2_X1 U499 ( .A(n402), .B(KEYINPUT14), .ZN(n403) );
  NAND2_X1 U500 ( .A1(G952), .A2(n403), .ZN(n627) );
  NOR2_X1 U501 ( .A1(n627), .A2(G953), .ZN(n543) );
  NAND2_X1 U502 ( .A1(n403), .A2(G902), .ZN(n405) );
  OR2_X1 U503 ( .A1(n735), .A2(n542), .ZN(n406) );
  XNOR2_X1 U504 ( .A(KEYINPUT98), .B(n406), .ZN(n407) );
  NOR2_X1 U505 ( .A1(G900), .A2(n407), .ZN(n408) );
  NOR2_X1 U506 ( .A1(n543), .A2(n408), .ZN(n493) );
  NOR2_X1 U507 ( .A1(n561), .A2(n493), .ZN(n410) );
  NAND2_X1 U508 ( .A1(G234), .A2(n735), .ZN(n411) );
  XOR2_X1 U509 ( .A(KEYINPUT8), .B(n411), .Z(n478) );
  NAND2_X1 U510 ( .A1(G221), .A2(n478), .ZN(n413) );
  XOR2_X1 U511 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n412) );
  XNOR2_X1 U512 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U513 ( .A(KEYINPUT88), .B(G110), .Z(n415) );
  XOR2_X1 U514 ( .A(n415), .B(n414), .Z(n416) );
  XNOR2_X1 U515 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U516 ( .A(G137), .B(G140), .Z(n429) );
  NAND2_X1 U517 ( .A1(n663), .A2(n454), .ZN(n425) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(KEYINPUT89), .Z(n422) );
  NAND2_X1 U519 ( .A1(n420), .A2(G217), .ZN(n421) );
  XNOR2_X1 U520 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U521 ( .A(n423), .B(KEYINPUT70), .ZN(n424) );
  XNOR2_X2 U522 ( .A(n425), .B(n424), .ZN(n576) );
  NAND2_X1 U523 ( .A1(n514), .A2(n576), .ZN(n426) );
  NOR2_X1 U524 ( .A1(n577), .A2(n426), .ZN(n428) );
  XNOR2_X1 U525 ( .A(KEYINPUT102), .B(KEYINPUT28), .ZN(n427) );
  XNOR2_X1 U526 ( .A(n428), .B(n427), .ZN(n440) );
  XOR2_X1 U527 ( .A(n429), .B(G110), .Z(n430) );
  NAND2_X1 U528 ( .A1(G227), .A2(n735), .ZN(n434) );
  XOR2_X1 U529 ( .A(G101), .B(G107), .Z(n435) );
  NOR2_X1 U530 ( .A1(G902), .A2(n655), .ZN(n439) );
  INV_X1 U531 ( .A(G469), .ZN(n438) );
  XNOR2_X1 U532 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n443) );
  XNOR2_X1 U533 ( .A(n445), .B(n446), .ZN(n452) );
  INV_X1 U534 ( .A(G113), .ZN(n447) );
  XNOR2_X1 U535 ( .A(n447), .B(G104), .ZN(n469) );
  XNOR2_X1 U536 ( .A(n448), .B(n469), .ZN(n451) );
  XNOR2_X1 U537 ( .A(G122), .B(G107), .ZN(n479) );
  XNOR2_X1 U538 ( .A(KEYINPUT16), .B(G110), .ZN(n449) );
  XNOR2_X1 U539 ( .A(n479), .B(n449), .ZN(n450) );
  XNOR2_X1 U540 ( .A(n451), .B(n450), .ZN(n725) );
  XNOR2_X1 U541 ( .A(n452), .B(n725), .ZN(n649) );
  NAND2_X1 U542 ( .A1(n454), .A2(n453), .ZN(n458) );
  NAND2_X1 U543 ( .A1(n458), .A2(G210), .ZN(n456) );
  INV_X1 U544 ( .A(KEYINPUT85), .ZN(n455) );
  XNOR2_X1 U545 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U546 ( .A1(n458), .A2(G214), .ZN(n614) );
  INV_X1 U547 ( .A(n614), .ZN(n459) );
  XNOR2_X2 U548 ( .A(n460), .B(KEYINPUT19), .ZN(n690) );
  XNOR2_X1 U549 ( .A(G143), .B(n461), .ZN(n473) );
  XOR2_X1 U550 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n463) );
  XNOR2_X1 U551 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n462) );
  XNOR2_X1 U552 ( .A(n463), .B(n462), .ZN(n468) );
  NAND2_X1 U553 ( .A1(G214), .A2(n464), .ZN(n465) );
  XNOR2_X1 U554 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U555 ( .A(n468), .B(n467), .ZN(n471) );
  XOR2_X1 U556 ( .A(G122), .B(n469), .Z(n470) );
  XOR2_X1 U557 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n475) );
  XNOR2_X1 U558 ( .A(G116), .B(KEYINPUT95), .ZN(n474) );
  XNOR2_X1 U559 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U560 ( .A(n477), .B(n476), .ZN(n483) );
  NAND2_X1 U561 ( .A1(G217), .A2(n478), .ZN(n481) );
  XNOR2_X1 U562 ( .A(n479), .B(G134), .ZN(n480) );
  XNOR2_X1 U563 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U564 ( .A(n483), .B(n482), .ZN(n715) );
  NOR2_X1 U565 ( .A1(G902), .A2(n715), .ZN(n484) );
  XNOR2_X1 U566 ( .A(G478), .B(n484), .ZN(n490) );
  NOR2_X1 U567 ( .A1(n501), .A2(n490), .ZN(n697) );
  NOR2_X1 U568 ( .A1(n697), .A2(n513), .ZN(n619) );
  INV_X1 U569 ( .A(n619), .ZN(n485) );
  NAND2_X1 U570 ( .A1(n690), .A2(n485), .ZN(n486) );
  NOR2_X1 U571 ( .A1(n692), .A2(n486), .ZN(n487) );
  NOR2_X1 U572 ( .A1(n488), .A2(n487), .ZN(n489) );
  NOR2_X1 U573 ( .A1(KEYINPUT47), .A2(n489), .ZN(n499) );
  INV_X1 U574 ( .A(n490), .ZN(n500) );
  NAND2_X1 U575 ( .A1(n501), .A2(n500), .ZN(n549) );
  NAND2_X1 U576 ( .A1(n606), .A2(n614), .ZN(n491) );
  XNOR2_X1 U577 ( .A(KEYINPUT30), .B(n491), .ZN(n492) );
  NOR2_X1 U578 ( .A1(n493), .A2(n492), .ZN(n496) );
  XNOR2_X1 U579 ( .A(n495), .B(KEYINPUT90), .ZN(n556) );
  NAND2_X1 U580 ( .A1(n496), .A2(n556), .ZN(n508) );
  NOR2_X1 U581 ( .A1(n508), .A2(n534), .ZN(n497) );
  XNOR2_X1 U582 ( .A(n497), .B(KEYINPUT101), .ZN(n498) );
  NOR2_X1 U583 ( .A1(n549), .A2(n498), .ZN(n689) );
  NOR2_X1 U584 ( .A1(n499), .A2(n385), .ZN(n512) );
  NOR2_X1 U585 ( .A1(n501), .A2(n500), .ZN(n503) );
  INV_X1 U586 ( .A(KEYINPUT96), .ZN(n502) );
  XNOR2_X1 U587 ( .A(n503), .B(n502), .ZN(n617) );
  XOR2_X1 U588 ( .A(KEYINPUT38), .B(n534), .Z(n507) );
  INV_X1 U589 ( .A(n507), .ZN(n615) );
  NAND2_X1 U590 ( .A1(n615), .A2(n614), .ZN(n618) );
  NOR2_X1 U591 ( .A1(n617), .A2(n618), .ZN(n504) );
  XNOR2_X1 U592 ( .A(KEYINPUT41), .B(n504), .ZN(n628) );
  OR2_X1 U593 ( .A1(n628), .A2(n692), .ZN(n506) );
  XOR2_X1 U594 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n505) );
  NOR2_X2 U595 ( .A1(n508), .A2(n507), .ZN(n510) );
  XOR2_X1 U596 ( .A(KEYINPUT68), .B(KEYINPUT39), .Z(n509) );
  XNOR2_X1 U597 ( .A(n510), .B(n509), .ZN(n530) );
  AND2_X1 U598 ( .A1(n530), .A2(n513), .ZN(n511) );
  XNOR2_X1 U599 ( .A(n511), .B(KEYINPUT40), .ZN(n744) );
  INV_X1 U600 ( .A(n570), .ZN(n515) );
  XOR2_X1 U601 ( .A(KEYINPUT97), .B(n513), .Z(n695) );
  INV_X1 U602 ( .A(n534), .ZN(n516) );
  NAND2_X1 U603 ( .A1(n352), .A2(n516), .ZN(n518) );
  XNOR2_X1 U604 ( .A(KEYINPUT105), .B(KEYINPUT36), .ZN(n517) );
  XNOR2_X1 U605 ( .A(n518), .B(n517), .ZN(n522) );
  INV_X1 U606 ( .A(KEYINPUT1), .ZN(n519) );
  INV_X1 U607 ( .A(n553), .ZN(n539) );
  NAND2_X1 U608 ( .A1(n522), .A2(n572), .ZN(n703) );
  NAND2_X1 U609 ( .A1(KEYINPUT74), .A2(n619), .ZN(n523) );
  NAND2_X1 U610 ( .A1(n690), .A2(n523), .ZN(n524) );
  OR2_X1 U611 ( .A1(n692), .A2(n524), .ZN(n525) );
  NAND2_X1 U612 ( .A1(n525), .A2(KEYINPUT47), .ZN(n526) );
  INV_X1 U613 ( .A(KEYINPUT48), .ZN(n527) );
  NAND2_X1 U614 ( .A1(n697), .A2(n530), .ZN(n704) );
  XOR2_X1 U615 ( .A(KEYINPUT43), .B(KEYINPUT100), .Z(n533) );
  XNOR2_X1 U616 ( .A(KEYINPUT99), .B(n352), .ZN(n531) );
  NOR2_X1 U617 ( .A1(n539), .A2(n531), .ZN(n532) );
  XNOR2_X1 U618 ( .A(n533), .B(n532), .ZN(n535) );
  NAND2_X1 U619 ( .A1(n535), .A2(n534), .ZN(n671) );
  AND2_X1 U620 ( .A1(n704), .A2(n671), .ZN(n593) );
  AND2_X1 U621 ( .A1(n593), .A2(KEYINPUT2), .ZN(n536) );
  NAND2_X1 U622 ( .A1(n594), .A2(n536), .ZN(n538) );
  INV_X1 U623 ( .A(KEYINPUT76), .ZN(n537) );
  XNOR2_X1 U624 ( .A(n538), .B(n537), .ZN(n592) );
  AND2_X1 U625 ( .A1(n570), .A2(n494), .ZN(n540) );
  NAND2_X1 U626 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U627 ( .A(G898), .B(KEYINPUT86), .Z(n722) );
  NAND2_X1 U628 ( .A1(G953), .A2(n722), .ZN(n726) );
  OR2_X1 U629 ( .A1(n542), .A2(n726), .ZN(n545) );
  INV_X1 U630 ( .A(n543), .ZN(n544) );
  NAND2_X1 U631 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U632 ( .A1(n690), .A2(n546), .ZN(n547) );
  XNOR2_X1 U633 ( .A(n548), .B(KEYINPUT34), .ZN(n551) );
  INV_X1 U634 ( .A(n549), .ZN(n550) );
  NAND2_X1 U635 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X2 U636 ( .A(n552), .B(KEYINPUT35), .ZN(n742) );
  NAND2_X1 U637 ( .A1(n742), .A2(KEYINPUT44), .ZN(n568) );
  NOR2_X1 U638 ( .A1(n598), .A2(n599), .ZN(n554) );
  NAND2_X1 U639 ( .A1(n554), .A2(n606), .ZN(n609) );
  OR2_X1 U640 ( .A1(n609), .A2(n563), .ZN(n555) );
  XNOR2_X1 U641 ( .A(n555), .B(KEYINPUT31), .ZN(n698) );
  AND2_X1 U642 ( .A1(n556), .A2(n577), .ZN(n558) );
  INV_X1 U643 ( .A(n563), .ZN(n557) );
  NOR2_X1 U644 ( .A1(n698), .A2(n386), .ZN(n559) );
  OR2_X1 U645 ( .A1(n559), .A2(n619), .ZN(n566) );
  NOR2_X1 U646 ( .A1(n570), .A2(n576), .ZN(n560) );
  NAND2_X1 U647 ( .A1(n598), .A2(n560), .ZN(n565) );
  OR2_X1 U648 ( .A1(n617), .A2(n561), .ZN(n562) );
  XNOR2_X1 U649 ( .A(KEYINPUT69), .B(KEYINPUT22), .ZN(n564) );
  OR2_X1 U650 ( .A1(n565), .A2(n579), .ZN(n669) );
  AND2_X1 U651 ( .A1(n566), .A2(n669), .ZN(n567) );
  NAND2_X1 U652 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U653 ( .A(n569), .B(KEYINPUT79), .ZN(n590) );
  NOR2_X1 U654 ( .A1(n570), .A2(n603), .ZN(n571) );
  XNOR2_X1 U655 ( .A(n573), .B(KEYINPUT72), .ZN(n574) );
  XNOR2_X1 U656 ( .A(n575), .B(KEYINPUT32), .ZN(n672) );
  AND2_X1 U657 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n598), .A2(n578), .ZN(n580) );
  OR2_X1 U659 ( .A1(n580), .A2(n579), .ZN(n670) );
  NAND2_X1 U660 ( .A1(n672), .A2(n670), .ZN(n582) );
  INV_X1 U661 ( .A(KEYINPUT80), .ZN(n581) );
  INV_X1 U662 ( .A(n585), .ZN(n584) );
  INV_X1 U663 ( .A(KEYINPUT44), .ZN(n583) );
  NAND2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X2 U668 ( .A(n591), .B(KEYINPUT45), .ZN(n641) );
  NAND2_X1 U669 ( .A1(n592), .A2(n641), .ZN(n645) );
  NAND2_X1 U670 ( .A1(n641), .A2(n733), .ZN(n596) );
  XNOR2_X1 U671 ( .A(KEYINPUT73), .B(KEYINPUT2), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n645), .A2(n597), .ZN(n633) );
  XNOR2_X1 U674 ( .A(KEYINPUT114), .B(KEYINPUT51), .ZN(n612) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U676 ( .A(KEYINPUT113), .B(n600), .Z(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT50), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U679 ( .A(KEYINPUT49), .B(n604), .Z(n605) );
  NOR2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n628), .A2(n613), .ZN(n624) );
  NOR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n622) );
  NOR2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U688 ( .A(KEYINPUT115), .B(n620), .Z(n621) );
  NOR2_X1 U689 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U690 ( .A1(n624), .A2(n356), .ZN(n625) );
  XNOR2_X1 U691 ( .A(n625), .B(KEYINPUT52), .ZN(n626) );
  NOR2_X1 U692 ( .A1(n627), .A2(n626), .ZN(n630) );
  NOR2_X1 U693 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U694 ( .A(n631), .B(KEYINPUT116), .ZN(n632) );
  NAND2_X1 U695 ( .A1(n633), .A2(n632), .ZN(n635) );
  NOR2_X1 U696 ( .A1(G953), .A2(n636), .ZN(n638) );
  XNOR2_X1 U697 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n637) );
  NAND2_X1 U698 ( .A1(n640), .A2(n381), .ZN(n642) );
  INV_X1 U699 ( .A(n641), .ZN(n719) );
  NOR2_X1 U700 ( .A1(n642), .A2(n719), .ZN(n644) );
  AND2_X1 U701 ( .A1(n381), .A2(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U702 ( .A1(n713), .A2(G210), .ZN(n651) );
  XOR2_X1 U703 ( .A(KEYINPUT82), .B(KEYINPUT55), .Z(n647) );
  XNOR2_X1 U704 ( .A(n647), .B(KEYINPUT54), .ZN(n648) );
  XNOR2_X1 U705 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U706 ( .A(n651), .B(n650), .ZN(n653) );
  INV_X1 U707 ( .A(G952), .ZN(n652) );
  AND2_X1 U708 ( .A1(n652), .A2(G953), .ZN(n718) );
  NOR2_X2 U709 ( .A1(n653), .A2(n718), .ZN(n654) );
  XNOR2_X1 U710 ( .A(n654), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U711 ( .A1(n713), .A2(G469), .ZN(n659) );
  XNOR2_X1 U712 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n657) );
  XNOR2_X1 U713 ( .A(n655), .B(KEYINPUT57), .ZN(n656) );
  XNOR2_X1 U714 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U715 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X2 U716 ( .A1(n660), .A2(n718), .ZN(n661) );
  XNOR2_X1 U717 ( .A(n661), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U718 ( .A1(n713), .A2(G217), .ZN(n665) );
  XNOR2_X1 U719 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n662) );
  XNOR2_X1 U720 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U721 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X2 U722 ( .A1(n666), .A2(n718), .ZN(n668) );
  XNOR2_X1 U723 ( .A(n668), .B(n667), .ZN(G66) );
  XNOR2_X1 U724 ( .A(n669), .B(G101), .ZN(G3) );
  XNOR2_X1 U725 ( .A(n670), .B(G110), .ZN(G12) );
  XNOR2_X1 U726 ( .A(n671), .B(G140), .ZN(G42) );
  XNOR2_X1 U727 ( .A(n672), .B(G119), .ZN(G21) );
  NAND2_X1 U728 ( .A1(n713), .A2(G472), .ZN(n675) );
  XOR2_X1 U729 ( .A(KEYINPUT62), .B(n673), .Z(n674) );
  XNOR2_X1 U730 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X2 U731 ( .A1(n676), .A2(n718), .ZN(n678) );
  XNOR2_X1 U732 ( .A(KEYINPUT81), .B(KEYINPUT63), .ZN(n677) );
  XNOR2_X1 U733 ( .A(n678), .B(n677), .ZN(G57) );
  NAND2_X1 U734 ( .A1(n386), .A2(n695), .ZN(n679) );
  XNOR2_X1 U735 ( .A(n679), .B(G104), .ZN(G6) );
  NAND2_X1 U736 ( .A1(n386), .A2(n697), .ZN(n685) );
  XOR2_X1 U737 ( .A(KEYINPUT108), .B(KEYINPUT27), .Z(n681) );
  XNOR2_X1 U738 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n681), .B(n680), .ZN(n683) );
  XOR2_X1 U740 ( .A(G107), .B(KEYINPUT26), .Z(n682) );
  XNOR2_X1 U741 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U742 ( .A(n685), .B(n684), .ZN(G9) );
  XOR2_X1 U743 ( .A(G128), .B(KEYINPUT29), .Z(n688) );
  NAND2_X1 U744 ( .A1(n690), .A2(n697), .ZN(n686) );
  OR2_X1 U745 ( .A1(n692), .A2(n686), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n688), .B(n687), .ZN(G30) );
  XOR2_X1 U747 ( .A(G143), .B(n689), .Z(G45) );
  NAND2_X1 U748 ( .A1(n690), .A2(n695), .ZN(n691) );
  NOR2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U750 ( .A(G146), .B(KEYINPUT109), .ZN(n693) );
  XNOR2_X1 U751 ( .A(n694), .B(n693), .ZN(G48) );
  NAND2_X1 U752 ( .A1(n695), .A2(n698), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n696), .B(G113), .ZN(G15) );
  XOR2_X1 U754 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n700) );
  NAND2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U756 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U757 ( .A(G116), .B(n701), .ZN(G18) );
  XOR2_X1 U758 ( .A(G125), .B(KEYINPUT37), .Z(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(n702), .ZN(G27) );
  XNOR2_X1 U760 ( .A(G134), .B(KEYINPUT112), .ZN(n705) );
  XNOR2_X1 U761 ( .A(n705), .B(n704), .ZN(G36) );
  NAND2_X1 U762 ( .A1(n713), .A2(G475), .ZN(n708) );
  XOR2_X1 U763 ( .A(n706), .B(KEYINPUT59), .Z(n707) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X2 U765 ( .A1(n709), .A2(n718), .ZN(n712) );
  XNOR2_X1 U766 ( .A(KEYINPUT65), .B(KEYINPUT121), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n710), .B(KEYINPUT60), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n712), .B(n711), .ZN(G60) );
  NAND2_X1 U769 ( .A1(n713), .A2(G478), .ZN(n714) );
  XNOR2_X1 U770 ( .A(n714), .B(KEYINPUT122), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n718), .A2(n717), .ZN(G63) );
  NOR2_X1 U773 ( .A1(n719), .A2(G953), .ZN(n724) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n720) );
  XOR2_X1 U775 ( .A(KEYINPUT61), .B(n720), .Z(n721) );
  NOR2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n730) );
  XOR2_X1 U778 ( .A(KEYINPUT127), .B(n725), .Z(n727) );
  NAND2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(KEYINPUT126), .ZN(n729) );
  XNOR2_X1 U781 ( .A(n730), .B(n729), .ZN(G69) );
  XNOR2_X1 U782 ( .A(n732), .B(n731), .ZN(n737) );
  INV_X1 U783 ( .A(n737), .ZN(n734) );
  XOR2_X1 U784 ( .A(n734), .B(n733), .Z(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(n735), .ZN(n741) );
  XOR2_X1 U786 ( .A(G227), .B(n737), .Z(n738) );
  NAND2_X1 U787 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U789 ( .A1(n741), .A2(n740), .ZN(G72) );
  XOR2_X1 U790 ( .A(n742), .B(G122), .Z(G24) );
  XOR2_X1 U791 ( .A(G137), .B(n743), .Z(G39) );
  XOR2_X1 U792 ( .A(n744), .B(G131), .Z(G33) );
endmodule

