

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734;

  INV_X1 U369 ( .A(G146), .ZN(n389) );
  NOR2_X1 U370 ( .A1(n576), .A2(n547), .ZN(n562) );
  XNOR2_X1 U371 ( .A(n470), .B(n660), .ZN(n528) );
  INV_X1 U372 ( .A(n437), .ZN(n725) );
  NOR2_X1 U373 ( .A1(n528), .A2(n484), .ZN(n347) );
  NOR2_X2 U374 ( .A1(n595), .A2(n594), .ZN(n616) );
  AND2_X2 U375 ( .A1(n484), .A2(n528), .ZN(n588) );
  OR2_X1 U376 ( .A1(n543), .A2(n548), .ZN(n544) );
  XNOR2_X1 U377 ( .A(n450), .B(n449), .ZN(n596) );
  AND2_X1 U378 ( .A1(n364), .A2(n382), .ZN(n366) );
  NOR2_X1 U379 ( .A1(n617), .A2(n598), .ZN(n691) );
  AND2_X1 U380 ( .A1(n381), .A2(n580), .ZN(n675) );
  NOR2_X1 U381 ( .A1(n596), .A2(n512), .ZN(n379) );
  XNOR2_X1 U382 ( .A(G113), .B(G131), .ZN(n454) );
  XOR2_X1 U383 ( .A(KEYINPUT4), .B(KEYINPUT68), .Z(n433) );
  OR2_X1 U384 ( .A1(n697), .A2(G902), .ZN(n376) );
  NAND2_X1 U385 ( .A1(n429), .A2(n531), .ZN(n430) );
  XNOR2_X1 U386 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n586) );
  NOR2_X1 U387 ( .A1(n607), .A2(KEYINPUT47), .ZN(n604) );
  INV_X1 U388 ( .A(G104), .ZN(n453) );
  NAND2_X1 U389 ( .A1(n373), .A2(n348), .ZN(n372) );
  XNOR2_X1 U390 ( .A(n389), .B(G125), .ZN(n432) );
  NOR2_X1 U391 ( .A1(n640), .A2(KEYINPUT81), .ZN(n384) );
  XNOR2_X1 U392 ( .A(n378), .B(n481), .ZN(n721) );
  XNOR2_X1 U393 ( .A(n387), .B(n388), .ZN(n378) );
  XNOR2_X1 U394 ( .A(G137), .B(G131), .ZN(n388) );
  INV_X1 U395 ( .A(n433), .ZN(n387) );
  XNOR2_X1 U396 ( .A(n376), .B(n352), .ZN(n531) );
  INV_X1 U397 ( .A(n376), .ZN(n546) );
  NOR2_X1 U398 ( .A1(n654), .A2(G902), .ZN(n399) );
  XNOR2_X1 U399 ( .A(n360), .B(n359), .ZN(n443) );
  XNOR2_X1 U400 ( .A(n393), .B(n395), .ZN(n359) );
  XNOR2_X1 U401 ( .A(n394), .B(n396), .ZN(n360) );
  XOR2_X1 U402 ( .A(G110), .B(G128), .Z(n408) );
  XNOR2_X1 U403 ( .A(n432), .B(n371), .ZN(n722) );
  XNOR2_X1 U404 ( .A(KEYINPUT10), .B(G140), .ZN(n371) );
  XNOR2_X1 U405 ( .A(n406), .B(n405), .ZN(n477) );
  NAND2_X1 U406 ( .A1(n725), .A2(G234), .ZN(n406) );
  XNOR2_X1 U407 ( .A(n721), .B(n389), .ZN(n421) );
  XOR2_X1 U408 ( .A(G140), .B(G101), .Z(n423) );
  INV_X1 U409 ( .A(G110), .ZN(n424) );
  XNOR2_X1 U410 ( .A(n716), .B(n356), .ZN(n647) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n436), .B(n435), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n440), .B(n439), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n367), .B(n574), .ZN(n614) );
  XNOR2_X1 U415 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n574) );
  NOR2_X1 U416 ( .A1(n524), .A2(n548), .ZN(n526) );
  OR2_X1 U417 ( .A1(n705), .A2(G902), .ZN(n370) );
  NOR2_X1 U418 ( .A1(n627), .A2(n375), .ZN(n374) );
  NAND2_X1 U419 ( .A1(n631), .A2(n351), .ZN(n375) );
  INV_X1 U420 ( .A(G902), .ZN(n446) );
  XNOR2_X1 U421 ( .A(n380), .B(KEYINPUT94), .ZN(n551) );
  NOR2_X1 U422 ( .A1(n688), .A2(n675), .ZN(n380) );
  AND2_X1 U423 ( .A1(n578), .A2(n577), .ZN(n590) );
  XNOR2_X1 U424 ( .A(G902), .B(KEYINPUT15), .ZN(n640) );
  XNOR2_X1 U425 ( .A(n613), .B(KEYINPUT48), .ZN(n629) );
  XOR2_X1 U426 ( .A(KEYINPUT96), .B(G122), .Z(n455) );
  XNOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n434) );
  XOR2_X1 U428 ( .A(G143), .B(G128), .Z(n435) );
  XNOR2_X1 U429 ( .A(G116), .B(G122), .ZN(n471) );
  XOR2_X1 U430 ( .A(KEYINPUT7), .B(G107), .Z(n472) );
  XNOR2_X1 U431 ( .A(KEYINPUT9), .B(KEYINPUT101), .ZN(n473) );
  XOR2_X1 U432 ( .A(KEYINPUT100), .B(KEYINPUT102), .Z(n474) );
  XNOR2_X1 U433 ( .A(n377), .B(G134), .ZN(n481) );
  XNOR2_X1 U434 ( .A(G143), .B(G128), .ZN(n377) );
  NAND2_X1 U435 ( .A1(n366), .A2(n365), .ZN(n645) );
  AND2_X1 U436 ( .A1(n572), .A2(n571), .ZN(n610) );
  NOR2_X1 U437 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U438 ( .A(n592), .ZN(n569) );
  XNOR2_X1 U439 ( .A(n444), .B(n443), .ZN(n716) );
  XNOR2_X1 U440 ( .A(KEYINPUT16), .B(G122), .ZN(n441) );
  XNOR2_X1 U441 ( .A(n409), .B(n385), .ZN(n414) );
  XNOR2_X1 U442 ( .A(n421), .B(n353), .ZN(n697) );
  AND2_X1 U443 ( .A1(n437), .A2(n650), .ZN(n709) );
  XNOR2_X1 U444 ( .A(n597), .B(KEYINPUT36), .ZN(n598) );
  XNOR2_X1 U445 ( .A(n530), .B(KEYINPUT35), .ZN(n732) );
  XNOR2_X1 U446 ( .A(n362), .B(n541), .ZN(n637) );
  NOR2_X1 U447 ( .A1(n601), .A2(n600), .ZN(n683) );
  OR2_X1 U448 ( .A1(n555), .A2(n542), .ZN(n361) );
  XNOR2_X1 U449 ( .A(n374), .B(KEYINPUT122), .ZN(n633) );
  AND2_X1 U450 ( .A1(n637), .A2(n361), .ZN(n348) );
  XOR2_X1 U451 ( .A(n399), .B(G472), .Z(n563) );
  AND2_X1 U452 ( .A1(n724), .A2(n384), .ZN(n349) );
  OR2_X1 U453 ( .A1(n372), .A2(KEYINPUT44), .ZN(n350) );
  NOR2_X1 U454 ( .A1(n632), .A2(n626), .ZN(n351) );
  XOR2_X1 U455 ( .A(n428), .B(KEYINPUT1), .Z(n352) );
  XOR2_X1 U456 ( .A(n427), .B(n426), .Z(n353) );
  XOR2_X1 U457 ( .A(n612), .B(KEYINPUT80), .Z(n354) );
  OR2_X2 U458 ( .A1(n577), .A2(n420), .ZN(n547) );
  XOR2_X1 U459 ( .A(n513), .B(KEYINPUT19), .Z(n355) );
  XOR2_X2 U460 ( .A(n588), .B(KEYINPUT105), .Z(n686) );
  INV_X1 U461 ( .A(n361), .ZN(n678) );
  NAND2_X1 U462 ( .A1(n363), .A2(n617), .ZN(n555) );
  NAND2_X1 U463 ( .A1(n363), .A2(n539), .ZN(n362) );
  XNOR2_X1 U464 ( .A(n538), .B(KEYINPUT22), .ZN(n363) );
  NAND2_X1 U465 ( .A1(n349), .A2(n711), .ZN(n364) );
  NAND2_X1 U466 ( .A1(n711), .A2(n724), .ZN(n639) );
  NAND2_X1 U467 ( .A1(n639), .A2(KEYINPUT81), .ZN(n365) );
  NAND2_X1 U468 ( .A1(n614), .A2(n588), .ZN(n575) );
  NAND2_X1 U469 ( .A1(n610), .A2(n573), .ZN(n367) );
  NAND2_X1 U470 ( .A1(n369), .A2(n368), .ZN(n613) );
  XNOR2_X1 U471 ( .A(n587), .B(n586), .ZN(n368) );
  AND2_X1 U472 ( .A1(n606), .A2(n354), .ZN(n369) );
  XNOR2_X2 U473 ( .A(n370), .B(n415), .ZN(n577) );
  NAND2_X1 U474 ( .A1(n372), .A2(KEYINPUT44), .ZN(n558) );
  INV_X1 U475 ( .A(n732), .ZN(n373) );
  INV_X1 U476 ( .A(n644), .ZN(n624) );
  NAND2_X1 U477 ( .A1(n630), .A2(n711), .ZN(n644) );
  XNOR2_X2 U478 ( .A(n561), .B(KEYINPUT45), .ZN(n711) );
  NAND2_X1 U479 ( .A1(n599), .A2(n522), .ZN(n523) );
  XNOR2_X1 U480 ( .A(n379), .B(n355), .ZN(n599) );
  XNOR2_X1 U481 ( .A(n550), .B(KEYINPUT92), .ZN(n381) );
  AND2_X1 U482 ( .A1(n643), .A2(n383), .ZN(n382) );
  NAND2_X1 U483 ( .A1(n640), .A2(KEYINPUT81), .ZN(n383) );
  INV_X2 U484 ( .A(n661), .ZN(n704) );
  NAND2_X1 U485 ( .A1(n645), .A2(n644), .ZN(n661) );
  XOR2_X1 U486 ( .A(n408), .B(n407), .Z(n385) );
  XNOR2_X1 U487 ( .A(n454), .B(n453), .ZN(n456) );
  XNOR2_X1 U488 ( .A(n456), .B(n455), .ZN(n458) );
  INV_X1 U489 ( .A(KEYINPUT8), .ZN(n405) );
  AND2_X1 U490 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U491 ( .A(G469), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n705), .B(KEYINPUT124), .ZN(n706) );
  XNOR2_X1 U493 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U494 ( .A(n635), .B(n634), .ZN(G75) );
  NAND2_X1 U495 ( .A1(G234), .A2(G237), .ZN(n386) );
  XNOR2_X1 U496 ( .A(n386), .B(KEYINPUT14), .ZN(n518) );
  NAND2_X1 U497 ( .A1(G952), .A2(n518), .ZN(n514) );
  XOR2_X1 U498 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n510) );
  XOR2_X1 U499 ( .A(KEYINPUT5), .B(KEYINPUT74), .Z(n391) );
  NOR2_X1 U500 ( .A1(G953), .A2(G237), .ZN(n461) );
  NAND2_X1 U501 ( .A1(n461), .A2(G210), .ZN(n390) );
  XNOR2_X1 U502 ( .A(n391), .B(n390), .ZN(n397) );
  INV_X1 U503 ( .A(G113), .ZN(n392) );
  XNOR2_X1 U504 ( .A(n392), .B(G101), .ZN(n394) );
  XNOR2_X1 U505 ( .A(G119), .B(G116), .ZN(n393) );
  XNOR2_X1 U506 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n396) );
  XNOR2_X1 U507 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n395) );
  XOR2_X1 U508 ( .A(n397), .B(n443), .Z(n398) );
  XNOR2_X1 U509 ( .A(n421), .B(n398), .ZN(n654) );
  XNOR2_X1 U510 ( .A(KEYINPUT6), .B(KEYINPUT104), .ZN(n400) );
  XNOR2_X1 U511 ( .A(n563), .B(n400), .ZN(n553) );
  INV_X1 U512 ( .A(n553), .ZN(n593) );
  XOR2_X1 U513 ( .A(KEYINPUT75), .B(KEYINPUT90), .Z(n403) );
  NAND2_X1 U514 ( .A1(n640), .A2(G234), .ZN(n401) );
  XNOR2_X1 U515 ( .A(n401), .B(KEYINPUT20), .ZN(n416) );
  NAND2_X1 U516 ( .A1(n416), .A2(G217), .ZN(n402) );
  XNOR2_X1 U517 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U518 ( .A(KEYINPUT25), .B(n404), .ZN(n415) );
  XNOR2_X2 U519 ( .A(KEYINPUT64), .B(G953), .ZN(n437) );
  NAND2_X1 U520 ( .A1(G221), .A2(n477), .ZN(n409) );
  XNOR2_X1 U521 ( .A(G119), .B(G137), .ZN(n407) );
  XOR2_X1 U522 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n411) );
  XNOR2_X1 U523 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n410) );
  XNOR2_X1 U524 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U525 ( .A(n722), .B(n412), .Z(n413) );
  XNOR2_X1 U526 ( .A(n414), .B(n413), .ZN(n705) );
  NAND2_X1 U527 ( .A1(n416), .A2(G221), .ZN(n418) );
  INV_X1 U528 ( .A(KEYINPUT21), .ZN(n417) );
  XNOR2_X1 U529 ( .A(n418), .B(n417), .ZN(n578) );
  INV_X1 U530 ( .A(KEYINPUT91), .ZN(n419) );
  XNOR2_X1 U531 ( .A(n578), .B(n419), .ZN(n535) );
  INV_X1 U532 ( .A(n535), .ZN(n420) );
  INV_X1 U533 ( .A(n547), .ZN(n429) );
  NAND2_X1 U534 ( .A1(G227), .A2(n725), .ZN(n422) );
  XNOR2_X1 U535 ( .A(n423), .B(n422), .ZN(n427) );
  XNOR2_X1 U536 ( .A(G104), .B(G107), .ZN(n425) );
  XNOR2_X1 U537 ( .A(n425), .B(n424), .ZN(n442) );
  INV_X1 U538 ( .A(n442), .ZN(n426) );
  INV_X1 U539 ( .A(n531), .ZN(n617) );
  NOR2_X1 U540 ( .A1(n553), .A2(n430), .ZN(n431) );
  XNOR2_X1 U541 ( .A(n431), .B(KEYINPUT33), .ZN(n524) );
  INV_X1 U542 ( .A(n524), .ZN(n491) );
  XNOR2_X1 U543 ( .A(n433), .B(n432), .ZN(n440) );
  XNOR2_X1 U544 ( .A(n434), .B(KEYINPUT76), .ZN(n436) );
  INV_X1 U545 ( .A(G224), .ZN(n438) );
  OR2_X1 U546 ( .A1(n437), .A2(n438), .ZN(n439) );
  XNOR2_X1 U547 ( .A(n442), .B(n441), .ZN(n444) );
  NAND2_X1 U548 ( .A1(n647), .A2(n640), .ZN(n450) );
  INV_X1 U549 ( .A(G237), .ZN(n445) );
  NAND2_X1 U550 ( .A1(n446), .A2(n445), .ZN(n451) );
  NAND2_X1 U551 ( .A1(n451), .A2(G210), .ZN(n448) );
  INV_X1 U552 ( .A(KEYINPUT85), .ZN(n447) );
  XNOR2_X1 U553 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U554 ( .A(n596), .B(KEYINPUT38), .ZN(n573) );
  NAND2_X1 U555 ( .A1(n451), .A2(G214), .ZN(n589) );
  NOR2_X1 U556 ( .A1(n573), .A2(n589), .ZN(n452) );
  XNOR2_X1 U557 ( .A(KEYINPUT119), .B(n452), .ZN(n483) );
  XNOR2_X1 U558 ( .A(KEYINPUT98), .B(KEYINPUT95), .ZN(n457) );
  XNOR2_X1 U559 ( .A(n458), .B(n457), .ZN(n460) );
  INV_X1 U560 ( .A(n722), .ZN(n459) );
  XNOR2_X1 U561 ( .A(n460), .B(n459), .ZN(n467) );
  XNOR2_X1 U562 ( .A(G143), .B(KEYINPUT12), .ZN(n463) );
  NAND2_X1 U563 ( .A1(G214), .A2(n461), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n463), .B(n462), .ZN(n465) );
  XOR2_X1 U565 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n464) );
  XNOR2_X1 U566 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n467), .B(n466), .ZN(n662) );
  NOR2_X1 U568 ( .A1(G902), .A2(n662), .ZN(n469) );
  XNOR2_X1 U569 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n468) );
  XNOR2_X1 U570 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U571 ( .A(G475), .ZN(n660) );
  XNOR2_X1 U572 ( .A(n472), .B(n471), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U574 ( .A(n476), .B(n475), .Z(n479) );
  NAND2_X1 U575 ( .A1(G217), .A2(n477), .ZN(n478) );
  XNOR2_X1 U576 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U577 ( .A(n481), .B(n480), .ZN(n701) );
  NOR2_X1 U578 ( .A1(G902), .A2(n701), .ZN(n482) );
  XNOR2_X1 U579 ( .A(G478), .B(n482), .ZN(n484) );
  INV_X1 U580 ( .A(n484), .ZN(n527) );
  OR2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n493) );
  INV_X1 U582 ( .A(n493), .ZN(n536) );
  NAND2_X1 U583 ( .A1(n483), .A2(n536), .ZN(n489) );
  NOR2_X1 U584 ( .A1(n347), .A2(n588), .ZN(n486) );
  INV_X1 U585 ( .A(KEYINPUT103), .ZN(n485) );
  XNOR2_X1 U586 ( .A(n486), .B(n485), .ZN(n602) );
  NAND2_X1 U587 ( .A1(n573), .A2(n589), .ZN(n492) );
  NOR2_X1 U588 ( .A1(n602), .A2(n492), .ZN(n487) );
  XOR2_X1 U589 ( .A(KEYINPUT120), .B(n487), .Z(n488) );
  NAND2_X1 U590 ( .A1(n489), .A2(n488), .ZN(n490) );
  NAND2_X1 U591 ( .A1(n491), .A2(n490), .ZN(n508) );
  NOR2_X1 U592 ( .A1(n493), .A2(n492), .ZN(n495) );
  XNOR2_X1 U593 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n494) );
  XNOR2_X1 U594 ( .A(n495), .B(n494), .ZN(n625) );
  INV_X1 U595 ( .A(n563), .ZN(n580) );
  NOR2_X1 U596 ( .A1(n617), .A2(n580), .ZN(n496) );
  NAND2_X1 U597 ( .A1(n496), .A2(n429), .ZN(n543) );
  INV_X1 U598 ( .A(n577), .ZN(n552) );
  NOR2_X1 U599 ( .A1(n552), .A2(n578), .ZN(n497) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(n497), .Z(n501) );
  NAND2_X1 U601 ( .A1(n547), .A2(n617), .ZN(n498) );
  XNOR2_X1 U602 ( .A(n498), .B(KEYINPUT117), .ZN(n499) );
  XNOR2_X1 U603 ( .A(KEYINPUT50), .B(n499), .ZN(n500) );
  NOR2_X1 U604 ( .A1(n501), .A2(n500), .ZN(n502) );
  NAND2_X1 U605 ( .A1(n502), .A2(n580), .ZN(n503) );
  NAND2_X1 U606 ( .A1(n543), .A2(n503), .ZN(n504) );
  XNOR2_X1 U607 ( .A(KEYINPUT51), .B(n504), .ZN(n505) );
  NOR2_X1 U608 ( .A1(n625), .A2(n505), .ZN(n506) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(n506), .Z(n507) );
  NAND2_X1 U610 ( .A1(n508), .A2(n507), .ZN(n509) );
  XOR2_X1 U611 ( .A(n510), .B(n509), .Z(n511) );
  NOR2_X1 U612 ( .A1(n514), .A2(n511), .ZN(n632) );
  INV_X1 U613 ( .A(n589), .ZN(n512) );
  INV_X1 U614 ( .A(KEYINPUT67), .ZN(n513) );
  NOR2_X1 U615 ( .A1(n514), .A2(G953), .ZN(n516) );
  INV_X1 U616 ( .A(KEYINPUT86), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n516), .B(n515), .ZN(n568) );
  INV_X1 U618 ( .A(G953), .ZN(n710) );
  NOR2_X1 U619 ( .A1(n710), .A2(G898), .ZN(n517) );
  XNOR2_X1 U620 ( .A(n517), .B(KEYINPUT87), .ZN(n717) );
  INV_X1 U621 ( .A(n717), .ZN(n520) );
  NAND2_X1 U622 ( .A1(G902), .A2(n518), .ZN(n565) );
  INV_X1 U623 ( .A(n565), .ZN(n519) );
  NAND2_X1 U624 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U625 ( .A1(n568), .A2(n521), .ZN(n522) );
  XNOR2_X2 U626 ( .A(n523), .B(KEYINPUT0), .ZN(n548) );
  XNOR2_X1 U627 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n525) );
  XNOR2_X1 U628 ( .A(n526), .B(n525), .ZN(n529) );
  AND2_X1 U629 ( .A1(n528), .A2(n527), .ZN(n608) );
  NAND2_X1 U630 ( .A1(n529), .A2(n608), .ZN(n530) );
  AND2_X1 U631 ( .A1(n531), .A2(n577), .ZN(n532) );
  NAND2_X1 U632 ( .A1(n532), .A2(n553), .ZN(n534) );
  INV_X1 U633 ( .A(KEYINPUT78), .ZN(n533) );
  XNOR2_X1 U634 ( .A(n534), .B(n533), .ZN(n539) );
  NAND2_X1 U635 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U636 ( .A1(n548), .A2(n537), .ZN(n538) );
  INV_X1 U637 ( .A(KEYINPUT77), .ZN(n540) );
  XNOR2_X1 U638 ( .A(n540), .B(KEYINPUT32), .ZN(n541) );
  NAND2_X1 U639 ( .A1(n580), .A2(n577), .ZN(n542) );
  XOR2_X1 U640 ( .A(KEYINPUT31), .B(KEYINPUT93), .Z(n545) );
  XNOR2_X1 U641 ( .A(n545), .B(n544), .ZN(n688) );
  XNOR2_X1 U642 ( .A(G469), .B(n546), .ZN(n576) );
  INV_X1 U643 ( .A(n562), .ZN(n549) );
  NOR2_X1 U644 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U645 ( .A1(n551), .A2(n602), .ZN(n556) );
  NAND2_X1 U646 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U647 ( .A1(n555), .A2(n554), .ZN(n669) );
  NOR2_X1 U648 ( .A1(n556), .A2(n669), .ZN(n557) );
  NAND2_X1 U649 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U650 ( .A(n559), .B(KEYINPUT83), .ZN(n560) );
  NAND2_X1 U651 ( .A1(n560), .A2(n350), .ZN(n561) );
  XNOR2_X1 U652 ( .A(n562), .B(KEYINPUT106), .ZN(n572) );
  NAND2_X1 U653 ( .A1(n563), .A2(n589), .ZN(n564) );
  XNOR2_X1 U654 ( .A(KEYINPUT30), .B(n564), .ZN(n570) );
  NOR2_X1 U655 ( .A1(G900), .A2(n565), .ZN(n566) );
  NAND2_X1 U656 ( .A1(n566), .A2(n437), .ZN(n567) );
  NAND2_X1 U657 ( .A1(n568), .A2(n567), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n575), .B(KEYINPUT40), .ZN(n733) );
  INV_X1 U659 ( .A(n576), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n590), .A2(n592), .ZN(n579) );
  NOR2_X1 U661 ( .A1(n580), .A2(n579), .ZN(n582) );
  XOR2_X1 U662 ( .A(KEYINPUT28), .B(KEYINPUT107), .Z(n581) );
  XNOR2_X1 U663 ( .A(n582), .B(n581), .ZN(n583) );
  NAND2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n601) );
  NOR2_X1 U665 ( .A1(n601), .A2(n625), .ZN(n585) );
  XOR2_X1 U666 ( .A(KEYINPUT42), .B(n585), .Z(n734) );
  NAND2_X1 U667 ( .A1(n733), .A2(n734), .ZN(n587) );
  NAND2_X1 U668 ( .A1(n686), .A2(n591), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n594) );
  INV_X1 U670 ( .A(n596), .ZN(n619) );
  NAND2_X1 U671 ( .A1(n616), .A2(n619), .ZN(n597) );
  INV_X1 U672 ( .A(n599), .ZN(n600) );
  INV_X1 U673 ( .A(n602), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n683), .A2(n603), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT73), .B(n604), .Z(n605) );
  NOR2_X1 U676 ( .A1(n691), .A2(n605), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(KEYINPUT47), .ZN(n611) );
  AND2_X1 U678 ( .A1(n608), .A2(n619), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n682) );
  NAND2_X1 U680 ( .A1(n611), .A2(n682), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n614), .A2(n347), .ZN(n694) );
  NAND2_X1 U682 ( .A1(KEYINPUT2), .A2(n694), .ZN(n615) );
  XNOR2_X1 U683 ( .A(KEYINPUT79), .B(n615), .ZN(n621) );
  NAND2_X1 U684 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U685 ( .A(KEYINPUT43), .B(n618), .Z(n620) );
  OR2_X1 U686 ( .A1(n620), .A2(n619), .ZN(n638) );
  NAND2_X1 U687 ( .A1(n621), .A2(n638), .ZN(n622) );
  NOR2_X1 U688 ( .A1(n629), .A2(n622), .ZN(n630) );
  INV_X1 U689 ( .A(KEYINPUT2), .ZN(n623) );
  NOR2_X1 U690 ( .A1(n624), .A2(n623), .ZN(n627) );
  NOR2_X1 U691 ( .A1(n625), .A2(n524), .ZN(n626) );
  NAND2_X1 U692 ( .A1(n694), .A2(n638), .ZN(n628) );
  NOR2_X2 U693 ( .A1(n629), .A2(n628), .ZN(n724) );
  OR2_X1 U694 ( .A1(n639), .A2(n630), .ZN(n631) );
  NAND2_X1 U695 ( .A1(n633), .A2(n710), .ZN(n635) );
  XNOR2_X1 U696 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n634) );
  XOR2_X1 U697 ( .A(G119), .B(KEYINPUT127), .Z(n636) );
  XNOR2_X1 U698 ( .A(n637), .B(n636), .ZN(G21) );
  XNOR2_X1 U699 ( .A(n638), .B(G140), .ZN(G42) );
  INV_X1 U700 ( .A(n640), .ZN(n641) );
  NAND2_X1 U701 ( .A1(n641), .A2(KEYINPUT2), .ZN(n642) );
  XNOR2_X1 U702 ( .A(n642), .B(KEYINPUT66), .ZN(n643) );
  NAND2_X1 U703 ( .A1(n704), .A2(G210), .ZN(n649) );
  XOR2_X1 U704 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n646) );
  XNOR2_X1 U705 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U706 ( .A(n649), .B(n648), .ZN(n651) );
  INV_X1 U707 ( .A(G952), .ZN(n650) );
  INV_X1 U708 ( .A(n709), .ZN(n665) );
  NAND2_X1 U709 ( .A1(n651), .A2(n665), .ZN(n653) );
  INV_X1 U710 ( .A(KEYINPUT56), .ZN(n652) );
  XNOR2_X1 U711 ( .A(n653), .B(n652), .ZN(G51) );
  NAND2_X1 U712 ( .A1(n704), .A2(G472), .ZN(n656) );
  XOR2_X1 U713 ( .A(n654), .B(KEYINPUT62), .Z(n655) );
  XNOR2_X1 U714 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U715 ( .A1(n657), .A2(n665), .ZN(n659) );
  XNOR2_X1 U716 ( .A(KEYINPUT84), .B(KEYINPUT63), .ZN(n658) );
  XNOR2_X1 U717 ( .A(n659), .B(n658), .ZN(G57) );
  NOR2_X1 U718 ( .A1(n661), .A2(n660), .ZN(n664) );
  XOR2_X1 U719 ( .A(n662), .B(KEYINPUT59), .Z(n663) );
  XNOR2_X1 U720 ( .A(n664), .B(n663), .ZN(n666) );
  NAND2_X1 U721 ( .A1(n666), .A2(n665), .ZN(n668) );
  INV_X1 U722 ( .A(KEYINPUT60), .ZN(n667) );
  XNOR2_X1 U723 ( .A(n668), .B(n667), .ZN(G60) );
  XNOR2_X1 U724 ( .A(G101), .B(n669), .ZN(n670) );
  XNOR2_X1 U725 ( .A(n670), .B(KEYINPUT109), .ZN(G3) );
  NAND2_X1 U726 ( .A1(n686), .A2(n675), .ZN(n671) );
  XNOR2_X1 U727 ( .A(n671), .B(G104), .ZN(G6) );
  XOR2_X1 U728 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n673) );
  XNOR2_X1 U729 ( .A(G107), .B(KEYINPUT26), .ZN(n672) );
  XNOR2_X1 U730 ( .A(n673), .B(n672), .ZN(n674) );
  XOR2_X1 U731 ( .A(KEYINPUT110), .B(n674), .Z(n677) );
  NAND2_X1 U732 ( .A1(n675), .A2(n347), .ZN(n676) );
  XNOR2_X1 U733 ( .A(n677), .B(n676), .ZN(G9) );
  XOR2_X1 U734 ( .A(G110), .B(n678), .Z(G12) );
  XOR2_X1 U735 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n680) );
  NAND2_X1 U736 ( .A1(n683), .A2(n347), .ZN(n679) );
  XNOR2_X1 U737 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U738 ( .A(G128), .B(n681), .ZN(G30) );
  XNOR2_X1 U739 ( .A(G143), .B(n682), .ZN(G45) );
  XOR2_X1 U740 ( .A(G146), .B(KEYINPUT113), .Z(n685) );
  NAND2_X1 U741 ( .A1(n683), .A2(n686), .ZN(n684) );
  XNOR2_X1 U742 ( .A(n685), .B(n684), .ZN(G48) );
  NAND2_X1 U743 ( .A1(n686), .A2(n688), .ZN(n687) );
  XNOR2_X1 U744 ( .A(n687), .B(G113), .ZN(G15) );
  NAND2_X1 U745 ( .A1(n688), .A2(n347), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n689), .B(KEYINPUT114), .ZN(n690) );
  XNOR2_X1 U747 ( .A(G116), .B(n690), .ZN(G18) );
  XOR2_X1 U748 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n693) );
  XNOR2_X1 U749 ( .A(G125), .B(n691), .ZN(n692) );
  XNOR2_X1 U750 ( .A(n693), .B(n692), .ZN(G27) );
  XNOR2_X1 U751 ( .A(G134), .B(KEYINPUT116), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n695), .B(n694), .ZN(G36) );
  NAND2_X1 U753 ( .A1(n704), .A2(G469), .ZN(n699) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n696) );
  XNOR2_X1 U755 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U756 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U757 ( .A1(n709), .A2(n700), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n704), .A2(G478), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U760 ( .A1(n709), .A2(n703), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n704), .A2(G217), .ZN(n707) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(G66) );
  NAND2_X1 U763 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U764 ( .A1(G953), .A2(G224), .ZN(n712) );
  XNOR2_X1 U765 ( .A(KEYINPUT61), .B(n712), .ZN(n713) );
  NAND2_X1 U766 ( .A1(n713), .A2(G898), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n720) );
  XNOR2_X1 U768 ( .A(n716), .B(KEYINPUT125), .ZN(n718) );
  NAND2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U770 ( .A(n720), .B(n719), .Z(G69) );
  XOR2_X1 U771 ( .A(n722), .B(n721), .Z(n723) );
  XOR2_X1 U772 ( .A(KEYINPUT126), .B(n723), .Z(n727) );
  XOR2_X1 U773 ( .A(n727), .B(n724), .Z(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n731) );
  XNOR2_X1 U775 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XOR2_X1 U779 ( .A(G122), .B(n732), .Z(G24) );
  XNOR2_X1 U780 ( .A(n733), .B(G131), .ZN(G33) );
  XNOR2_X1 U781 ( .A(G137), .B(n734), .ZN(G39) );
endmodule

