//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n453), .B2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n465), .A3(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT69), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G137), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(G160));
  AND2_X1   g058(.A1(new_n480), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n486));
  OAI211_X1 g061(.A(G2105), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT72), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n485), .A2(new_n486), .B1(new_n488), .B2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n479), .B2(new_n494), .ZN(new_n495));
  OR3_X1    g070(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(new_n469), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(new_n474), .B2(G114), .ZN(new_n500));
  NOR2_X1   g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n487), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G126), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT73), .B1(new_n516), .B2(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(new_n514), .A3(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G543), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n517), .A2(new_n519), .B1(new_n516), .B2(G651), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(new_n512), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT75), .B(G88), .Z(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n515), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n515), .A2(new_n524), .A3(new_n528), .A4(KEYINPUT76), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n525), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n510), .A2(new_n511), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n535), .B1(new_n536), .B2(new_n522), .C1(new_n537), .C2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT77), .B(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n526), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n523), .A2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n538), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G651), .B1(new_n523), .B2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n526), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  XOR2_X1   g134(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n560));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n522), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n525), .A2(G91), .A3(new_n512), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n525), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n510), .B2(new_n511), .ZN(new_n570));
  AND2_X1   g145(.A1(G78), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n572), .ZN(G299));
  XNOR2_X1  g148(.A(new_n548), .B(KEYINPUT79), .ZN(G301));
  INV_X1    g149(.A(G166), .ZN(G303));
  OAI21_X1  g150(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n576));
  INV_X1    g151(.A(G49), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n525), .A2(new_n512), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI221_X1 g154(.A(new_n576), .B1(new_n522), .B2(new_n577), .C1(new_n578), .C2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n526), .A2(G86), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n523), .A2(G48), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n510), .B2(new_n511), .ZN(new_n584));
  AND2_X1   g159(.A1(G73), .A2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n581), .A2(new_n582), .A3(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(new_n514), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n526), .A2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n523), .A2(G47), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND3_X1  g171(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n578), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n597), .A2(new_n600), .B1(G54), .B2(new_n523), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n512), .A2(G66), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT81), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n548), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n610), .B2(new_n607), .ZN(G284));
  OAI21_X1  g186(.A(new_n608), .B1(new_n610), .B2(new_n607), .ZN(G321));
  NAND2_X1  g187(.A1(G299), .A2(new_n607), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G168), .B2(new_n607), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(G168), .B2(new_n607), .ZN(G280));
  INV_X1    g190(.A(new_n606), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  OR3_X1    g193(.A1(new_n606), .A2(KEYINPUT82), .A3(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT82), .B1(new_n606), .B2(G559), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g199(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2100), .Z(new_n628));
  INV_X1    g203(.A(G135), .ZN(new_n629));
  NOR2_X1   g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n631));
  OAI22_X1  g206(.A1(new_n479), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n488), .B2(G123), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n628), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2435), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2438), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2443), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2096), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n653), .B2(new_n654), .ZN(new_n660));
  AOI21_X1  g235(.A(KEYINPUT18), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n658), .B(new_n661), .Z(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n668), .B1(KEYINPUT20), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n671), .B(new_n672), .C1(KEYINPUT20), .C2(new_n670), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G35), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G162), .B2(new_n681), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT29), .B(G2090), .Z(new_n684));
  XOR2_X1   g259(.A(new_n683), .B(new_n684), .Z(new_n685));
  XOR2_X1   g260(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G34), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(G29), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G160), .B2(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G2084), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT95), .ZN(new_n691));
  NOR2_X1   g266(.A1(G29), .A2(G32), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n472), .A2(G105), .ZN(new_n693));
  INV_X1    g268(.A(G141), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n479), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n488), .B2(G129), .ZN(new_n696));
  NAND3_X1  g271(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT26), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n692), .B1(new_n701), .B2(G29), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT27), .B(G1996), .Z(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n681), .A2(G33), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT25), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n472), .A2(G103), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(G115), .A2(G2104), .ZN(new_n710));
  INV_X1    g285(.A(G127), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n469), .B2(new_n711), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n480), .A2(G139), .B1(new_n712), .B2(G2105), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n705), .B1(new_n715), .B2(new_n681), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n704), .B1(G2072), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n691), .B(new_n717), .C1(G2072), .C2(new_n716), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT96), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n488), .A2(G128), .ZN(new_n720));
  OR2_X1    g295(.A1(G104), .A2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT90), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n480), .A2(G140), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(new_n681), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n681), .A2(G26), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT28), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(KEYINPUT28), .B2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G2067), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(G171), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G5), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n681), .B1(new_n738), .B2(G28), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT97), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n738), .B2(G28), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n633), .B2(G29), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n736), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G11), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n689), .A2(G2084), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n556), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G1341), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(G4), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n616), .B2(new_n746), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G1348), .Z(new_n753));
  INV_X1    g328(.A(KEYINPUT23), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n746), .A2(G20), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n754), .B(new_n755), .C1(G299), .C2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT98), .B(G1956), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n748), .A2(G1341), .ZN(new_n761));
  NOR2_X1   g336(.A1(G168), .A2(new_n746), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n746), .B2(G21), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n681), .A2(G27), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G164), .B2(new_n681), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n702), .A2(new_n703), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n765), .A2(new_n766), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n750), .A2(new_n760), .A3(new_n761), .A4(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n719), .A2(new_n732), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n488), .A2(G119), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT85), .ZN(new_n776));
  OR2_X1    g351(.A1(G95), .A2(G2105), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n778));
  INV_X1    g353(.A(G131), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n776), .B(new_n778), .C1(new_n779), .C2(new_n479), .ZN(new_n780));
  MUX2_X1   g355(.A(G25), .B(new_n780), .S(G29), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT86), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT35), .B(G1991), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n746), .A2(G23), .ZN(new_n785));
  INV_X1    g360(.A(G288), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n746), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT33), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1976), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n790));
  INV_X1    g365(.A(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(G16), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n746), .A2(KEYINPUT89), .A3(G22), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n792), .B(new_n793), .C1(G166), .C2(new_n746), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G6), .B(G305), .S(G16), .Z(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT32), .B(G1981), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT88), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n797), .B(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n789), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n803));
  NOR2_X1   g378(.A1(G16), .A2(G24), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT87), .ZN(new_n805));
  XNOR2_X1  g380(.A(G290), .B(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n804), .B1(new_n806), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n802), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(KEYINPUT36), .B1(new_n784), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n810), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n813));
  INV_X1    g388(.A(new_n783), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n782), .B(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI211_X1 g391(.A(new_n685), .B(new_n774), .C1(new_n811), .C2(new_n816), .ZN(G311));
  AOI21_X1  g392(.A(new_n774), .B1(new_n816), .B2(new_n811), .ZN(new_n818));
  INV_X1    g393(.A(new_n685), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(G150));
  NAND2_X1  g395(.A1(G80), .A2(G543), .ZN(new_n821));
  INV_X1    g396(.A(G67), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n538), .B2(new_n822), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n823), .A2(G651), .B1(new_n523), .B2(G55), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT99), .B(G93), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n526), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n616), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n556), .A2(new_n827), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n555), .A2(new_n824), .A3(new_n826), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT39), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n831), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n829), .B1(new_n836), .B2(G860), .ZN(G145));
  XOR2_X1   g412(.A(new_n492), .B(new_n633), .Z(new_n838));
  INV_X1    g413(.A(G160), .ZN(new_n839));
  INV_X1    g414(.A(G142), .ZN(new_n840));
  NOR2_X1   g415(.A1(G106), .A2(G2105), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(new_n474), .B2(G118), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n479), .A2(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n488), .B2(G130), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n780), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n780), .A2(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n700), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n700), .B1(new_n845), .B2(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n839), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n851), .A2(G160), .A3(new_n847), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n726), .B(new_n505), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n714), .A2(KEYINPUT100), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n714), .A2(KEYINPUT100), .ZN(new_n855));
  INV_X1    g430(.A(new_n626), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n853), .B(new_n859), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n850), .A2(new_n852), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n850), .B2(new_n852), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n838), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  INV_X1    g439(.A(new_n860), .ZN(new_n865));
  AOI21_X1  g440(.A(G160), .B1(new_n851), .B2(new_n847), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n848), .A2(new_n839), .A3(new_n849), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n838), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n850), .A2(new_n852), .A3(new_n860), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n863), .A2(new_n864), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT40), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n863), .A2(new_n871), .A3(new_n874), .A4(new_n864), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(G395));
  NOR2_X1   g451(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n606), .B(G299), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n555), .B(new_n827), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n834), .A2(KEYINPUT101), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n621), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n882), .A2(new_n883), .A3(new_n620), .A4(new_n619), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n879), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n879), .A2(KEYINPUT41), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  INV_X1    g465(.A(G299), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n606), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n606), .B(new_n891), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(new_n890), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n889), .B1(new_n894), .B2(KEYINPUT41), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n886), .A3(new_n885), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n878), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n885), .A2(new_n886), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT103), .B1(new_n899), .B2(new_n895), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n877), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n877), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n896), .A2(new_n878), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n887), .B1(new_n899), .B2(new_n895), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n902), .B(new_n903), .C1(new_n904), .C2(new_n878), .ZN(new_n905));
  NAND2_X1  g480(.A1(G290), .A2(new_n786), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n594), .A2(G288), .A3(new_n595), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(G305), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(G166), .B(G305), .Z(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(KEYINPUT104), .A3(new_n908), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n901), .A2(new_n905), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n901), .B2(new_n905), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n827), .A2(new_n607), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(G295));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n921), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT106), .B1(new_n610), .B2(G286), .ZN(new_n925));
  NAND2_X1  g500(.A1(G171), .A2(G286), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(G301), .A2(new_n927), .A3(G168), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n834), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n925), .A2(new_n928), .A3(new_n880), .A4(new_n926), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(KEYINPUT107), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n933), .A3(new_n834), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n895), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(new_n893), .A3(new_n931), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n916), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n864), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n916), .B1(new_n935), .B2(new_n936), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n924), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n916), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n893), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT108), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n894), .A2(KEYINPUT41), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n944), .A2(new_n945), .B1(new_n930), .B2(new_n931), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n879), .B1(new_n932), .B2(new_n934), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(KEYINPUT43), .A3(new_n864), .A4(new_n937), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT44), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT43), .B1(new_n938), .B2(new_n939), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n948), .A2(new_n924), .A3(new_n864), .A4(new_n937), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(G397));
  XOR2_X1   g532(.A(KEYINPUT109), .B(G1384), .Z(new_n958));
  AOI21_X1  g533(.A(KEYINPUT45), .B1(new_n505), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n473), .A2(G40), .A3(new_n481), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n726), .B(G2067), .ZN(new_n964));
  INV_X1    g539(.A(G1996), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n700), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n967), .A2(KEYINPUT110), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n964), .A2(new_n966), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(KEYINPUT110), .A3(new_n962), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n780), .A2(new_n783), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n726), .A2(new_n731), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n963), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n970), .ZN(new_n975));
  INV_X1    g550(.A(new_n971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n780), .A2(new_n783), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n963), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n963), .A2(G290), .A3(G1986), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT48), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n975), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n962), .A2(new_n965), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT46), .Z(new_n983));
  NAND2_X1  g558(.A1(new_n964), .A2(new_n701), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n984), .B2(new_n962), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT47), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n974), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G2084), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n475), .B1(new_n465), .B2(G2104), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n466), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n991), .A2(G138), .A3(new_n474), .A4(new_n476), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n497), .B1(new_n992), .B2(KEYINPUT4), .ZN(new_n993));
  INV_X1    g568(.A(G126), .ZN(new_n994));
  OAI22_X1  g569(.A1(new_n487), .A2(new_n994), .B1(new_n501), .B2(new_n500), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n960), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n499), .B2(new_n504), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1000), .B(new_n989), .C1(new_n993), .C2(new_n995), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(KEYINPUT111), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n988), .B(new_n997), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n961), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT45), .B(new_n989), .C1(new_n993), .C2(new_n995), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n764), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G8), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G286), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1002), .B(KEYINPUT111), .ZN(new_n1013));
  INV_X1    g588(.A(G2090), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n997), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n960), .B1(new_n996), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1971), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1012), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n531), .A2(G8), .A3(new_n532), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1022), .B(KEYINPUT55), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n961), .B1(new_n999), .B2(new_n1000), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1002), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1027), .A2(G2090), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n1029), .B2(new_n1019), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1012), .B1(new_n961), .B2(new_n999), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(G288), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  INV_X1    g610(.A(G48), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n586), .B1(new_n1036), .B2(new_n522), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT112), .B(G86), .Z(new_n1038));
  NOR2_X1   g613(.A1(new_n578), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n581), .A2(new_n582), .A3(new_n1041), .A4(new_n586), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1042), .A3(KEYINPUT49), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1032), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1033), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1032), .B(new_n1048), .C1(new_n1033), .C2(G288), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1035), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1011), .A2(new_n1025), .A3(new_n1031), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT63), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1035), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(KEYINPUT114), .A3(new_n1011), .A4(new_n1031), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1050), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1054), .B1(new_n1059), .B2(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1050), .B(new_n1061), .C1(new_n1021), .C2(new_n1024), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(new_n1025), .A3(new_n1011), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1050), .A2(new_n1024), .A3(new_n1021), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1047), .A2(new_n1033), .A3(new_n786), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1042), .B(KEYINPUT113), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1032), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G286), .A2(G8), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT122), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1010), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1012), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT123), .B1(new_n1075), .B2(new_n1072), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(KEYINPUT51), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1009), .A2(new_n1072), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT123), .B(new_n1079), .C1(new_n1075), .C2(new_n1072), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .A4(KEYINPUT124), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1017), .A2(new_n769), .A3(new_n1006), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1085), .A2(KEYINPUT125), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(KEYINPUT125), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1013), .A2(new_n997), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n735), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1017), .A2(new_n769), .A3(new_n1018), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1088), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT62), .B(new_n610), .C1(new_n1089), .C2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1083), .A2(new_n1084), .A3(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1056), .A2(new_n1031), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1956), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(KEYINPUT116), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(KEYINPUT116), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT117), .Z(new_n1104));
  AND3_X1   g679(.A1(G299), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(G299), .B2(new_n1102), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1017), .A2(new_n1018), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1100), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1348), .B1(new_n1013), .B2(new_n997), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n961), .A2(new_n999), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(G2067), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1110), .B(new_n616), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1017), .A2(new_n1018), .A3(new_n1108), .ZN(new_n1116));
  AOI21_X1  g691(.A(G1956), .B1(new_n997), .B2(new_n1002), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1017), .A2(new_n965), .A3(new_n1018), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT118), .B(G1341), .Z(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT58), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1112), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n556), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT119), .B1(new_n1125), .B2(KEYINPUT120), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1127), .A3(new_n556), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(KEYINPUT59), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  OAI211_X1 g705(.A(KEYINPUT119), .B(new_n1130), .C1(new_n1125), .C2(KEYINPUT120), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1118), .A2(new_n1110), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT61), .B1(new_n1132), .B2(KEYINPUT121), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  AOI211_X1 g710(.A(new_n1134), .B(new_n1135), .C1(new_n1118), .C2(new_n1110), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1129), .B(new_n1131), .C1(new_n1133), .C2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT60), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n616), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1119), .B1(new_n1137), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1089), .A2(new_n1094), .A3(new_n610), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1090), .A2(new_n735), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n959), .A2(new_n1088), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1148), .A2(new_n769), .A3(new_n961), .A4(new_n1018), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n548), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT54), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n610), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1147), .A2(G301), .A3(new_n1149), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1145), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1152), .A2(KEYINPUT62), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1069), .B1(new_n1098), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n975), .A2(new_n978), .ZN(new_n1162));
  XNOR2_X1  g737(.A(G290), .B(new_n808), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n963), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n987), .B1(new_n1161), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g740(.A(G227), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n649), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g742(.A(new_n677), .B(new_n678), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1169), .A2(G319), .ZN(new_n1170));
  OAI21_X1  g744(.A(KEYINPUT126), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g745(.A1(G229), .A2(new_n462), .ZN(new_n1172));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n1173));
  NAND4_X1  g747(.A1(new_n1172), .A2(new_n1173), .A3(new_n649), .A4(new_n1167), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  AND3_X1   g749(.A1(new_n1175), .A2(new_n872), .A3(new_n954), .ZN(G308));
  NAND3_X1  g750(.A1(new_n1175), .A2(new_n872), .A3(new_n954), .ZN(G225));
endmodule


