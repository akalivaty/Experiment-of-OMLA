//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT31), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G228gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT79), .A2(G155gat), .A3(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(KEYINPUT2), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(KEYINPUT80), .ZN(new_n219));
  AND2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G155gat), .B(G162gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n212), .A2(new_n224), .A3(KEYINPUT2), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n219), .A2(new_n222), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n218), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(G211gat), .A2(G218gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(G211gat), .A2(G218gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G197gat), .A2(G204gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(G197gat), .B(G204gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n237), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n242), .A3(KEYINPUT76), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(new_n233), .C1(new_n236), .C2(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n218), .A2(new_n226), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT29), .B1(new_n238), .B2(new_n242), .ZN(new_n249));
  INV_X1    g048(.A(new_n227), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n209), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n243), .A2(new_n229), .A3(new_n245), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n248), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT83), .ZN(new_n258));
  INV_X1    g057(.A(new_n209), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n230), .B2(new_n246), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n257), .B2(new_n260), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n253), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G22gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n206), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n209), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n218), .A2(new_n226), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n254), .B2(new_n255), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT83), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n252), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G22gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n264), .A2(KEYINPUT84), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  AND4_X1   g076(.A1(KEYINPUT85), .A2(new_n275), .A3(new_n277), .A4(new_n206), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n205), .B1(new_n263), .B2(new_n274), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT85), .B1(new_n279), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n273), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n284), .B2(KEYINPUT26), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n289), .B2(KEYINPUT26), .ZN(new_n290));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT27), .B(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(KEYINPUT28), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n297));
  NOR2_X1   g096(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT66), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n298), .B1(new_n303), .B2(KEYINPUT27), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n297), .B1(new_n304), .B2(G190gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n296), .B1(new_n305), .B2(KEYINPUT68), .ZN(new_n306));
  INV_X1    g105(.A(new_n298), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT66), .B(G183gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT27), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT28), .B1(new_n310), .B2(new_n294), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n292), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT64), .B(G176gat), .Z(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(KEYINPUT23), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n291), .A2(KEYINPUT24), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n282), .B1(new_n284), .B2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n317), .A2(new_n322), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n286), .A2(KEYINPUT23), .A3(new_n288), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n325), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n300), .A2(new_n302), .A3(new_n294), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n321), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n321), .A3(KEYINPUT67), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n328), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n326), .B1(new_n334), .B2(new_n323), .ZN(new_n335));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n314), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(KEYINPUT29), .ZN(new_n339));
  INV_X1    g138(.A(new_n292), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n295), .B1(new_n311), .B2(new_n312), .ZN(new_n341));
  AOI211_X1 g140(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n310), .C2(new_n294), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AND4_X1   g142(.A1(new_n323), .A2(new_n317), .A3(new_n322), .A4(new_n325), .ZN(new_n344));
  INV_X1    g143(.A(new_n333), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT67), .B1(new_n329), .B2(new_n321), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n325), .B(new_n327), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n344), .B1(new_n347), .B2(KEYINPUT25), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n339), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n246), .B1(new_n338), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n351));
  OAI22_X1  g150(.A1(new_n314), .A2(new_n335), .B1(KEYINPUT29), .B2(new_n337), .ZN(new_n352));
  INV_X1    g151(.A(new_n246), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n348), .A3(new_n336), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n352), .A2(KEYINPUT77), .A3(new_n353), .A4(new_n354), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G64gat), .ZN(new_n360));
  INV_X1    g159(.A(G92gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(KEYINPUT30), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n358), .A2(new_n362), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n358), .A2(new_n369), .A3(new_n362), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n366), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G113gat), .ZN(new_n374));
  INV_X1    g173(.A(G120gat), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT1), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G113gat), .A2(G120gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G127gat), .B(G134gat), .Z(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT69), .B(G134gat), .Z(new_n381));
  INV_X1    g180(.A(G127gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT70), .B(G127gat), .ZN(new_n383));
  INV_X1    g182(.A(G134gat), .ZN(new_n384));
  OAI22_X1  g183(.A1(new_n381), .A2(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n380), .B1(new_n385), .B2(new_n378), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n228), .C1(new_n255), .C2(new_n267), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n267), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n389), .A2(KEYINPUT4), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n386), .B2(new_n267), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n388), .B(new_n392), .C1(new_n393), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT5), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n385), .A2(new_n378), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n248), .B1(new_n398), .B2(new_n380), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n389), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n400), .B2(new_n391), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n389), .B(KEYINPUT4), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n391), .A2(KEYINPUT5), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n388), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT82), .B(KEYINPUT0), .Z(new_n406));
  XNOR2_X1  g205(.A(G1gat), .B(G29gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G57gat), .B(G85gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n402), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n402), .A2(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(new_n410), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n413), .B(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n281), .B1(new_n373), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n390), .B1(new_n403), .B2(new_n388), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT39), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n390), .A3(new_n389), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n423), .B2(KEYINPUT87), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(KEYINPUT87), .B2(new_n423), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n422), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT40), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n416), .A2(KEYINPUT40), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n369), .B1(new_n358), .B2(new_n362), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT78), .B(new_n364), .C1(new_n356), .C2(new_n357), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n372), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n363), .A2(new_n365), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n281), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n413), .B(new_n416), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n431), .B2(new_n432), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT38), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n362), .B1(new_n358), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n356), .A2(KEYINPUT37), .A3(new_n357), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT88), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n350), .A2(new_n355), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT38), .B1(new_n449), .B2(KEYINPUT37), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n444), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n448), .B1(new_n444), .B2(new_n450), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n439), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n419), .B1(new_n438), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  INV_X1    g255(.A(G227gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(new_n208), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n314), .A2(new_n386), .A3(new_n335), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n387), .B1(new_n343), .B2(new_n348), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n456), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT74), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT34), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n386), .B1(new_n314), .B2(new_n335), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n343), .A2(new_n387), .A3(new_n348), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n458), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT74), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n456), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n463), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(new_n458), .A3(new_n467), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G43gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT71), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(G71gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G99gat), .ZN(new_n476));
  INV_X1    g275(.A(G71gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n474), .B(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G99gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT73), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT33), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n481), .A2(KEYINPUT73), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT32), .B(new_n472), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT32), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT33), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n487), .B1(new_n490), .B2(new_n482), .ZN(new_n491));
  AOI211_X1 g290(.A(KEYINPUT72), .B(new_n481), .C1(new_n472), .C2(new_n489), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n471), .B(new_n486), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n486), .B1(new_n491), .B2(new_n492), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n463), .A2(new_n470), .A3(new_n465), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT75), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(KEYINPUT75), .A3(new_n495), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT36), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n281), .A2(new_n493), .A3(new_n496), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n373), .A2(new_n504), .A3(new_n418), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n436), .A2(new_n437), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n418), .A2(new_n508), .A3(new_n281), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n500), .B2(new_n498), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n455), .A2(new_n503), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT91), .B(KEYINPUT17), .ZN(new_n513));
  XOR2_X1   g312(.A(G43gat), .B(G50gat), .Z(new_n514));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT89), .B(G29gat), .Z(new_n518));
  OR3_X1    g317(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n518), .A2(G36gat), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n514), .B2(new_n515), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n517), .B1(new_n521), .B2(new_n523), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n513), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT16), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(G1gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G15gat), .B(G22gat), .Z(new_n533));
  INV_X1    g332(.A(G1gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n528), .B(KEYINPUT92), .C1(new_n529), .C2(G1gat), .ZN(new_n536));
  XOR2_X1   g335(.A(KEYINPUT93), .B(G8gat), .Z(new_n537));
  NAND4_X1  g336(.A1(new_n532), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n530), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G8gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT94), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n521), .A2(new_n523), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(KEYINPUT17), .A3(new_n524), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n538), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n527), .A2(new_n542), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n524), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n541), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n548), .A2(KEYINPUT18), .A3(new_n549), .A4(new_n551), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n550), .B(new_n541), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n549), .B(KEYINPUT13), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G113gat), .B(G141gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT11), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G169gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G197gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(new_n316), .ZN(new_n564));
  INV_X1    g363(.A(G197gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n563), .A2(new_n566), .A3(KEYINPUT12), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT12), .B1(new_n563), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n552), .A2(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(new_n569), .A3(new_n555), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT97), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT41), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n361), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n587), .A2(new_n588), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n587), .A2(KEYINPUT99), .A3(new_n588), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n581), .B1(new_n596), .B2(new_n550), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n527), .A2(new_n545), .A3(new_n595), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n577), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n577), .A3(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n580), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n599), .B2(KEYINPUT100), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G71gat), .B(G78gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT9), .ZN(new_n613));
  INV_X1    g412(.A(G78gat), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n613), .B1(new_n477), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G57gat), .B(G64gat), .Z(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT21), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n538), .B(new_n540), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT96), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT95), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n623), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n621), .ZN(new_n629));
  XOR2_X1   g428(.A(G127gat), .B(G155gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n628), .B(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n610), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G230gat), .A2(G233gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n595), .A2(new_n620), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  INV_X1    g438(.A(new_n588), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n587), .A2(KEYINPUT101), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n583), .A2(new_n642), .A3(new_n586), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n640), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT102), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n620), .A2(new_n592), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n644), .B2(KEYINPUT102), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n638), .B(new_n639), .C1(new_n646), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n591), .A2(new_n594), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n620), .A2(new_n592), .A3(new_n639), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n637), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n638), .B1(new_n646), .B2(new_n648), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n655), .A2(new_n637), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT103), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n654), .A2(new_n656), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n654), .B2(new_n656), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n635), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n512), .A2(new_n575), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n440), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  INV_X1    g468(.A(new_n507), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(G8gat), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND3_X1  g473(.A1(new_n667), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n675), .A2(KEYINPUT104), .A3(new_n673), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT104), .B1(new_n675), .B2(new_n673), .ZN(new_n677));
  OAI221_X1 g476(.A(new_n672), .B1(new_n673), .B2(new_n675), .C1(new_n676), .C2(new_n677), .ZN(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n498), .A2(new_n500), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n667), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n503), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n501), .A2(KEYINPUT105), .A3(new_n502), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n667), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n681), .B1(new_n686), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n667), .A2(new_n439), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n512), .A2(new_n575), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n665), .A2(new_n634), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n609), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT106), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(new_n418), .A3(new_n518), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT45), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT44), .B1(new_n512), .B2(new_n609), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n511), .A2(new_n506), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n373), .A2(new_n418), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n439), .ZN(new_n701));
  INV_X1    g500(.A(new_n430), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT30), .B1(new_n368), .B2(new_n370), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT86), .B1(new_n703), .B2(new_n366), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n444), .A2(new_n445), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT38), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n440), .A3(new_n371), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n444), .A2(new_n450), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT88), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n444), .A2(new_n448), .A3(new_n450), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n281), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n701), .B1(new_n706), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n699), .B1(new_n685), .B2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n610), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n698), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n692), .A2(new_n575), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n518), .B1(new_n723), .B2(new_n418), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n696), .A2(KEYINPUT45), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n697), .A2(new_n724), .A3(new_n725), .ZN(G1328gat));
  OAI21_X1  g525(.A(G36gat), .B1(new_n723), .B2(new_n507), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n507), .A2(G36gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n695), .A2(KEYINPUT108), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT108), .B1(new_n695), .B2(new_n729), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n730), .B2(new_n732), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(G1329gat));
  NAND3_X1  g534(.A1(new_n721), .A2(new_n685), .A3(new_n722), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G43gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n680), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n695), .A2(G43gat), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n737), .A2(new_n739), .A3(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1330gat));
  NAND3_X1  g543(.A1(new_n721), .A2(new_n439), .A3(new_n722), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n691), .A2(new_n204), .A3(new_n439), .A4(new_n694), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT48), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1331gat));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n507), .A2(new_n510), .B1(new_n505), .B2(KEYINPUT35), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n501), .A2(KEYINPUT105), .A3(new_n502), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT105), .B1(new_n501), .B2(new_n502), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(new_n455), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n635), .A2(new_n575), .A3(new_n664), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n753), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n759), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n716), .A2(KEYINPUT109), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n418), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT110), .B(G57gat), .Z(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1332gat));
  OAI22_X1  g565(.A1(new_n763), .A2(new_n507), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT49), .B(G64gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n760), .A2(new_n762), .A3(new_n670), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n763), .B2(new_n757), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n680), .A2(new_n477), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n763), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n771), .B(KEYINPUT50), .C1(new_n763), .C2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1334gat));
  NOR2_X1   g576(.A1(new_n763), .A2(new_n281), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT111), .B(G78gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1335gat));
  NAND2_X1  g579(.A1(new_n575), .A2(new_n634), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT112), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n664), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n698), .B2(new_n720), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(G85gat), .B1(new_n785), .B2(new_n418), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n610), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT51), .B1(new_n758), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  INV_X1    g588(.A(new_n787), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n716), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n791), .A3(new_n664), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n440), .A2(new_n585), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n786), .B1(new_n792), .B2(new_n793), .ZN(G1336gat));
  INV_X1    g593(.A(new_n783), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n501), .A2(new_n502), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n699), .B1(new_n715), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n610), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n758), .A2(new_n718), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n670), .B(new_n795), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n507), .A2(G92gat), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n791), .A3(new_n664), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT52), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n802), .A2(new_n803), .A3(new_n808), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1337gat));
  OAI21_X1  g609(.A(new_n479), .B1(new_n792), .B2(new_n738), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n685), .A2(G99gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n785), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n811), .B(KEYINPUT114), .C1(new_n785), .C2(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1338gat));
  OAI211_X1 g616(.A(new_n439), .B(new_n795), .C1(new_n799), .C2(new_n800), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G106gat), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n281), .A2(G106gat), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n788), .A2(new_n791), .A3(new_n664), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  XOR2_X1   g623(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(new_n819), .ZN(new_n828));
  INV_X1    g627(.A(G106gat), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n829), .B1(new_n784), .B2(new_n439), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n826), .A3(KEYINPUT116), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n823), .B1(new_n828), .B2(new_n831), .ZN(G1339gat));
  NOR2_X1   g631(.A1(new_n666), .A2(new_n574), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n563), .A2(new_n566), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n549), .B1(new_n548), .B2(new_n551), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n556), .A2(new_n557), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n573), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT117), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n636), .B1(new_n651), .B2(new_n652), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n649), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n649), .A2(new_n653), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n637), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n660), .B1(new_n654), .B2(new_n840), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT55), .ZN(new_n846));
  AND4_X1   g645(.A1(new_n607), .A2(new_n846), .A3(new_n608), .A4(new_n662), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT55), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n839), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n573), .A2(new_n837), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n664), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT118), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n849), .A2(new_n574), .A3(new_n662), .A4(new_n846), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n664), .A3(new_n855), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n850), .B1(new_n857), .B2(new_n610), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n833), .B1(new_n858), .B2(new_n634), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(new_n439), .A3(new_n738), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n440), .A3(new_n507), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(new_n374), .A3(new_n575), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n859), .A2(new_n418), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n507), .A2(new_n504), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n574), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n862), .A2(new_n867), .ZN(G1340gat));
  NOR3_X1   g667(.A1(new_n861), .A2(new_n375), .A3(new_n665), .ZN(new_n869));
  AOI21_X1  g668(.A(G120gat), .B1(new_n866), .B2(new_n664), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(G1341gat));
  OAI21_X1  g670(.A(new_n383), .B1(new_n861), .B2(new_n634), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n634), .A2(new_n383), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n865), .B2(new_n873), .ZN(G1342gat));
  OR3_X1    g673(.A1(new_n865), .A2(new_n381), .A3(new_n609), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n861), .B2(new_n609), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G1343gat));
  INV_X1    g678(.A(new_n634), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  AND4_X1   g680(.A1(new_n569), .A2(new_n554), .A3(new_n555), .A4(new_n558), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n569), .B1(new_n572), .B2(new_n555), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n662), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT55), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(new_n848), .ZN(new_n886));
  INV_X1    g685(.A(new_n852), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n574), .A2(new_n662), .A3(new_n846), .ZN(new_n889));
  OAI211_X1 g688(.A(KEYINPUT119), .B(new_n852), .C1(new_n889), .C2(new_n848), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n609), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n880), .B1(new_n891), .B2(new_n850), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n439), .B1(new_n892), .B2(new_n833), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(new_n859), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n281), .A2(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n685), .A2(new_n418), .A3(new_n670), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G141gat), .B1(new_n899), .B2(new_n575), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n859), .A2(KEYINPUT120), .A3(new_n418), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT120), .B1(new_n859), .B2(new_n418), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n685), .A2(new_n670), .A3(new_n281), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n575), .A2(G141gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n908), .B(G148gat), .C1(new_n899), .C2(new_n665), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n892), .B2(new_n833), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n890), .A2(new_n609), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT119), .B1(new_n854), .B2(new_n852), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n850), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n634), .ZN(new_n916));
  INV_X1    g715(.A(new_n833), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(KEYINPUT121), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n912), .A2(new_n918), .A3(new_n896), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT57), .B1(new_n859), .B2(new_n281), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n919), .A2(new_n664), .A3(new_n898), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G148gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n910), .B1(new_n922), .B2(KEYINPUT59), .ZN(new_n923));
  AOI211_X1 g722(.A(KEYINPUT122), .B(new_n908), .C1(new_n921), .C2(G148gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n909), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OR3_X1    g724(.A1(new_n904), .A2(G148gat), .A3(new_n665), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1345gat));
  INV_X1    g726(.A(new_n904), .ZN(new_n928));
  AOI21_X1  g727(.A(G155gat), .B1(new_n928), .B2(new_n880), .ZN(new_n929));
  INV_X1    g728(.A(new_n899), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n880), .A2(G155gat), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT123), .Z(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n930), .B2(new_n932), .ZN(G1346gat));
  OAI21_X1  g732(.A(G162gat), .B1(new_n899), .B2(new_n609), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n609), .A2(G162gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n904), .B2(new_n935), .ZN(G1347gat));
  NAND2_X1  g735(.A1(new_n670), .A2(new_n418), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n860), .A2(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n316), .A3(new_n575), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n895), .A2(new_n504), .A3(new_n938), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n574), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n316), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT124), .ZN(G1348gat));
  NOR3_X1   g743(.A1(new_n939), .A2(new_n315), .A3(new_n665), .ZN(new_n945));
  AOI21_X1  g744(.A(G176gat), .B1(new_n941), .B2(new_n664), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(new_n303), .B1(new_n939), .B2(new_n634), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n941), .A2(new_n293), .A3(new_n880), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n941), .A2(new_n294), .A3(new_n610), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n860), .A2(new_n610), .A3(new_n938), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G190gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n953), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n955), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n952), .B1(new_n959), .B2(new_n960), .ZN(G1351gat));
  NAND2_X1  g760(.A1(new_n895), .A2(new_n439), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n938), .A2(new_n757), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n574), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n963), .B(KEYINPUT126), .Z(new_n966));
  NOR3_X1   g765(.A1(new_n966), .A2(new_n565), .A3(new_n575), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n919), .A2(new_n920), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G1352gat));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n664), .ZN(new_n970));
  OAI21_X1  g769(.A(G204gat), .B1(new_n970), .B2(new_n966), .ZN(new_n971));
  NOR4_X1   g770(.A1(new_n962), .A2(new_n963), .A3(G204gat), .A4(new_n665), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(G1353gat));
  NOR2_X1   g775(.A1(new_n963), .A2(new_n634), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n919), .A3(new_n920), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n962), .A2(G211gat), .ZN(new_n981));
  AOI22_X1  g780(.A1(new_n979), .A2(new_n980), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n979), .A2(new_n980), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  AOI21_X1  g784(.A(G218gat), .B1(new_n964), .B2(new_n610), .ZN(new_n986));
  INV_X1    g785(.A(G218gat), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n966), .A2(new_n987), .A3(new_n609), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n986), .B1(new_n988), .B2(new_n968), .ZN(G1355gat));
endmodule


