//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n197), .A3(new_n201), .A4(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n206), .B(new_n208), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(G107), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G104), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n206), .A2(new_n208), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n219), .A2(G104), .ZN(new_n226));
  OAI21_X1  g040(.A(G101), .B1(new_n212), .B2(new_n226), .ZN(new_n227));
  AND4_X1   g041(.A1(new_n210), .A2(new_n222), .A3(new_n225), .A4(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT10), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT0), .A4(G128), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n206), .A2(new_n208), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G128), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n215), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n217), .B1(new_n212), .B2(new_n214), .ZN(new_n237));
  OAI21_X1  g051(.A(G101), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n235), .B1(new_n238), .B2(KEYINPUT4), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n226), .B1(new_n220), .B2(new_n218), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n216), .B1(new_n242), .B2(new_n215), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n240), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n238), .A2(KEYINPUT82), .A3(KEYINPUT4), .A4(new_n222), .ZN(new_n245));
  AOI211_X1 g059(.A(KEYINPUT83), .B(new_n239), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n245), .ZN(new_n248));
  INV_X1    g062(.A(new_n239), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n204), .B(new_n230), .C1(new_n246), .C2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G140), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n253), .A2(G227), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n230), .B1(new_n246), .B2(new_n250), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n203), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n225), .A2(new_n210), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n222), .B2(new_n227), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n203), .B1(new_n262), .B2(new_n228), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT12), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n251), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n257), .A2(new_n259), .B1(new_n266), .B2(new_n255), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n192), .B1(new_n267), .B2(G469), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n256), .B1(new_n259), .B2(new_n251), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n251), .A2(new_n265), .A3(new_n256), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n190), .B(new_n191), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n189), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G214), .B1(G237), .B2(G902), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT84), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT71), .B(G125), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n225), .A2(new_n210), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G125), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT71), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G125), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n231), .B(new_n281), .C1(new_n232), .C2(new_n233), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n253), .A2(G224), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT2), .B(G113), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(G116), .B(G119), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g104(.A(G116), .B(G119), .Z(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n287), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(new_n238), .B2(KEYINPUT4), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n244), .B2(new_n245), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n296));
  INV_X1    g110(.A(G119), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(G116), .ZN(new_n298));
  OAI211_X1 g112(.A(G113), .B(new_n298), .C1(new_n291), .C2(new_n296), .ZN(new_n299));
  AND4_X1   g113(.A1(new_n290), .A2(new_n299), .A3(new_n222), .A4(new_n227), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n286), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(G110), .B(G122), .Z(new_n302));
  AND2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n294), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n300), .B1(new_n248), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT85), .ZN(new_n306));
  INV_X1    g120(.A(new_n302), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n303), .A2(new_n306), .B1(KEYINPUT6), .B2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n306), .A2(KEYINPUT6), .A3(new_n301), .A4(new_n302), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n285), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G210), .B1(G237), .B2(G902), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n295), .A2(new_n300), .A3(new_n302), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n302), .B(new_n315), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n290), .A2(new_n299), .B1(new_n222), .B2(new_n227), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n300), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n284), .A2(KEYINPUT7), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n276), .A2(new_n282), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n319), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT87), .B1(new_n283), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n283), .A2(KEYINPUT87), .A3(new_n321), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n318), .B(new_n320), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n191), .B1(new_n314), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(KEYINPUT88), .B(new_n191), .C1(new_n314), .C2(new_n324), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n312), .A2(new_n313), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n313), .ZN(new_n331));
  INV_X1    g145(.A(new_n285), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n306), .A2(new_n302), .A3(new_n301), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n308), .A2(KEYINPUT6), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n332), .B1(new_n335), .B2(new_n310), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n328), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n274), .B1(new_n330), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n272), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT16), .ZN(new_n342));
  INV_X1    g156(.A(G140), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n281), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n278), .B2(new_n280), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n277), .A2(new_n343), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n345), .B(KEYINPUT16), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n347), .B1(new_n275), .B2(new_n343), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n345), .B1(new_n351), .B2(KEYINPUT16), .ZN(new_n352));
  OAI211_X1 g166(.A(G146), .B(new_n344), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n348), .B1(new_n281), .B2(G140), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT72), .B1(new_n355), .B2(new_n342), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n349), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G146), .A4(new_n344), .ZN(new_n359));
  INV_X1    g173(.A(G237), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n253), .A3(G214), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(new_n207), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G131), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n361), .B(G143), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n201), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT19), .ZN(new_n367));
  NAND2_X1  g181(.A1(G125), .A2(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n347), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT76), .B1(new_n347), .B2(new_n368), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n355), .A2(KEYINPUT19), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n205), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n354), .A2(new_n359), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n371), .A2(new_n372), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n378), .A2(KEYINPUT77), .A3(G146), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT77), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n369), .B(new_n370), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(new_n205), .ZN(new_n382));
  OAI22_X1  g196(.A1(new_n379), .A2(new_n382), .B1(new_n205), .B2(new_n351), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT18), .A2(G131), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n362), .B(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n377), .A2(KEYINPUT90), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT90), .B1(new_n377), .B2(new_n386), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n341), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT73), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n353), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n357), .A2(KEYINPUT73), .A3(G146), .A4(new_n344), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n344), .B1(new_n350), .B2(new_n352), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n205), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n362), .A2(KEYINPUT17), .A3(G131), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n366), .B2(KEYINPUT17), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n386), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n401), .A2(new_n389), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n377), .A2(new_n386), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n405), .A2(KEYINPUT91), .A3(new_n389), .A4(new_n387), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n392), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT92), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n409), .A2(KEYINPUT20), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n401), .B(new_n389), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n191), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G475), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT94), .B(KEYINPUT13), .Z(new_n421));
  NAND2_X1  g235(.A1(new_n209), .A2(G143), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n209), .A2(G143), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n194), .B1(new_n426), .B2(KEYINPUT95), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT95), .ZN(new_n428));
  INV_X1    g242(.A(new_n425), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n427), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n422), .A3(new_n194), .ZN(new_n432));
  INV_X1    g246(.A(G116), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G122), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT93), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(G122), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(G107), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n431), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n440), .B(KEYINPUT96), .Z(new_n441));
  OAI21_X1  g255(.A(new_n435), .B1(KEYINPUT14), .B2(new_n436), .ZN(new_n442));
  OAI21_X1  g256(.A(G107), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G134), .B1(new_n423), .B2(new_n425), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n432), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n443), .B(new_n445), .C1(G107), .C2(new_n437), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G217), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n187), .A2(new_n448), .A3(G953), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n447), .B(new_n449), .Z(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n191), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT97), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(KEYINPUT15), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(KEYINPUT15), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n451), .B(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G952), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n459), .A2(KEYINPUT98), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(KEYINPUT98), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n253), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(G234), .A2(G237), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(G902), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n458), .A2(new_n470), .ZN(new_n471));
  AND4_X1   g285(.A1(new_n340), .A2(new_n417), .A3(new_n420), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n448), .B1(G234), .B2(new_n191), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n379), .A2(new_n382), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n297), .A2(G128), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n297), .A2(G128), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n478), .B(new_n479), .C1(new_n480), .C2(KEYINPUT23), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT24), .B(G110), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n209), .A2(G119), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n484), .A2(new_n478), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n481), .A2(G110), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n477), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n354), .A2(new_n359), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n481), .A2(G110), .B1(new_n483), .B2(new_n485), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n398), .A2(KEYINPUT74), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT74), .B1(new_n398), .B2(new_n490), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT78), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n495), .B(new_n489), .C1(new_n491), .C2(new_n492), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT79), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT22), .B(G137), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n492), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n398), .A2(KEYINPUT74), .A3(new_n490), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n503), .A2(new_n504), .B1(new_n488), .B2(new_n487), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n505), .B2(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n476), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n502), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n474), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT65), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n194), .B2(G137), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n196), .A2(KEYINPUT65), .A3(G134), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n198), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G131), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n261), .A2(KEYINPUT66), .A3(new_n202), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT64), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n231), .B(new_n520), .C1(new_n232), .C2(new_n233), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n203), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT66), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n202), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n523), .B1(new_n524), .B2(new_n260), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT67), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n260), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n529), .B2(new_n524), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n235), .A2(new_n203), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(KEYINPUT30), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(new_n533), .A3(new_n293), .ZN(new_n534));
  INV_X1    g348(.A(new_n293), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n360), .A2(new_n253), .A3(G210), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n538), .B(KEYINPUT27), .Z(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT26), .B(G101), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n539), .B(new_n540), .Z(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n537), .A2(new_n542), .B1(KEYINPUT68), .B2(KEYINPUT31), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n526), .A2(new_n293), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n536), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n542), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT68), .B(KEYINPUT31), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n534), .A2(new_n541), .A3(new_n536), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n543), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(G472), .A2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT32), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n537), .A2(new_n541), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT29), .ZN(new_n558));
  AOI21_X1  g372(.A(G902), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n545), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n531), .A2(new_n532), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n293), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(KEYINPUT69), .B2(new_n536), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n536), .A2(KEYINPUT69), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT28), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n558), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n545), .A2(new_n547), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n541), .B1(new_n568), .B2(KEYINPUT29), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n559), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n554), .A2(new_n556), .B1(new_n570), .B2(G472), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n505), .A2(new_n500), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n473), .A2(G902), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n502), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n512), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n472), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  INV_X1    g391(.A(new_n470), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n551), .A2(new_n191), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(G472), .B1(new_n551), .B2(new_n552), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n272), .A2(new_n339), .A3(new_n578), .A4(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n512), .A2(new_n581), .A3(new_n574), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(KEYINPUT99), .ZN(new_n585));
  MUX2_X1   g399(.A(new_n583), .B(new_n585), .S(new_n450), .Z(new_n586));
  NOR2_X1   g400(.A1(new_n452), .A2(G902), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT100), .B(G478), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n586), .A2(new_n587), .B1(new_n451), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n417), .B2(new_n420), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT34), .B(G104), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT101), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(G6));
  NAND3_X1  g408(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n413), .A2(new_n415), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n420), .ZN(new_n597));
  INV_X1    g411(.A(new_n458), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n582), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G107), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  INV_X1    g417(.A(new_n573), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n501), .A2(KEYINPUT36), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n494), .B2(new_n496), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n494), .A2(new_n496), .A3(new_n605), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT103), .B1(new_n512), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n611));
  INV_X1    g425(.A(new_n609), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n502), .A2(new_n506), .A3(new_n510), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n510), .B1(new_n502), .B2(new_n506), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n613), .A2(new_n614), .A3(new_n476), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n611), .B(new_n612), .C1(new_n615), .C2(new_n474), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n420), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n414), .B1(new_n409), .B2(new_n411), .ZN(new_n619));
  AOI211_X1 g433(.A(KEYINPUT92), .B(new_n410), .C1(new_n407), .C2(new_n408), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n618), .B1(new_n621), .B2(new_n416), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n622), .A2(new_n340), .A3(new_n471), .A4(new_n580), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT37), .B(G110), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G12));
  NAND2_X1  g440(.A1(new_n507), .A2(new_n508), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n511), .A3(new_n475), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n473), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n611), .B1(new_n629), .B2(new_n612), .ZN(new_n630));
  AOI211_X1 g444(.A(KEYINPUT103), .B(new_n609), .C1(new_n628), .C2(new_n473), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n571), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n465), .B1(G900), .B2(new_n468), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT104), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n597), .A2(new_n598), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n632), .A2(new_n633), .A3(new_n340), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  AOI21_X1  g452(.A(new_n313), .B1(new_n312), .B2(new_n329), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n336), .A2(new_n337), .A3(new_n331), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT38), .Z(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n564), .A2(new_n565), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n191), .B1(new_n644), .B2(new_n541), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n542), .B1(new_n534), .B2(new_n536), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n554), .A2(new_n556), .B1(new_n647), .B2(G472), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n643), .A2(new_n274), .A3(new_n598), .A4(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n622), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n512), .A2(new_n609), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n635), .B(KEYINPUT39), .Z(new_n652));
  NAND2_X1  g466(.A1(new_n272), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT40), .Z(new_n654));
  NAND4_X1  g468(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  INV_X1    g470(.A(new_n589), .ZN(new_n657));
  INV_X1    g471(.A(new_n635), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n409), .A2(KEYINPUT20), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n619), .A2(new_n620), .A3(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n657), .B(new_n658), .C1(new_n660), .C2(new_n618), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n632), .A2(new_n633), .A3(new_n340), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G146), .ZN(G48));
  OR2_X1    g478(.A1(new_n269), .A2(new_n270), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n190), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n191), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n191), .B1(new_n269), .B2(new_n270), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n667), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n669), .A2(new_n188), .A3(new_n671), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n512), .A2(new_n571), .A3(new_n574), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n274), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n639), .B2(new_n640), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n470), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n590), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT41), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G113), .ZN(G15));
  NAND3_X1  g493(.A1(new_n673), .A2(new_n599), .A3(new_n676), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  NOR2_X1   g495(.A1(new_n672), .A2(new_n675), .ZN(new_n682));
  AND4_X1   g496(.A1(new_n417), .A2(new_n682), .A3(new_n420), .A4(new_n471), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n633), .A3(new_n610), .A4(new_n616), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  NOR2_X1   g499(.A1(new_n622), .A2(new_n598), .ZN(new_n686));
  INV_X1    g500(.A(new_n672), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n676), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n512), .B2(new_n574), .ZN(new_n691));
  INV_X1    g505(.A(new_n574), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n692), .B(KEYINPUT107), .C1(new_n615), .C2(new_n474), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n579), .A2(G472), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n552), .B(KEYINPUT106), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n541), .B1(new_n561), .B2(new_n566), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n543), .A2(new_n550), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT108), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n703), .B(new_n700), .C1(new_n691), .C2(new_n693), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n689), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n661), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n590), .A2(KEYINPUT109), .A3(new_n658), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n651), .A2(new_n700), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n682), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  AOI21_X1  g526(.A(new_n574), .B1(new_n628), .B2(new_n473), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n641), .A2(new_n674), .ZN(new_n714));
  INV_X1    g528(.A(new_n272), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n713), .A2(new_n633), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n708), .A2(new_n717), .A3(new_n709), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n571), .B1(new_n691), .B2(new_n693), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n714), .A2(new_n715), .A3(new_n719), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n708), .A3(new_n709), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G131), .ZN(G33));
  NAND2_X1  g539(.A1(new_n717), .A2(new_n636), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT110), .B(G134), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G36));
  NAND2_X1  g542(.A1(new_n622), .A2(new_n657), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT112), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n622), .A2(KEYINPUT43), .A3(new_n657), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n734), .A3(new_n730), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n651), .A2(new_n580), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(KEYINPUT44), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n267), .B2(KEYINPUT45), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(KEYINPUT45), .B2(new_n267), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n192), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n271), .B1(new_n741), .B2(KEYINPUT46), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n188), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n714), .B(KEYINPUT113), .Z(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n652), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n738), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT44), .B1(new_n736), .B2(new_n737), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G137), .ZN(G39));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n754));
  XOR2_X1   g568(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n755));
  MUX2_X1   g569(.A(new_n754), .B(new_n755), .S(new_n744), .Z(new_n756));
  OR4_X1    g570(.A1(new_n633), .A2(new_n661), .A3(new_n713), .A4(new_n714), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  NAND3_X1  g573(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n597), .A2(new_n458), .A3(new_n635), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n633), .A3(new_n610), .A4(new_n616), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n716), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n724), .A3(new_n726), .ZN(new_n765));
  INV_X1    g579(.A(new_n581), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n713), .A2(new_n622), .A3(new_n766), .A4(new_n458), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n617), .B2(new_n623), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(KEYINPUT115), .B(new_n767), .C1(new_n617), .C2(new_n623), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n575), .A2(new_n472), .B1(new_n582), .B2(new_n590), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n673), .B(new_n676), .C1(new_n599), .C2(new_n590), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n773), .A2(new_n774), .A3(new_n684), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n705), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n765), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n715), .A2(new_n648), .A3(new_n635), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n686), .A2(new_n778), .A3(new_n339), .A4(new_n651), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n637), .A2(new_n663), .A3(new_n711), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n617), .A2(new_n571), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n783), .B(new_n340), .C1(new_n636), .C2(new_n662), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(KEYINPUT52), .A3(new_n711), .A4(new_n779), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n781), .A2(KEYINPUT116), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n790));
  NAND4_X1  g604(.A1(new_n784), .A2(new_n711), .A3(new_n779), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT53), .B1(new_n777), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n787), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g609(.A(KEYINPUT117), .B(KEYINPUT53), .C1(new_n777), .C2(new_n792), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT54), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n782), .A2(new_n785), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n773), .A2(new_n774), .A3(new_n684), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n694), .A2(new_n701), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n703), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n694), .A2(KEYINPUT108), .A3(new_n701), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n800), .B1(new_n804), .B2(new_n689), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n720), .A2(new_n723), .B1(new_n636), .B2(new_n717), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n772), .A3(new_n764), .A4(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n798), .B1(new_n799), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT118), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n808), .A2(new_n813), .A3(new_n810), .A4(new_n809), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n797), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n714), .A2(new_n672), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT120), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n648), .A2(new_n466), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n817), .A2(new_n713), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n622), .A3(new_n589), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n736), .A2(new_n466), .A3(new_n817), .ZN(new_n822));
  INV_X1    g636(.A(new_n710), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n804), .A2(new_n466), .A3(new_n736), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n642), .A2(new_n674), .A3(new_n672), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n736), .A2(new_n466), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT50), .A3(new_n804), .A4(new_n827), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n824), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n826), .B2(new_n746), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n830), .A2(KEYINPUT119), .A3(new_n804), .A4(new_n745), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n669), .A2(new_n671), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n756), .B1(new_n188), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n832), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT51), .B1(new_n832), .B2(new_n838), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT48), .ZN(new_n841));
  INV_X1    g655(.A(new_n721), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n822), .A2(KEYINPUT121), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n830), .A2(new_n682), .A3(new_n804), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT121), .B(KEYINPUT48), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n822), .B2(new_n842), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n462), .B1(new_n820), .B2(new_n590), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OR4_X1    g662(.A1(new_n839), .A2(new_n840), .A3(new_n843), .A4(new_n848), .ZN(new_n849));
  OAI22_X1  g663(.A1(new_n815), .A2(new_n849), .B1(G952), .B2(G953), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n657), .A2(new_n674), .A3(new_n188), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n836), .B2(KEYINPUT49), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n643), .A2(new_n852), .A3(new_n648), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n622), .A3(new_n694), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n850), .A2(new_n855), .ZN(G75));
  NOR2_X1   g670(.A1(new_n253), .A2(G952), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n808), .A2(new_n810), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(G210), .A3(G902), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n309), .A2(new_n311), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n332), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n312), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n858), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT56), .B1(new_n860), .B2(KEYINPUT122), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(KEYINPUT122), .B2(new_n860), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n869), .B2(new_n865), .ZN(G51));
  XNOR2_X1  g684(.A(new_n192), .B(KEYINPUT57), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n809), .B1(new_n808), .B2(new_n810), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(KEYINPUT123), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n665), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n859), .A2(G902), .A3(new_n740), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n857), .B1(new_n878), .B2(new_n879), .ZN(G54));
  INV_X1    g694(.A(new_n407), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n859), .A2(G902), .ZN(new_n882));
  NAND2_X1  g696(.A1(KEYINPUT58), .A2(G475), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n858), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n882), .A2(new_n881), .A3(new_n883), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(G60));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n888));
  NAND2_X1  g702(.A1(G478), .A2(G902), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT59), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n586), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n777), .B2(new_n786), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n894), .B2(new_n811), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n888), .B1(new_n895), .B2(new_n857), .ZN(new_n896));
  INV_X1    g710(.A(new_n891), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n872), .B2(new_n873), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(KEYINPUT124), .A3(new_n858), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n586), .B1(new_n815), .B2(new_n890), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(G63));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n903));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n892), .A2(new_n893), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n905), .B(new_n906), .C1(new_n608), .C2(new_n607), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n905), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n502), .A2(new_n572), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n858), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n903), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  INV_X1    g726(.A(new_n608), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n908), .B1(new_n913), .B2(new_n606), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n914), .A3(KEYINPUT61), .A4(new_n858), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(new_n915), .ZN(G66));
  INV_X1    g730(.A(G224), .ZN(new_n917));
  OAI21_X1  g731(.A(G953), .B1(new_n467), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n776), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n862), .B1(G898), .B2(new_n253), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT125), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n920), .B(new_n922), .ZN(G69));
  AOI21_X1  g737(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n751), .A2(new_n758), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n784), .A2(new_n711), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n744), .A2(new_n747), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n339), .A3(new_n686), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n726), .B1(new_n929), .B2(new_n842), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n720), .B2(new_n723), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n925), .A2(new_n253), .A3(new_n927), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n528), .A2(new_n533), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n373), .A2(new_n374), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(G900), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n253), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n924), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n717), .A2(new_n652), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n590), .B1(new_n622), .B2(new_n458), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n927), .A2(new_n655), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n927), .A2(KEYINPUT62), .A3(new_n655), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(G953), .B1(new_n947), .B2(new_n925), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n939), .B(KEYINPUT126), .C1(new_n935), .C2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n935), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n751), .A2(new_n931), .A3(new_n758), .A4(new_n927), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n938), .B1(new_n952), .B2(G953), .ZN(new_n953));
  INV_X1    g767(.A(new_n924), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n950), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n949), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n932), .A2(new_n958), .A3(new_n938), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n959), .B(new_n960), .C1(new_n935), .C2(new_n948), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n924), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n957), .A2(new_n962), .ZN(G72));
  AND3_X1   g777(.A1(new_n947), .A2(new_n925), .A3(new_n919), .ZN(new_n964));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n646), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n952), .B2(new_n776), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n857), .B1(new_n969), .B2(new_n557), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n795), .A2(new_n796), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n557), .A2(new_n646), .A3(new_n967), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G57));
endmodule


