//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT64), .B(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT2), .B(G226), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G68), .B(G77), .ZN(new_n234));
  INV_X1    g0034(.A(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT65), .B(G50), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G351));
  AND2_X1   g0043(.A1(G1), .A2(G13), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  INV_X1    g0047(.A(G45), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n246), .A2(G274), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G226), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n255), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1698), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n259), .B1(G222), .B2(new_n264), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n250), .B1(new_n251), .B2(new_n254), .C1(new_n265), .C2(new_n246), .ZN(new_n266));
  INV_X1    g0066(.A(G169), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT69), .B(KEYINPUT8), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n210), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n211), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  INV_X1    g0083(.A(G20), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n283), .A2(new_n284), .A3(G1), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n277), .A2(new_n282), .B1(new_n202), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n281), .B1(G1), .B2(new_n284), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n202), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n268), .B(new_n288), .C1(G179), .C2(new_n266), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n266), .A2(G200), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT72), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n291), .A2(KEYINPUT10), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT71), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n288), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n288), .B(KEYINPUT71), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n290), .B1(new_n301), .B2(new_n266), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n293), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  AOI211_X1 g0104(.A(new_n292), .B(new_n302), .C1(new_n296), .C2(new_n299), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n289), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n271), .A2(new_n285), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n271), .B2(new_n287), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n250), .B1(new_n254), .B2(new_n226), .ZN(new_n310));
  INV_X1    g0110(.A(G1698), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n257), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n251), .A2(G1698), .ZN(new_n313));
  AND2_X1   g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n246), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n301), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G200), .B2(new_n319), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT75), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n314), .A2(new_n315), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n210), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n262), .A2(new_n284), .A3(new_n263), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n327), .A3(G68), .ZN(new_n328));
  AND2_X1   g0128(.A1(G58), .A2(G68), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n329), .B2(new_n201), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n275), .A2(G159), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AND4_X1   g0133(.A1(new_n322), .A2(new_n328), .A3(KEYINPUT16), .A4(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G68), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n326), .B2(KEYINPUT7), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n336), .B2(new_n325), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n322), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n284), .A2(KEYINPUT64), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT64), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G20), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT7), .B1(new_n343), .B2(new_n255), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n323), .A2(new_n324), .A3(new_n284), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(G68), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n333), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n279), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n309), .B(new_n321), .C1(new_n339), .C2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT17), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n314), .A2(new_n315), .A3(G20), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n354), .B2(new_n324), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n323), .A2(new_n210), .A3(new_n324), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT16), .B(new_n333), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT75), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n337), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n279), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n347), .B2(new_n348), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n308), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT17), .A3(new_n321), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n353), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n318), .ZN(new_n366));
  INV_X1    g0166(.A(G179), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n247), .A2(new_n248), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n252), .A2(new_n368), .B1(new_n244), .B2(new_n245), .ZN(new_n369));
  INV_X1    g0169(.A(G274), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n244), .B2(new_n245), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n369), .A2(G232), .B1(new_n371), .B2(new_n249), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n366), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n267), .B1(new_n310), .B2(new_n318), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n366), .A2(new_n372), .A3(new_n376), .A4(new_n367), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n360), .A2(new_n362), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n309), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT77), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT18), .B1(new_n363), .B2(new_n378), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n383), .B1(new_n382), .B2(new_n384), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n365), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n273), .A2(G77), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n275), .A2(G50), .B1(G20), .B2(new_n335), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n281), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(KEYINPUT11), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(KEYINPUT11), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n283), .A2(G1), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G20), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n394), .A2(KEYINPUT12), .A3(G68), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT12), .B1(new_n394), .B2(G68), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n285), .A2(new_n279), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n335), .B1(new_n252), .B2(G20), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n395), .A2(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n391), .A2(new_n392), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n251), .A2(new_n311), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n226), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n314), .C2(new_n315), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n246), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT73), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n246), .A2(G238), .A3(new_n253), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT74), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n250), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n250), .B2(new_n409), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n404), .A2(new_n405), .ZN(new_n416));
  INV_X1    g0216(.A(new_n245), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n211), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n407), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI211_X1 g0219(.A(KEYINPUT73), .B(new_n246), .C1(new_n404), .C2(new_n405), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n419), .A2(new_n420), .B1(new_n411), .B2(new_n412), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT13), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n415), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(G169), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(new_n422), .A3(G179), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n423), .B2(G169), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n401), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n415), .A2(new_n422), .A3(G190), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n415), .A2(new_n422), .ZN(new_n431));
  INV_X1    g0231(.A(G200), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n400), .B(new_n430), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT8), .B(G58), .ZN(new_n434));
  INV_X1    g0234(.A(new_n275), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n258), .A2(new_n210), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n273), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n361), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n361), .A2(new_n394), .ZN(new_n441));
  OAI21_X1  g0241(.A(G77), .B1(new_n284), .B2(G1), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n441), .A2(new_n442), .B1(G77), .B2(new_n394), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G244), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n250), .B1(new_n254), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n264), .A2(G232), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  INV_X1    g0249(.A(G238), .ZN(new_n450));
  OAI221_X1 g0250(.A(new_n448), .B1(new_n449), .B2(new_n255), .C1(new_n450), .C2(new_n256), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(KEYINPUT70), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n246), .B1(new_n451), .B2(KEYINPUT70), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n445), .B1(new_n454), .B2(G190), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n432), .B2(new_n454), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n454), .A2(G169), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n444), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n367), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n429), .A2(new_n433), .A3(new_n456), .A4(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n306), .A2(new_n387), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT87), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT85), .ZN(new_n464));
  OAI211_X1 g0264(.A(G257), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT83), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT83), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n255), .A2(new_n467), .A3(G257), .A4(G1698), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT84), .B(G294), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G33), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n255), .A2(G250), .A3(new_n311), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n418), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n248), .A2(G1), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n477), .A2(G264), .A3(new_n246), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n464), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  AOI211_X1 g0280(.A(KEYINPUT85), .B(new_n478), .C1(new_n472), .C2(new_n418), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n371), .A2(new_n474), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT86), .B1(new_n485), .B2(G200), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n473), .A2(new_n479), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT85), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n478), .B1(new_n472), .B2(new_n418), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n464), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n483), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT86), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(new_n432), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n483), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G190), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n486), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n210), .A2(new_n255), .A3(G87), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT22), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT24), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT23), .A2(G107), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(G20), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT23), .A2(G107), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n343), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n499), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n500), .B1(new_n499), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n279), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n285), .A2(new_n449), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n509), .B(KEYINPUT25), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n261), .A2(G1), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n285), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n281), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n513), .B2(G107), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n497), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n488), .A2(G179), .A3(new_n483), .A4(new_n490), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n494), .A2(G169), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n515), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n463), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n518), .A2(new_n519), .B1(new_n508), .B2(new_n514), .ZN(new_n523));
  AOI211_X1 g0323(.A(KEYINPUT87), .B(new_n523), .C1(new_n497), .C2(new_n516), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n340), .A2(new_n342), .A3(G33), .A4(G97), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR3_X1    g0328(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n405), .A2(new_n527), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n343), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n210), .A2(new_n255), .A3(G68), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n279), .B1(new_n285), .B2(new_n437), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n281), .A2(G87), .A3(new_n512), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n255), .A2(G238), .A3(new_n311), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  OAI211_X1 g0338(.A(G244), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n418), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n246), .A2(G274), .A3(new_n474), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n252), .A2(G45), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n543), .B(G250), .C1(new_n417), .C2(new_n211), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n540), .B2(new_n418), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G190), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n536), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n513), .A2(new_n438), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(new_n534), .B1(new_n367), .B2(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(new_n267), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n418), .B1(new_n474), .B2(new_n482), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n484), .B1(G257), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(new_n311), .C1(new_n314), .C2(new_n315), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  OAI211_X1 g0363(.A(G250), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n559), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT78), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(new_n418), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n566), .B1(new_n565), .B2(new_n418), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n367), .B(new_n558), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n563), .B(new_n564), .C1(new_n560), .C2(new_n561), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT4), .B1(new_n264), .B2(G244), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n418), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n558), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n267), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n281), .A2(G97), .A3(new_n512), .ZN(new_n576));
  INV_X1    g0376(.A(G97), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n285), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n344), .A2(G107), .A3(new_n345), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n583), .A2(new_n577), .A3(G107), .ZN(new_n584));
  XNOR2_X1  g0384(.A(G97), .B(G107), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n586), .A2(new_n210), .B1(new_n258), .B2(new_n435), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n279), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n580), .A2(new_n588), .A3(KEYINPUT79), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT79), .B1(new_n580), .B2(new_n588), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n570), .B(new_n575), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n583), .ZN(new_n592));
  INV_X1    g0392(.A(new_n584), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n343), .B1(G77), .B2(new_n275), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n361), .B1(new_n595), .B2(new_n581), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n579), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n558), .A2(new_n573), .A3(G190), .ZN(new_n598));
  INV_X1    g0398(.A(new_n558), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n573), .A2(KEYINPUT78), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n567), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n597), .B(new_n598), .C1(new_n601), .C2(new_n432), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n556), .A2(new_n591), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(G116), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n511), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n441), .A2(new_n606), .B1(G116), .B2(new_n394), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(G20), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n563), .B1(new_n577), .B2(G33), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n279), .B(new_n608), .C1(new_n343), .C2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT20), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n607), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n477), .A2(G270), .A3(new_n246), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n483), .ZN(new_n616));
  OAI211_X1 g0416(.A(G257), .B(new_n311), .C1(new_n314), .C2(new_n315), .ZN(new_n617));
  OAI211_X1 g0417(.A(G264), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n618));
  INV_X1    g0418(.A(G303), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n255), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n616), .B1(new_n418), .B2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n614), .B(KEYINPUT81), .C1(new_n621), .C2(new_n432), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT81), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n615), .A2(new_n483), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n620), .A2(new_n418), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n432), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n397), .A2(new_n605), .B1(new_n604), .B2(new_n285), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n610), .A2(new_n611), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n610), .A2(new_n611), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n623), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n625), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n622), .B(new_n631), .C1(new_n301), .C2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n267), .B1(new_n624), .B2(new_n625), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n630), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT80), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n632), .A2(KEYINPUT21), .A3(G169), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n624), .A2(new_n625), .A3(G179), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n641), .B2(new_n630), .ZN(new_n642));
  AOI211_X1 g0442(.A(KEYINPUT80), .B(new_n614), .C1(new_n639), .C2(new_n640), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n633), .B(new_n637), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT82), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n634), .A2(KEYINPUT21), .B1(new_n621), .B2(G179), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT80), .B1(new_n646), .B2(new_n614), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n641), .A2(new_n638), .A3(new_n630), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT82), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(new_n633), .A4(new_n637), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n603), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n462), .A2(new_n525), .A3(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n289), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n304), .A2(new_n305), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n433), .A2(new_n458), .A3(new_n459), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n429), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n365), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n382), .A2(new_n384), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n654), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n462), .ZN(new_n663));
  INV_X1    g0463(.A(new_n597), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n664), .A2(new_n570), .A3(new_n575), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n542), .A2(new_n667), .A3(new_n544), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n542), .B2(new_n544), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n541), .ZN(new_n672));
  OAI21_X1  g0472(.A(G200), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n536), .A2(new_n666), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n534), .A2(new_n535), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n545), .A2(KEYINPUT88), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n668), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n432), .B1(new_n677), .B2(new_n541), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT89), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n674), .A2(new_n679), .A3(new_n550), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n676), .A2(new_n668), .B1(new_n418), .B2(new_n540), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n553), .B1(G169), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n665), .A2(new_n680), .A3(new_n681), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n551), .A2(new_n555), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT26), .B1(new_n591), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n684), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n591), .A2(new_n680), .A3(new_n602), .A4(new_n683), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n517), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n641), .A2(new_n630), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n637), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n521), .A2(KEYINPUT90), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT90), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n523), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n692), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n687), .B1(new_n690), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n662), .B1(new_n663), .B2(new_n698), .ZN(G369));
  NAND2_X1  g0499(.A1(new_n210), .A2(new_n393), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT91), .Z(new_n701));
  INV_X1    g0501(.A(KEYINPUT27), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(G213), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n525), .B1(new_n516), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n523), .A2(new_n707), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n645), .A2(new_n651), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n614), .B2(new_n708), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n692), .A2(new_n630), .A3(new_n707), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n693), .A2(new_n695), .A3(new_n708), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n647), .A2(new_n648), .B1(new_n636), .B2(new_n635), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n707), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n525), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n207), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n529), .A2(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n215), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n491), .A2(new_n432), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n495), .B1(new_n730), .B2(KEYINPUT86), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n515), .B1(new_n731), .B2(new_n493), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT87), .B1(new_n732), .B2(new_n523), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n517), .A2(new_n463), .A3(new_n521), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n652), .A4(new_n708), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n480), .A2(new_n481), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n574), .A2(new_n640), .A3(new_n547), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT30), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n558), .B1(new_n568), .B2(new_n569), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n682), .A2(new_n621), .A3(G179), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n491), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n707), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT31), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n735), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(KEYINPUT92), .B1(new_n748), .B2(G330), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT92), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n750), .B(new_n712), .C1(new_n735), .C2(new_n747), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n534), .B(new_n535), .C1(new_n682), .C2(new_n432), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n550), .B1(new_n753), .B2(KEYINPUT89), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n666), .B1(new_n536), .B2(new_n673), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n683), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n601), .A2(new_n367), .B1(new_n267), .B2(new_n574), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n664), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT26), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n589), .A2(new_n590), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n556), .A2(new_n760), .A3(new_n681), .A4(new_n757), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(new_n683), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT94), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n637), .B1(new_n642), .B2(new_n643), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n523), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n719), .A2(new_n521), .A3(KEYINPUT94), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n688), .B1(new_n516), .B2(new_n497), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n707), .ZN(new_n770));
  INV_X1    g0570(.A(new_n692), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n520), .A2(new_n694), .A3(new_n515), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n694), .B1(new_n520), .B2(new_n515), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n707), .B1(new_n775), .B2(new_n687), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n778));
  AOI22_X1  g0578(.A1(new_n770), .A2(KEYINPUT29), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n752), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n729), .B1(new_n780), .B2(G1), .ZN(G364));
  NOR2_X1   g0581(.A1(new_n343), .A2(new_n283), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G45), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n784), .A2(new_n252), .A3(new_n724), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n716), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n714), .A2(new_n715), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(G330), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n284), .B1(KEYINPUT96), .B2(new_n267), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n267), .A2(KEYINPUT96), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n211), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n432), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(G20), .A3(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G87), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n255), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G179), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n343), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n796), .B1(G97), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n801));
  NOR2_X1   g0601(.A1(new_n210), .A2(G190), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n797), .ZN(new_n803));
  INV_X1    g0603(.A(G159), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n367), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n800), .B(new_n805), .C1(new_n258), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n367), .A2(new_n432), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n343), .A2(G190), .A3(new_n809), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n811), .A2(G68), .B1(G50), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n802), .A2(new_n792), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G107), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n343), .A2(G190), .A3(new_n806), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n814), .B(new_n817), .C1(new_n235), .C2(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n803), .A2(new_n804), .A3(new_n801), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n808), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n803), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G283), .A2(new_n816), .B1(new_n822), .B2(G329), .ZN(new_n823));
  XOR2_X1   g0623(.A(KEYINPUT33), .B(G317), .Z(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n810), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n818), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G322), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n255), .B1(new_n794), .B2(G303), .ZN(new_n828));
  INV_X1    g0628(.A(new_n469), .ZN(new_n829));
  INV_X1    g0629(.A(new_n799), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  INV_X1    g0632(.A(G326), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n807), .A2(new_n832), .B1(new_n833), .B2(new_n812), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n825), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n791), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n785), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n255), .A2(new_n207), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(KEYINPUT95), .B2(G355), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(KEYINPUT95), .B2(G355), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n238), .A2(G45), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n723), .A2(new_n255), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(G45), .B2(new_n215), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n840), .B1(G116), .B2(new_n207), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(G13), .A2(G33), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(G20), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n791), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n837), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n847), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n836), .B(new_n849), .C1(new_n787), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n788), .A2(new_n851), .ZN(G396));
  NOR2_X1   g0652(.A1(new_n791), .A2(new_n845), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n785), .B1(new_n854), .B2(G77), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n458), .A2(new_n459), .A3(new_n708), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n456), .B1(new_n444), .B2(new_n708), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n460), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(new_n846), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n816), .A2(G87), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n860), .B1(new_n619), .B2(new_n812), .C1(new_n832), .C2(new_n803), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n255), .B1(new_n794), .B2(G107), .ZN(new_n862));
  INV_X1    g0662(.A(G283), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n862), .B1(new_n830), .B2(new_n577), .C1(new_n863), .C2(new_n810), .ZN(new_n864));
  INV_X1    g0664(.A(G294), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n807), .A2(new_n604), .B1(new_n865), .B2(new_n818), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n861), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT98), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n822), .A2(G132), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n816), .A2(G68), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n799), .A2(G58), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n323), .B1(new_n794), .B2(G50), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n870), .A2(new_n871), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G137), .A2(new_n813), .B1(new_n826), .B2(G143), .ZN(new_n875));
  INV_X1    g0675(.A(G150), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n875), .B1(new_n876), .B2(new_n810), .C1(new_n804), .C2(new_n807), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT34), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n869), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n881), .A2(KEYINPUT99), .ZN(new_n882));
  INV_X1    g0682(.A(new_n791), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n881), .B2(KEYINPUT99), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n855), .B(new_n859), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n752), .ZN(new_n886));
  INV_X1    g0686(.A(new_n858), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n777), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n697), .A2(new_n708), .A3(new_n858), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n785), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n752), .A2(new_n888), .A3(new_n889), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n885), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(G384));
  NAND2_X1  g0694(.A1(new_n779), .A2(new_n462), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n662), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT108), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n377), .A2(new_n375), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n376), .B1(new_n319), .B2(new_n367), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n282), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n358), .B2(new_n359), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n902), .B2(new_n308), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT102), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n351), .A3(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n703), .A2(new_n704), .A3(G213), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n902), .B2(new_n308), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n904), .B1(new_n903), .B2(new_n351), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT103), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT103), .B(KEYINPUT37), .C1(new_n908), .C2(new_n909), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n379), .A2(new_n309), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT104), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n906), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT104), .B1(new_n363), .B2(new_n705), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n380), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n351), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n912), .A2(new_n913), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n907), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n387), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n921), .A2(KEYINPUT38), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n401), .A2(new_n707), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n429), .A2(new_n433), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT14), .B1(new_n431), .B2(new_n267), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n433), .A2(new_n931), .A3(new_n426), .A4(new_n425), .ZN(new_n932));
  INV_X1    g0732(.A(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n930), .A2(KEYINPUT101), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT101), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n429), .A2(new_n936), .A3(new_n433), .A4(new_n929), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n856), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n889), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n928), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n659), .A2(new_n705), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n918), .A2(new_n351), .ZN(new_n944));
  AOI211_X1 g0744(.A(KEYINPUT106), .B(new_n380), .C1(new_n916), .C2(new_n917), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n944), .B1(new_n945), .B2(new_n919), .ZN(new_n946));
  INV_X1    g0746(.A(new_n919), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n918), .A2(KEYINPUT106), .A3(new_n351), .A4(new_n947), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n382), .A2(new_n353), .A3(new_n364), .A4(new_n384), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n916), .A3(new_n917), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n925), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n927), .A2(new_n952), .A3(KEYINPUT107), .A4(new_n953), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n921), .A2(KEYINPUT38), .A3(new_n923), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT107), .B1(new_n951), .B2(new_n925), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n921), .B2(new_n923), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n954), .B1(new_n958), .B2(new_n953), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n429), .A2(new_n707), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n943), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n897), .B(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT109), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n927), .A2(new_n952), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n935), .A2(new_n858), .A3(new_n937), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n748), .A2(new_n966), .A3(KEYINPUT40), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n964), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n935), .A2(new_n858), .A3(new_n937), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n735), .B2(new_n747), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n927), .A2(new_n952), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT109), .A4(KEYINPUT40), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT40), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n970), .B1(new_n955), .B2(new_n957), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n968), .A2(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n462), .A2(new_n748), .ZN(new_n977));
  OAI21_X1  g0777(.A(G330), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n977), .B2(new_n976), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n963), .A2(new_n979), .B1(new_n252), .B2(new_n782), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n963), .B2(new_n979), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n982), .A2(G116), .A3(new_n212), .A4(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  OR3_X1    g0786(.A1(new_n215), .A2(new_n258), .A3(new_n329), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n202), .A2(G68), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n252), .B(G13), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  OR3_X1    g0789(.A1(new_n981), .A2(new_n986), .A3(new_n989), .ZN(G367));
  NAND2_X1  g0790(.A1(new_n707), .A2(new_n675), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(new_n683), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n683), .A3(new_n680), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(KEYINPUT43), .B2(new_n994), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n708), .A2(new_n597), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n591), .B2(new_n602), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n757), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n1000), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n721), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT42), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n591), .B1(new_n1004), .B2(new_n521), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n708), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  MUX2_X1   g0809(.A(new_n998), .B(new_n999), .S(new_n1009), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n717), .B2(new_n1004), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n1010), .A2(new_n717), .A3(new_n1004), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n724), .B(KEYINPUT41), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n721), .A2(new_n718), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n1004), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1004), .ZN(new_n1017));
  XOR2_X1   g0817(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n717), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n721), .B1(new_n711), .B2(new_n720), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(new_n716), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(new_n780), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1013), .B1(new_n1025), .B2(new_n780), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n784), .A2(new_n252), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1011), .B(new_n1012), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n842), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n232), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n848), .B1(new_n207), .B2(new_n437), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n785), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n794), .A2(G116), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT46), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n816), .A2(G97), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n807), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(G283), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n811), .A2(new_n469), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n323), .B1(new_n812), .B2(new_n832), .C1(new_n830), .C2(new_n449), .ZN(new_n1041));
  INV_X1    g0841(.A(G317), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n803), .A2(new_n1042), .B1(new_n619), .B2(new_n818), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT112), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n793), .A2(new_n235), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n830), .A2(new_n335), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(G159), .C2(new_n811), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1037), .A2(G50), .B1(G150), .B2(new_n826), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n822), .A2(G137), .B1(G143), .B2(new_n813), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n816), .A2(G77), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n255), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT113), .Z(new_n1054));
  OAI21_X1  g0854(.A(new_n1045), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT47), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1033), .B1(new_n1056), .B2(new_n791), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n850), .B2(new_n994), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1029), .A2(new_n1058), .ZN(G387));
  NAND3_X1  g0859(.A1(new_n709), .A2(new_n710), .A3(new_n847), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n726), .A2(new_n838), .B1(G107), .B2(new_n207), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n229), .A2(new_n248), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n726), .ZN(new_n1063));
  AOI211_X1 g0863(.A(G45), .B(new_n1063), .C1(G68), .C2(G77), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n434), .A2(G50), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT50), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1030), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1061), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n848), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n785), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n803), .A2(new_n876), .B1(new_n258), .B2(new_n793), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT114), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n799), .A2(new_n438), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1036), .A2(new_n255), .A3(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n811), .A2(new_n271), .B1(G159), .B2(new_n813), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1037), .A2(G68), .B1(G50), .B2(new_n826), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n830), .A2(new_n863), .B1(new_n829), .B2(new_n793), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G317), .A2(new_n826), .B1(new_n813), .B2(G322), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n619), .B2(new_n807), .C1(new_n832), .C2(new_n810), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT48), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1081), .B2(new_n1080), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT115), .Z(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT49), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n255), .B1(new_n822), .B2(G326), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n604), .C2(new_n815), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1084), .A2(KEYINPUT49), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1077), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1070), .B1(new_n1089), .B2(new_n791), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1023), .A2(new_n1028), .B1(new_n1060), .B2(new_n1090), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1024), .A2(new_n725), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1023), .A2(new_n780), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(G393));
  AOI21_X1  g0894(.A(new_n725), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1024), .B2(new_n1021), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n202), .A2(new_n810), .B1(new_n807), .B2(new_n434), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n799), .A2(G77), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n323), .B1(new_n794), .B2(G68), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n860), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1097), .B(new_n1100), .C1(G143), .C2(new_n822), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n876), .A2(new_n812), .B1(new_n818), .B2(new_n804), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n832), .A2(new_n818), .B1(new_n812), .B2(new_n1042), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G303), .A2(new_n811), .B1(new_n822), .B2(G322), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n865), .B2(new_n807), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n255), .B1(new_n794), .B2(G283), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n817), .B(new_n1108), .C1(new_n604), .C2(new_n830), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1101), .A2(new_n1103), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1111), .A2(new_n883), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n242), .A2(new_n842), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1069), .B1(G97), .B2(new_n723), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n837), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT116), .Z(new_n1116));
  AOI211_X1 g0916(.A(new_n1112), .B(new_n1116), .C1(new_n1004), .C2(new_n847), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n1021), .B2(new_n1028), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1096), .A2(new_n1118), .ZN(G390));
  INV_X1    g0919(.A(new_n938), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n752), .A2(KEYINPUT119), .A3(new_n858), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT31), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n746), .B(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n603), .B(new_n707), .C1(new_n645), .C2(new_n651), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n525), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n750), .B1(new_n1125), .B2(new_n712), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n748), .A2(KEYINPUT92), .A3(G330), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n858), .A4(new_n1120), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT119), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1121), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT117), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n857), .A2(new_n460), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n769), .A2(new_n707), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1132), .B1(new_n1135), .B2(new_n856), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n767), .A2(new_n768), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n708), .B(new_n1133), .C1(new_n1137), .C2(new_n762), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(KEYINPUT117), .A3(new_n939), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(new_n1120), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n965), .A2(new_n961), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT39), .B1(new_n928), .B2(new_n956), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT118), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n940), .B2(new_n961), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n856), .B1(new_n776), .B2(new_n858), .ZN(new_n1146));
  OAI211_X1 g0946(.A(KEYINPUT118), .B(new_n960), .C1(new_n1146), .C2(new_n938), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1143), .A2(new_n954), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1131), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1142), .B1(new_n959), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n748), .A2(new_n966), .A3(G330), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1028), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n271), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n837), .B1(new_n1157), .B2(new_n853), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n811), .A2(G107), .B1(G283), .B2(new_n813), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n865), .B2(new_n803), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n871), .A2(new_n323), .A3(new_n795), .A4(new_n1098), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n807), .A2(new_n577), .B1(new_n604), .B2(new_n818), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n794), .A2(G150), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT122), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT53), .Z(new_n1166));
  INV_X1    g0966(.A(G132), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n255), .B1(new_n818), .B2(new_n1167), .C1(new_n830), .C2(new_n804), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n202), .A2(new_n815), .B1(new_n807), .B2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1166), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(G125), .ZN(new_n1172));
  INV_X1    g0972(.A(G128), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n803), .A2(new_n1172), .B1(new_n1173), .B2(new_n812), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G137), .B2(new_n811), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1163), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1158), .B1(new_n883), .B2(new_n1176), .C1(new_n959), .C2(new_n846), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1156), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1146), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1126), .A2(new_n1127), .A3(new_n858), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(KEYINPUT120), .A3(new_n938), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1152), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT120), .B1(new_n1181), .B2(new_n938), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n748), .A2(G330), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n938), .B1(new_n1187), .B2(new_n887), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1131), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n663), .A2(new_n1187), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n896), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1194));
  OAI211_X1 g0994(.A(KEYINPUT121), .B(new_n724), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1192), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n725), .B1(new_n1199), .B2(new_n1155), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(KEYINPUT121), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1179), .B1(new_n1197), .B2(new_n1201), .ZN(G378));
  OAI22_X1  g1002(.A1(new_n830), .A2(new_n876), .B1(new_n793), .B2(new_n1169), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1037), .A2(G137), .B1(G128), .B2(new_n826), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1172), .B2(new_n812), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G132), .C2(new_n811), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n261), .B(new_n247), .C1(new_n815), .C2(new_n804), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G124), .B2(new_n822), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n807), .A2(new_n437), .B1(new_n449), .B2(new_n818), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n323), .A2(new_n247), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1214), .B(new_n1047), .C1(G77), .C2(new_n794), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G58), .A2(new_n816), .B1(new_n822), .B2(G283), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n577), .C2(new_n810), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1213), .B(new_n1217), .C1(G116), .C2(new_n813), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT58), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(KEYINPUT58), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1214), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1221));
  AND4_X1   g1021(.A1(new_n1212), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n785), .B1(G50), .B2(new_n854), .C1(new_n1222), .C2(new_n883), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n297), .A2(new_n705), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n306), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n306), .A2(new_n1226), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1225), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1226), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n655), .A2(new_n289), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n306), .A2(new_n1226), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1224), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1223), .B1(new_n1235), .B2(new_n845), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n962), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n968), .A2(new_n972), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n974), .A2(new_n973), .ZN(new_n1239));
  AND4_X1   g1039(.A1(G330), .A2(new_n1234), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1234), .B1(new_n975), .B2(G330), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1237), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1238), .A2(G330), .A3(new_n1239), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1235), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n975), .A2(G330), .A3(new_n1234), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n962), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1236), .B1(new_n1247), .B2(new_n1028), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1244), .A2(new_n962), .A3(new_n1245), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n962), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1198), .B1(new_n1155), .B2(new_n1190), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n724), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1121), .B2(new_n1130), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT120), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n749), .A2(new_n751), .A3(new_n887), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(new_n1120), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n1152), .A3(new_n1182), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1255), .B1(new_n1259), .B2(new_n1180), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1192), .B1(new_n1260), .B2(new_n1194), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT57), .B1(new_n1261), .B2(new_n1247), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1248), .B1(new_n1253), .B2(new_n1262), .ZN(G375));
  NAND3_X1  g1063(.A1(new_n1185), .A2(new_n1189), .A3(new_n1198), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT123), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1260), .A2(KEYINPUT123), .A3(new_n1198), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1013), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1193), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n837), .B1(new_n335), .B2(new_n853), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n255), .B1(new_n804), .B2(new_n793), .C1(new_n830), .C2(new_n202), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G128), .A2(new_n822), .B1(new_n1037), .B2(G150), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n826), .A2(G137), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1272), .B(new_n1273), .C1(new_n810), .C2(new_n1169), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1271), .B(new_n1274), .C1(G58), .C2(new_n816), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n813), .A2(G132), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT124), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n604), .A2(new_n810), .B1(new_n803), .B2(new_n619), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G294), .B2(new_n813), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1037), .A2(G107), .B1(G283), .B2(new_n826), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n255), .B1(new_n794), .B2(G97), .ZN(new_n1281));
  AND4_X1   g1081(.A1(new_n1052), .A2(new_n1280), .A3(new_n1073), .A4(new_n1281), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1275), .A2(new_n1277), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n1270), .B1(new_n883), .B2(new_n1283), .C1(new_n1120), .C2(new_n846), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1260), .B2(new_n1027), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1269), .A2(new_n1286), .ZN(G381));
  OR2_X1    g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  OR4_X1    g1088(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1288), .ZN(new_n1289));
  OR4_X1    g1089(.A1(G378), .A2(new_n1289), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1090(.A(G375), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1200), .A2(KEYINPUT121), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1200), .A2(KEYINPUT121), .B1(new_n1194), .B2(new_n1193), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1178), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(G213), .A3(new_n706), .A4(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(G407), .A2(G213), .A3(new_n1295), .ZN(G409));
  NAND3_X1  g1096(.A1(new_n1261), .A2(new_n1268), .A3(new_n1247), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1248), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1298), .B(new_n1179), .C1(new_n1197), .C2(new_n1201), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1294), .B2(G375), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n706), .A2(G213), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n706), .A2(G213), .A3(G2897), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT60), .B1(new_n1260), .B2(new_n1198), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1185), .A2(new_n1189), .A3(KEYINPUT60), .A4(new_n1198), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1307), .A2(new_n724), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G384), .B1(new_n1309), .B2(new_n1286), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n893), .B(new_n1285), .C1(new_n1306), .C2(new_n1308), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1304), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT126), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1303), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1316), .B(new_n1304), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1302), .A2(new_n1313), .A3(new_n1315), .A4(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1300), .A2(new_n1301), .A3(new_n1314), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT62), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1300), .A2(new_n1322), .A3(new_n1301), .A4(new_n1314), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1318), .A2(new_n1319), .A3(new_n1321), .A4(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(G390), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1029), .B2(new_n1058), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(G393), .B(G396), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1328), .B1(new_n1029), .B2(new_n1058), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1325), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G387), .A2(new_n1329), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1333), .B(G390), .C1(new_n1327), .C2(new_n1329), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1324), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  OR2_X1    g1137(.A1(new_n1320), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1338), .A2(new_n1339), .A3(new_n1319), .A4(new_n1318), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1320), .A2(new_n1337), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(KEYINPUT125), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT125), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1320), .A2(new_n1343), .A3(new_n1337), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1336), .B1(new_n1340), .B2(new_n1345), .ZN(G405));
  NOR2_X1   g1146(.A1(new_n1291), .A2(G378), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1294), .A2(G375), .ZN(new_n1348));
  OR3_X1    g1148(.A1(new_n1347), .A2(new_n1348), .A3(new_n1314), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1314), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1335), .B(new_n1351), .ZN(G402));
endmodule


