//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1392, new_n1393;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G20), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n212), .B1(KEYINPUT1), .B2(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G200), .ZN(new_n243));
  INV_X1    g0043(.A(G41), .ZN(new_n244));
  INV_X1    g0044(.A(G45), .ZN(new_n245));
  AOI21_X1  g0045(.A(G1), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  AND4_X1   g0048(.A1(KEYINPUT66), .A2(new_n246), .A3(new_n248), .A4(G274), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n250), .B1(new_n222), .B2(new_n247), .ZN(new_n251));
  AOI21_X1  g0051(.A(KEYINPUT66), .B1(new_n251), .B2(new_n246), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n248), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n246), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n253), .B1(G226), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G222), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n263), .B1(new_n213), .B2(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n254), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n243), .B1(new_n256), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n256), .A2(G190), .A3(new_n267), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n203), .A2(G20), .ZN(new_n273));
  INV_X1    g0073(.A(G150), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n273), .B1(new_n274), .B2(new_n276), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G1), .A2(G13), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT67), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT67), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n281), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(new_n277), .A3(G1), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n280), .A2(new_n287), .B1(new_n202), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n284), .A2(new_n292), .A3(new_n286), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT68), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n293), .A2(new_n294), .B1(new_n296), .B2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n290), .B1(new_n298), .B2(new_n202), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT9), .Z(new_n300));
  NOR2_X1   g0100(.A1(new_n272), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n270), .A4(new_n271), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n302), .B(new_n303), .C1(new_n272), .C2(new_n300), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n256), .A2(new_n308), .A3(new_n267), .ZN(new_n309));
  XOR2_X1   g0109(.A(new_n309), .B(KEYINPUT69), .Z(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n256), .A2(new_n267), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n314), .A2(new_n299), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n310), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n310), .B2(new_n315), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n253), .B1(G244), .B2(new_n255), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n261), .A2(G232), .A3(new_n262), .ZN(new_n320));
  INV_X1    g0120(.A(G238), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n320), .B1(new_n206), .B2(new_n261), .C1(new_n264), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n254), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n243), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT71), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n277), .A2(new_n213), .B1(new_n326), .B2(new_n278), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n279), .A2(new_n276), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n283), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n289), .A2(new_n283), .ZN(new_n330));
  INV_X1    g0130(.A(G77), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n296), .B2(G20), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n330), .A2(new_n332), .B1(new_n213), .B2(new_n289), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  OR3_X1    g0134(.A1(new_n324), .A2(new_n325), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n325), .B1(new_n324), .B2(new_n334), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n319), .A2(new_n323), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n338), .A2(new_n313), .B1(new_n329), .B2(new_n333), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n319), .A2(new_n308), .A3(new_n323), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n307), .A2(new_n318), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G58), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n347), .B2(new_n201), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n275), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(KEYINPUT80), .A2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(KEYINPUT80), .A2(G33), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT3), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n259), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n355), .A2(new_n356), .A3(G20), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n258), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT80), .A2(G33), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n257), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n361), .A2(KEYINPUT81), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT81), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n354), .B2(new_n259), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n277), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n357), .B1(new_n366), .B2(new_n356), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT16), .B(new_n351), .C1(new_n367), .C2(new_n346), .ZN(new_n368));
  INV_X1    g0168(.A(new_n283), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n259), .A2(new_n277), .A3(new_n260), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n359), .A2(new_n257), .A3(new_n360), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n277), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n356), .A2(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n351), .B1(new_n373), .B2(new_n346), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n369), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n279), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n289), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n298), .B2(new_n378), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n265), .A2(new_n262), .ZN(new_n382));
  INV_X1    g0182(.A(G226), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G1698), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n384), .C1(new_n361), .C2(new_n362), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G87), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n248), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n246), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(G232), .A3(new_n248), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n249), .B2(new_n252), .ZN(new_n390));
  OAI21_X1  g0190(.A(G200), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n246), .A2(new_n248), .A3(G274), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT66), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n251), .A2(KEYINPUT66), .A3(new_n246), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n394), .A2(new_n395), .B1(new_n255), .B2(G232), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n382), .A2(new_n384), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n354), .B2(new_n259), .ZN(new_n398));
  INV_X1    g0198(.A(new_n386), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n254), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(new_n400), .A3(G190), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n377), .A2(new_n381), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n380), .B1(new_n368), .B2(new_n376), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n396), .A2(new_n400), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G169), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n396), .A2(G179), .A3(new_n400), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT18), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  INV_X1    g0214(.A(new_n376), .ZN(new_n415));
  INV_X1    g0215(.A(new_n357), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT81), .B1(new_n361), .B2(new_n362), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n354), .A2(new_n364), .A3(new_n259), .ZN(new_n418));
  AOI21_X1  g0218(.A(G20), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(KEYINPUT7), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n350), .B1(new_n420), .B2(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n414), .B(new_n411), .C1(new_n422), .C2(new_n380), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n403), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n406), .A2(new_n413), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT75), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n346), .B1(new_n296), .B2(G20), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n330), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n296), .A2(new_n346), .A3(G13), .A4(G20), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT76), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT12), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n369), .A2(new_n292), .A3(new_n427), .A4(new_n428), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n430), .A2(new_n435), .A3(KEYINPUT77), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT77), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n433), .A2(new_n434), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT12), .B1(new_n431), .B2(new_n432), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n438), .B1(new_n441), .B2(new_n429), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n346), .A2(G20), .ZN(new_n443));
  OAI221_X1 g0243(.A(new_n443), .B1(new_n278), .B2(new_n331), .C1(new_n276), .C2(new_n202), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n287), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT11), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT11), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(new_n287), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n437), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT78), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n437), .A2(new_n442), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n394), .A2(new_n395), .B1(new_n255), .B2(G238), .ZN(new_n455));
  AND2_X1   g0255(.A1(KEYINPUT3), .A2(G33), .ZN(new_n456));
  OAI211_X1 g0256(.A(G232), .B(G1698), .C1(new_n456), .C2(new_n362), .ZN(new_n457));
  OAI211_X1 g0257(.A(G226), .B(new_n262), .C1(new_n456), .C2(new_n362), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G97), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT74), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n460), .A2(new_n461), .A3(new_n254), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n460), .B2(new_n254), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT13), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT13), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n455), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n337), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(G200), .B1(new_n465), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n454), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT79), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n460), .A2(new_n254), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT74), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n460), .A2(new_n461), .A3(new_n254), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n466), .B1(new_n477), .B2(new_n455), .ZN(new_n478));
  INV_X1    g0278(.A(new_n467), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n243), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n468), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(KEYINPUT79), .A3(new_n454), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(G169), .B1(new_n478), .B2(new_n479), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT14), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n465), .A2(G179), .A3(new_n467), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n465), .A2(new_n467), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT14), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(G169), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n454), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n344), .A2(new_n426), .A3(new_n483), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n289), .A2(new_n206), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n495), .B(KEYINPUT25), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n296), .A2(G33), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n284), .A2(new_n292), .A3(new_n286), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n499), .B2(G107), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n352), .A2(new_n353), .ZN(new_n502));
  INV_X1    g0302(.A(G116), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT87), .B1(new_n206), .B2(G20), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT23), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n504), .A2(new_n277), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n277), .B(G87), .C1(new_n361), .C2(new_n362), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(G20), .B1(new_n354), .B2(new_n259), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(KEYINPUT86), .A3(G87), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT22), .ZN(new_n516));
  INV_X1    g0316(.A(new_n261), .ZN(new_n517));
  INV_X1    g0317(.A(G87), .ZN(new_n518));
  OR4_X1    g0318(.A1(KEYINPUT22), .A2(new_n517), .A3(G20), .A4(new_n518), .ZN(new_n519));
  AOI211_X1 g0319(.A(KEYINPUT24), .B(new_n510), .C1(new_n516), .C2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT22), .B1(new_n511), .B2(new_n512), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT86), .B1(new_n514), .B2(G87), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n521), .B1(new_n524), .B2(new_n509), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n283), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT88), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT88), .B(new_n283), .C1(new_n520), .C2(new_n525), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n501), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT5), .B(G41), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n245), .A2(G1), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n248), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(KEYINPUT90), .A3(G264), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT90), .ZN(new_n537));
  INV_X1    g0337(.A(G264), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n359), .A2(new_n360), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n362), .B1(new_n540), .B2(KEYINPUT3), .ZN(new_n541));
  INV_X1    g0341(.A(G250), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n262), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(G257), .B2(new_n262), .ZN(new_n544));
  INV_X1    g0344(.A(G294), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n541), .A2(new_n544), .B1(new_n545), .B2(new_n502), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n536), .A2(new_n539), .B1(new_n254), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n251), .A2(new_n532), .A3(new_n531), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n308), .ZN(new_n550));
  INV_X1    g0350(.A(new_n548), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n536), .B2(new_n539), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(KEYINPUT89), .A3(new_n254), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n546), .A2(new_n254), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n554), .A2(KEYINPUT89), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n550), .B1(new_n556), .B2(G169), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n530), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n549), .A2(new_n243), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n556), .B2(G190), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n530), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G270), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n548), .B1(new_n534), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n538), .A2(G1698), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G257), .B2(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(G303), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n541), .A2(new_n566), .B1(new_n567), .B2(new_n261), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n254), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n308), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G283), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n277), .C1(G33), .C2(new_n205), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n573), .B(new_n283), .C1(new_n277), .C2(G116), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT20), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n330), .A2(G116), .A3(new_n497), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n291), .A2(G20), .A3(new_n503), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n571), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n579), .A2(new_n570), .A3(KEYINPUT21), .A4(G169), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n570), .ZN(new_n583));
  OAI21_X1  g0383(.A(G169), .B1(new_n575), .B2(new_n578), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n579), .B1(G200), .B2(new_n570), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n337), .B2(new_n570), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n535), .A2(G257), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n572), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n355), .A2(G244), .A3(new_n262), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n548), .B(new_n591), .C1(new_n597), .C2(new_n248), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n292), .A2(G97), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n499), .B2(G97), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G97), .A2(G107), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT6), .B1(new_n207), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n605));
  OAI21_X1  g0405(.A(G20), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n275), .A2(G77), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n371), .A2(new_n372), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n370), .A2(new_n356), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n206), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n283), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT82), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n607), .B(new_n606), .C1(new_n373), .C2(new_n206), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n283), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n602), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n599), .B(new_n617), .C1(new_n337), .C2(new_n598), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n612), .A2(KEYINPUT82), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n615), .B1(new_n614), .B2(new_n283), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n601), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n598), .A2(new_n313), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n596), .A2(new_n595), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n254), .B1(new_n623), .B2(new_n594), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(new_n308), .A3(new_n548), .A4(new_n591), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n321), .A2(G1698), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n541), .A2(new_n629), .B1(new_n503), .B2(new_n502), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n214), .B(new_n262), .C1(new_n354), .C2(new_n259), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n254), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n532), .A2(new_n542), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n248), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT83), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT83), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n636), .A3(new_n248), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n635), .A2(new_n637), .B1(new_n251), .B2(new_n532), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n243), .B1(new_n632), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n277), .A2(G33), .A3(G97), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT19), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n644));
  NOR2_X1   g0444(.A1(G97), .A2(G107), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n277), .A2(new_n644), .B1(new_n645), .B2(new_n518), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n641), .A2(new_n640), .A3(new_n642), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI211_X1 g0449(.A(G20), .B(new_n346), .C1(new_n354), .C2(new_n259), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n283), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n326), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n292), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n498), .A2(new_n518), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n651), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT85), .B1(new_n639), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n504), .B1(new_n355), .B2(new_n628), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n355), .A2(G244), .A3(G1698), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n248), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n635), .A2(new_n637), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n251), .A2(new_n532), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(G200), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n648), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n666), .A2(new_n643), .A3(new_n646), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n355), .A2(new_n277), .A3(G68), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n369), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n669), .A2(new_n653), .A3(new_n655), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT85), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n665), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n632), .A2(new_n638), .A3(G190), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n658), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n313), .B1(new_n661), .B2(new_n664), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n632), .A2(new_n638), .A3(new_n308), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n499), .A2(new_n652), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n651), .A2(new_n654), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n590), .A2(new_n627), .A3(new_n680), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n494), .A2(new_n561), .A3(new_n681), .ZN(G372));
  INV_X1    g0482(.A(new_n307), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n413), .A2(new_n423), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n342), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n490), .A2(new_n491), .B1(new_n471), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n406), .A2(new_n424), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n318), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n679), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n665), .A2(new_n670), .A3(new_n673), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n679), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n626), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n613), .A2(new_n616), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n697), .A2(new_n601), .B1(new_n598), .B2(new_n313), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n674), .A2(new_n698), .A3(new_n625), .A4(new_n679), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT26), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n587), .B1(new_n530), .B2(new_n557), .ZN(new_n702));
  INV_X1    g0502(.A(new_n693), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n618), .A3(new_n626), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n530), .B2(new_n560), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n701), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n690), .B1(new_n493), .B2(new_n706), .ZN(G369));
  INV_X1    g0507(.A(new_n291), .ZN(new_n708));
  OR3_X1    g0508(.A1(new_n708), .A2(KEYINPUT27), .A3(G20), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT27), .B1(new_n708), .B2(G20), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G213), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G343), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n558), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n525), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n524), .A2(new_n521), .A3(new_n509), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT88), .B1(new_n717), .B2(new_n283), .ZN(new_n718));
  INV_X1    g0518(.A(new_n529), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n500), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n557), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n500), .B(new_n560), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n713), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n530), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n714), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(KEYINPUT91), .B(G330), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n580), .A3(new_n581), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n579), .A2(new_n713), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n590), .B2(new_n731), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n713), .B(KEYINPUT92), .Z(new_n735));
  NAND2_X1  g0535(.A1(new_n558), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n587), .A2(new_n713), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n723), .B(new_n737), .C1(new_n557), .C2(new_n530), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(G399));
  INV_X1    g0539(.A(new_n210), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G41), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(G1), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n224), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n681), .A2(new_n722), .A3(new_n723), .A4(new_n735), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n661), .A2(new_n664), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n571), .A2(new_n547), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n624), .A2(new_n591), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT30), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n750), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n748), .A2(new_n547), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n752), .A2(new_n753), .A3(new_n754), .A4(new_n571), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n748), .ZN(new_n757));
  AOI21_X1  g0557(.A(G179), .B1(new_n564), .B2(new_n569), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n549), .A2(new_n757), .A3(new_n598), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT31), .B1(new_n760), .B2(new_n713), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n751), .B2(new_n755), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT31), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n763), .A2(new_n764), .A3(new_n735), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n747), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n728), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n696), .A2(new_n700), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n730), .B1(new_n720), .B2(new_n721), .ZN(new_n771));
  INV_X1    g0571(.A(new_n704), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n723), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT93), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n775), .A3(new_n735), .ZN(new_n776));
  INV_X1    g0576(.A(new_n735), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT93), .B1(new_n706), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT29), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n691), .B1(new_n702), .B2(new_n705), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n699), .A2(new_n695), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(KEYINPUT94), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n694), .A2(KEYINPUT26), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT94), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n699), .A2(new_n785), .A3(new_n695), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n713), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT29), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n769), .B1(new_n780), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n746), .B1(new_n790), .B2(G1), .ZN(G364));
  NOR2_X1   g0591(.A1(new_n288), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n296), .B1(new_n792), .B2(G45), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n741), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n733), .B2(new_n728), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n728), .B2(new_n733), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n261), .A2(new_n210), .ZN(new_n798));
  INV_X1    g0598(.A(G355), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n798), .A2(new_n799), .B1(G116), .B2(new_n210), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n363), .A2(new_n365), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n740), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n224), .A2(G45), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n241), .B2(G45), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n800), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n282), .B1(G20), .B2(new_n313), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n277), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n795), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(G20), .A2(G179), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n813), .A2(G190), .A3(G200), .ZN(new_n814));
  INV_X1    g0614(.A(G326), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n337), .A2(G179), .A3(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n277), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n517), .B1(new_n814), .B2(new_n815), .C1(new_n817), .C2(new_n545), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n277), .A2(G179), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n819), .A2(G190), .A3(G200), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n818), .B1(G303), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G190), .A2(G200), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n812), .A2(new_n243), .A3(G190), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT33), .B(G317), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n825), .A2(G311), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G322), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n813), .A2(G190), .A3(new_n243), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n822), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n819), .A2(new_n337), .A3(G200), .ZN(new_n832));
  INV_X1    g0632(.A(G283), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n819), .A2(new_n823), .ZN(new_n834));
  INV_X1    g0634(.A(G329), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n832), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT96), .Z(new_n837));
  NOR2_X1   g0637(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n838), .A2(KEYINPUT97), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(KEYINPUT97), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n814), .A2(new_n202), .B1(new_n824), .B2(new_n213), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n517), .B(new_n841), .C1(G68), .C2(new_n826), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n820), .A2(new_n518), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n832), .A2(new_n206), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT32), .ZN(new_n845));
  INV_X1    g0645(.A(G159), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n834), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT95), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n830), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G58), .ZN(new_n851));
  INV_X1    g0651(.A(new_n847), .ZN(new_n852));
  INV_X1    g0652(.A(new_n817), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n852), .A2(KEYINPUT32), .B1(new_n853), .B2(G97), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n842), .A2(new_n848), .A3(new_n851), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n839), .A2(new_n840), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n811), .B1(new_n856), .B2(new_n806), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n809), .B(KEYINPUT98), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n733), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n797), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G396));
  INV_X1    g0661(.A(new_n808), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n807), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n801), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n853), .A2(G58), .B1(new_n821), .B2(G50), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n865), .B1(new_n346), .B2(new_n832), .C1(new_n866), .C2(new_n834), .ZN(new_n867));
  INV_X1    g0667(.A(new_n814), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n868), .A2(G137), .B1(new_n825), .B2(G159), .ZN(new_n869));
  INV_X1    g0669(.A(new_n826), .ZN(new_n870));
  INV_X1    g0670(.A(new_n850), .ZN(new_n871));
  INV_X1    g0671(.A(G143), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n869), .B1(new_n274), .B2(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT34), .Z(new_n874));
  AOI211_X1 g0674(.A(new_n864), .B(new_n867), .C1(new_n874), .C2(KEYINPUT100), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n874), .A2(KEYINPUT100), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n868), .A2(G303), .B1(new_n825), .B2(G116), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n833), .B2(new_n870), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT99), .ZN(new_n879));
  INV_X1    g0679(.A(G311), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n517), .B1(new_n834), .B2(new_n880), .C1(new_n830), .C2(new_n545), .ZN(new_n881));
  INV_X1    g0681(.A(new_n832), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(G87), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n205), .B2(new_n817), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n881), .B(new_n884), .C1(G107), .C2(new_n821), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n875), .A2(new_n876), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n795), .B1(G77), .B2(new_n863), .C1(new_n886), .C2(new_n807), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT101), .Z(new_n888));
  INV_X1    g0688(.A(new_n334), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n339), .B1(new_n889), .B2(new_n725), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n342), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n342), .A2(new_n713), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n888), .B1(new_n808), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n776), .A2(new_n778), .A3(new_n894), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n892), .B1(new_n890), .B2(new_n342), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n774), .A2(new_n735), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n769), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n898), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n795), .B1(new_n900), .B2(new_n768), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n895), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(G384));
  NOR3_X1   g0703(.A1(new_n213), .A2(new_n224), .A3(new_n347), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n202), .B2(G68), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n905), .A2(new_n296), .A3(G13), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT102), .Z(new_n907));
  INV_X1    g0707(.A(KEYINPUT36), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n604), .A2(new_n605), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n503), .B(new_n223), .C1(new_n910), .C2(KEYINPUT35), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(KEYINPUT35), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n907), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n908), .B2(new_n912), .ZN(new_n914));
  INV_X1    g0714(.A(new_n690), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n493), .B1(KEYINPUT29), .B2(new_n788), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(new_n780), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n368), .A2(new_n287), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n421), .A2(KEYINPUT16), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n381), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n711), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n425), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT37), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n380), .B(new_n402), .C1(new_n368), .C2(new_n376), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n921), .B2(new_n922), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n921), .A2(new_n411), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n377), .A2(new_n381), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n411), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n922), .ZN(new_n932));
  AND4_X1   g0732(.A1(new_n925), .A2(new_n931), .A3(new_n932), .A4(new_n404), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n924), .B(KEYINPUT38), .C1(new_n929), .C2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n932), .A3(new_n404), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT37), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n926), .B1(new_n930), .B2(new_n411), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n925), .A3(new_n932), .ZN(new_n938));
  INV_X1    g0738(.A(new_n932), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n936), .A2(new_n938), .B1(new_n425), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n934), .B1(new_n940), .B2(KEYINPUT38), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n489), .A2(new_n486), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n488), .B1(new_n487), .B2(G169), .ZN(new_n945));
  OAI211_X1 g0745(.A(KEYINPUT103), .B(new_n491), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT103), .B1(new_n490), .B2(new_n491), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n713), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n924), .B1(new_n929), .B2(new_n933), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT38), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(KEYINPUT39), .A3(new_n934), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n943), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n934), .ZN(new_n956));
  INV_X1    g0756(.A(new_n948), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n454), .A2(new_n725), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n454), .B2(new_n481), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n946), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n490), .B1(new_n473), .B2(new_n482), .ZN(new_n961));
  INV_X1    g0761(.A(new_n958), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n961), .A2(KEYINPUT104), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT104), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n944), .A2(new_n945), .ZN(new_n965));
  AOI221_X4 g0765(.A(new_n472), .B1(new_n451), .B2(new_n453), .C1(new_n480), .C2(new_n468), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT79), .B1(new_n481), .B2(new_n454), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n964), .B1(new_n968), .B2(new_n958), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n960), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n706), .A2(new_n777), .A3(new_n894), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n956), .B(new_n970), .C1(new_n971), .C2(new_n892), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n685), .A2(new_n922), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n955), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT105), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT104), .B1(new_n961), .B2(new_n962), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n968), .A2(new_n964), .A3(new_n958), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n977), .A2(new_n978), .B1(new_n949), .B2(new_n959), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n898), .B2(new_n893), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n973), .B1(new_n980), .B2(new_n956), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT105), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n982), .A3(new_n955), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n976), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n918), .B(new_n984), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n763), .A2(new_n764), .A3(new_n725), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n761), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n747), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n941), .A2(new_n970), .A3(new_n897), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT40), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n979), .A2(new_n894), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT40), .B1(new_n953), .B2(new_n934), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n992), .A3(new_n988), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n494), .A2(new_n988), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n728), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n985), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n296), .B2(new_n792), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n985), .A2(new_n997), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n914), .B1(new_n999), .B2(new_n1000), .ZN(G367));
  INV_X1    g0801(.A(new_n795), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n802), .A2(new_n234), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n810), .B1(new_n740), .B2(new_n652), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n657), .A2(new_n713), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n703), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n679), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n817), .A2(new_n346), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n870), .A2(new_n846), .B1(new_n830), .B2(new_n274), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G58), .C2(new_n821), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n261), .B1(new_n832), .B2(new_n213), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT113), .Z(new_n1013));
  INV_X1    g0813(.A(G137), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n834), .A2(new_n1014), .B1(new_n824), .B2(new_n202), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G143), .B2(new_n868), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n850), .A2(G303), .B1(G311), .B2(new_n868), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT112), .ZN(new_n1019));
  INV_X1    g0819(.A(G317), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n834), .A2(new_n1020), .B1(new_n824), .B2(new_n833), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n817), .A2(new_n206), .B1(new_n832), .B2(new_n205), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G294), .C2(new_n826), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT46), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n820), .B2(new_n503), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n821), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1023), .A2(new_n864), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1017), .B1(new_n1019), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT114), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT47), .Z(new_n1030));
  OAI221_X1 g0830(.A(new_n1005), .B1(new_n858), .B2(new_n1008), .C1(new_n1030), .C2(new_n807), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT115), .Z(new_n1032));
  OAI211_X1 g0832(.A(new_n618), .B(new_n626), .C1(new_n617), .C2(new_n735), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n698), .A2(new_n625), .A3(new_n777), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n738), .A2(new_n736), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT45), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n738), .A2(new_n736), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1035), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT44), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT44), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1043), .B(new_n1035), .C1(new_n738), .C2(new_n736), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1038), .A2(new_n1039), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n734), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1035), .B1(new_n738), .B2(new_n736), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT44), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1036), .B(new_n1037), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n734), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1047), .A2(new_n1051), .B1(KEYINPUT110), .B2(new_n1045), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1045), .A2(KEYINPUT110), .A3(new_n734), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n733), .A2(new_n728), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n561), .A2(new_n737), .B1(new_n1054), .B2(KEYINPUT111), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n737), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n714), .B(new_n1056), .C1(new_n724), .C2(new_n726), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1054), .A2(KEYINPUT111), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1055), .B(new_n1057), .C1(KEYINPUT111), .C2(new_n1054), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1053), .A2(new_n790), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n790), .B1(new_n1052), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n741), .B(new_n1065), .Z(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n794), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n734), .A2(new_n1041), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n561), .A2(KEYINPUT42), .A3(new_n737), .A4(new_n1035), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT42), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n738), .B2(new_n1041), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n626), .B1(new_n722), .B2(new_n1033), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1070), .A2(new_n1072), .B1(new_n1073), .B2(new_n735), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT108), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1008), .B(KEYINPUT43), .Z(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  OR3_X1    g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1075), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT107), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1074), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1081), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1069), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1080), .A2(new_n1085), .A3(new_n1069), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1032), .B1(new_n1068), .B2(new_n1089), .ZN(G387));
  OAI22_X1  g0890(.A1(new_n798), .A2(new_n743), .B1(G107), .B2(new_n210), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n231), .A2(G45), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n743), .B(new_n245), .C1(new_n346), .C2(new_n331), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT50), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n279), .B2(G50), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n378), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1097), .A2(new_n740), .A3(new_n801), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1091), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n795), .B1(new_n1099), .B2(new_n810), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n870), .A2(new_n279), .B1(new_n824), .B2(new_n346), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G97), .B2(new_n882), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n830), .A2(new_n202), .B1(new_n834), .B2(new_n274), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G159), .B2(new_n868), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n820), .A2(new_n213), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n652), .B2(new_n853), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1102), .A2(new_n1104), .A3(new_n801), .A4(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n853), .A2(G283), .B1(new_n821), .B2(G294), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n825), .A2(G303), .B1(G311), .B2(new_n826), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n829), .B2(new_n814), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G317), .B2(new_n850), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT116), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1108), .B1(new_n1113), .B2(KEYINPUT48), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(KEYINPUT48), .B2(new_n1113), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT117), .Z(new_n1116));
  INV_X1    g0916(.A(KEYINPUT49), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n832), .A2(new_n503), .B1(new_n834), .B2(new_n815), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n801), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1107), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1100), .B1(new_n1122), .B2(new_n806), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n727), .B2(new_n858), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1062), .A2(new_n794), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n790), .A2(new_n1062), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n790), .A2(new_n1062), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n741), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1124), .B(new_n1125), .C1(new_n1126), .C2(new_n1128), .ZN(G393));
  NAND2_X1  g0929(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n742), .B1(new_n1130), .B2(new_n1127), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1052), .B2(new_n1063), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1047), .A2(new_n1051), .A3(new_n794), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n830), .A2(new_n846), .B1(new_n814), .B2(new_n274), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT51), .Z(new_n1135));
  AOI22_X1  g0935(.A1(new_n825), .A2(new_n378), .B1(G50), .B2(new_n826), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n872), .B2(new_n834), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n883), .B1(new_n346), .B2(new_n820), .C1(new_n331), .C2(new_n817), .ZN(new_n1138));
  OR4_X1    g0938(.A1(new_n864), .A2(new_n1135), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n517), .B1(new_n834), .B2(new_n829), .C1(new_n545), .C2(new_n824), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n844), .B(new_n1140), .C1(G283), .C2(new_n821), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n817), .A2(new_n503), .B1(new_n870), .B2(new_n567), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT118), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n830), .A2(new_n880), .B1(new_n814), .B2(new_n1020), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT52), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1141), .A2(new_n1144), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n807), .B1(new_n1139), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n802), .A2(new_n238), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n810), .B1(G97), .B2(new_n740), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1002), .B(new_n1149), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1035), .B2(new_n809), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1133), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1132), .A2(new_n1154), .ZN(G390));
  AND3_X1   g0955(.A1(new_n953), .A2(KEYINPUT39), .A3(new_n934), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n925), .B1(new_n937), .B2(new_n932), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(new_n933), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n425), .A2(new_n939), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n952), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT39), .B1(new_n1160), .B2(new_n934), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n980), .A2(new_n950), .B1(new_n1156), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n950), .B1(new_n1160), .B2(new_n934), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n892), .B1(new_n788), .B2(new_n891), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n979), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n767), .A2(new_n728), .A3(new_n897), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1166), .A2(new_n979), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1162), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(G330), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n747), .B2(new_n987), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n991), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n808), .B1(new_n1156), .B2(new_n1161), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n795), .B1(new_n378), .B2(new_n863), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n261), .B(new_n843), .C1(G283), .C2(new_n868), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n830), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1177), .A2(G116), .B1(new_n825), .B2(G97), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n834), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1179), .A2(G294), .B1(G107), .B2(new_n826), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n853), .A2(G77), .B1(new_n882), .B2(G68), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1176), .A2(new_n1178), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n517), .B1(new_n1179), .B2(G125), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n202), .B2(new_n832), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT120), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n820), .A2(new_n274), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT53), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n870), .A2(new_n1014), .B1(new_n830), .B2(new_n866), .ZN(new_n1188));
  INV_X1    g0988(.A(G128), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT54), .B(G143), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n814), .A2(new_n1189), .B1(new_n824), .B2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1187), .B(new_n1192), .C1(new_n846), .C2(new_n817), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1182), .B1(new_n1185), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1175), .B1(new_n1194), .B2(new_n806), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1173), .A2(new_n794), .B1(new_n1174), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n780), .A2(new_n494), .A3(new_n789), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n494), .A2(new_n1170), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n690), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT119), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n917), .A2(KEYINPUT119), .A3(new_n1198), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n971), .A2(new_n892), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n991), .A2(new_n1170), .B1(new_n1166), .B2(new_n979), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1164), .B1(new_n979), .B2(new_n1166), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n970), .B1(new_n1170), .B2(new_n897), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1203), .A2(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1201), .A2(new_n1202), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n741), .B1(new_n1208), .B2(new_n1173), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1172), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1162), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1201), .A2(new_n1202), .A3(new_n1207), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1196), .B1(new_n1209), .B2(new_n1214), .ZN(G378));
  NAND2_X1  g1015(.A1(new_n310), .A2(new_n315), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n305), .A2(new_n306), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n299), .A3(new_n922), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n299), .A2(new_n922), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n305), .A2(new_n306), .A3(new_n1216), .A4(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n808), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n795), .B1(G50), .B2(new_n863), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n868), .A2(G125), .B1(G132), .B2(new_n826), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n1189), .B2(new_n830), .C1(new_n1014), .C2(new_n824), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n817), .A2(new_n274), .B1(new_n820), .B2(new_n1190), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n882), .A2(G159), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n1179), .C2(G124), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G283), .A2(new_n1179), .B1(new_n825), .B2(new_n652), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n503), .B2(new_n814), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n870), .A2(new_n205), .B1(new_n830), .B2(new_n206), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n832), .A2(new_n345), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1240), .A2(new_n1009), .A3(new_n1105), .A4(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1239), .A2(new_n1242), .A3(new_n244), .A4(new_n864), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(KEYINPUT58), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G50), .B1(new_n258), .B2(new_n244), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n801), .B2(G41), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(KEYINPUT58), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1236), .A2(new_n1245), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1226), .B1(new_n1249), .B2(new_n806), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1225), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1224), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n994), .B2(G330), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1169), .B(new_n1224), .C1(new_n990), .C2(new_n993), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n975), .A2(KEYINPUT105), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n982), .B1(new_n981), .B2(new_n955), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1253), .A2(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n970), .A2(new_n897), .A3(new_n988), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1258), .A2(new_n992), .B1(new_n989), .B2(KEYINPUT40), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1224), .B1(new_n1259), .B2(new_n1169), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n994), .A2(G330), .A3(new_n1252), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n983), .A4(new_n976), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1251), .B1(new_n1263), .B2(new_n793), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1257), .A2(KEYINPUT57), .A3(new_n1262), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1207), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1266), .B1(new_n1212), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n742), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT57), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1173), .B2(new_n1207), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1272), .B2(new_n1263), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1264), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(G375));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1267), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1067), .A3(new_n1213), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(KEYINPUT121), .Z(new_n1278));
  NOR2_X1   g1078(.A1(new_n871), .A2(new_n1014), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1241), .B1(G50), .B2(new_n853), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n846), .B2(new_n820), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n870), .A2(new_n1190), .B1(new_n834), .B2(new_n1189), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n814), .A2(new_n866), .B1(new_n824), .B2(new_n274), .ZN(new_n1283));
  NOR4_X1   g1083(.A1(new_n1279), .A2(new_n1281), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n830), .A2(new_n833), .B1(new_n824), .B2(new_n206), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n261), .B1(G116), .B2(new_n826), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n1286), .B1(new_n331), .B2(new_n832), .C1(new_n326), .C2(new_n817), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1285), .B(new_n1287), .C1(G294), .C2(new_n868), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n820), .A2(new_n205), .B1(new_n834), .B2(new_n567), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(KEYINPUT122), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1284), .A2(new_n801), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n795), .B1(G68), .B2(new_n863), .C1(new_n1291), .C2(new_n807), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n979), .B2(new_n808), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1207), .B2(new_n794), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1278), .A2(new_n1294), .ZN(G381));
  INV_X1    g1095(.A(G381), .ZN(new_n1296));
  INV_X1    g1096(.A(G378), .ZN(new_n1297));
  INV_X1    g1097(.A(G390), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n902), .ZN(new_n1299));
  NOR4_X1   g1099(.A1(new_n1299), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1296), .A2(new_n1297), .A3(new_n1274), .A4(new_n1300), .ZN(G407));
  NAND3_X1  g1101(.A1(new_n1274), .A2(new_n712), .A3(new_n1297), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(G407), .A2(G213), .A3(new_n1302), .ZN(G409));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(G393), .B(new_n860), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1088), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1307), .A2(new_n1086), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1045), .A2(KEYINPUT110), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n734), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1309), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1127), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1312), .A2(new_n1313), .A3(new_n1053), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1066), .B1(new_n1314), .B2(new_n790), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1308), .B1(new_n1315), .B2(new_n794), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G390), .B1(new_n1316), .B2(new_n1032), .ZN(new_n1317));
  OAI211_X1 g1117(.A(G390), .B(new_n1032), .C1(new_n1068), .C2(new_n1089), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1306), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G387), .A2(new_n1298), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(new_n1305), .A3(new_n1318), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT62), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT124), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n712), .A2(G213), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1251), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1329), .B2(new_n794), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT57), .B1(new_n1329), .B2(new_n1268), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1257), .A2(new_n1262), .A3(KEYINPUT57), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n741), .B1(new_n1332), .B2(new_n1272), .ZN(new_n1333));
  OAI211_X1 g1133(.A(G378), .B(new_n1330), .C1(new_n1331), .C2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT123), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1268), .A2(KEYINPUT57), .A3(new_n1262), .A4(new_n1257), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(new_n1273), .A3(new_n741), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1338), .A2(KEYINPUT123), .A3(G378), .A4(new_n1330), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1329), .A2(new_n1067), .A3(new_n1268), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G378), .B1(new_n1330), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1327), .B1(new_n1340), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1213), .A2(KEYINPUT60), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1345), .A2(new_n1276), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1271), .A2(new_n1267), .A3(KEYINPUT60), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n741), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1294), .B1(new_n1346), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n902), .ZN(new_n1350));
  OAI211_X1 g1150(.A(G384), .B(new_n1294), .C1(new_n1346), .C2(new_n1348), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1325), .B1(new_n1344), .B2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1342), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1355));
  NOR4_X1   g1155(.A1(new_n1355), .A2(new_n1352), .A3(KEYINPUT124), .A4(new_n1327), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1324), .B1(new_n1354), .B2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1327), .A2(G2897), .ZN(new_n1358));
  XNOR2_X1  g1158(.A(new_n1358), .B(KEYINPUT125), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1350), .A2(new_n1351), .A3(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1359), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1362), .B1(new_n1355), .B2(new_n1327), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT61), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1324), .B1(new_n1344), .B2(new_n1353), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1323), .B1(new_n1357), .B2(new_n1367), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1344), .A2(KEYINPUT63), .A3(new_n1353), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1320), .A2(new_n1364), .A3(new_n1322), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(new_n1370), .B(KEYINPUT126), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1369), .A2(new_n1371), .A3(new_n1363), .ZN(new_n1372));
  NOR2_X1   g1172(.A1(new_n1354), .A2(new_n1356), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT63), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1372), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1304), .B1(new_n1368), .B2(new_n1375), .ZN(new_n1376));
  AOI21_X1  g1176(.A(KEYINPUT123), .B1(new_n1274), .B2(G378), .ZN(new_n1377));
  NOR2_X1   g1177(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1343), .B1(new_n1377), .B2(new_n1378), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1379), .A2(new_n1353), .A3(new_n1326), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1380), .A2(KEYINPUT124), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1344), .A2(new_n1325), .A3(new_n1353), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1381), .A2(new_n1374), .A3(new_n1382), .ZN(new_n1383));
  AND2_X1   g1183(.A1(new_n1371), .A2(new_n1363), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1383), .A2(new_n1369), .A3(new_n1384), .ZN(new_n1385));
  NOR3_X1   g1185(.A1(new_n1355), .A2(new_n1352), .A3(new_n1327), .ZN(new_n1386));
  OAI211_X1 g1186(.A(new_n1364), .B(new_n1363), .C1(new_n1386), .C2(new_n1324), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1387), .B1(new_n1388), .B2(new_n1324), .ZN(new_n1389));
  OAI211_X1 g1189(.A(KEYINPUT127), .B(new_n1385), .C1(new_n1389), .C2(new_n1323), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1376), .A2(new_n1390), .ZN(G405));
  OAI21_X1  g1191(.A(new_n1340), .B1(G378), .B2(new_n1274), .ZN(new_n1392));
  XNOR2_X1  g1192(.A(new_n1392), .B(new_n1352), .ZN(new_n1393));
  XNOR2_X1  g1193(.A(new_n1393), .B(new_n1323), .ZN(G402));
endmodule


