//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT70), .B(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(KEYINPUT16), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n192), .B(G146), .C1(KEYINPUT16), .C2(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n200), .A2(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n201), .B(new_n203), .C1(new_n204), .C2(KEYINPUT23), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT24), .B(G110), .Z(new_n206));
  XNOR2_X1  g020(.A(G119), .B(G128), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n205), .A2(G110), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n199), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT72), .B(G110), .Z(new_n210));
  OAI22_X1  g024(.A1(new_n205), .A2(new_n210), .B1(new_n206), .B2(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n191), .A2(new_n196), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n198), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(KEYINPUT73), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G137), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n209), .A2(new_n213), .A3(new_n219), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n188), .A3(new_n222), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n190), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n189), .A2(G902), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n223), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n231));
  NOR2_X1   g045(.A1(G472), .A2(G902), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT31), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(new_n239), .A3(new_n242), .A4(new_n237), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n196), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT64), .B(G143), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G146), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT64), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n256), .A3(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n196), .A2(G143), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n249), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n244), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n238), .A2(G134), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n235), .A2(G137), .ZN(new_n262));
  OAI21_X1  g076(.A(G131), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n243), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n202), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n255), .A2(G143), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n253), .A2(KEYINPUT64), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n196), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n268), .B2(new_n246), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n257), .A2(new_n258), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n264), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n200), .A2(G116), .ZN(new_n273));
  INV_X1    g087(.A(G116), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G119), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT2), .B(G113), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n260), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT26), .B(G101), .Z(new_n283));
  INV_X1    g097(.A(G237), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(new_n215), .A3(G210), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n241), .A2(new_n243), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n254), .A2(new_n256), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n245), .B1(new_n291), .B2(new_n196), .ZN(new_n292));
  INV_X1    g106(.A(new_n251), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n259), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n243), .A2(new_n263), .ZN(new_n296));
  INV_X1    g110(.A(new_n265), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n248), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n258), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n247), .B2(G146), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n270), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n296), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT30), .B1(new_n295), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n260), .A2(new_n272), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n279), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n278), .B(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT66), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n260), .A2(new_n272), .A3(new_n304), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n304), .B1(new_n260), .B2(new_n272), .ZN(new_n311));
  OAI211_X1 g125(.A(KEYINPUT66), .B(new_n308), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n233), .B(new_n289), .C1(new_n309), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n308), .B1(new_n295), .B2(new_n302), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(new_n281), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n281), .A2(new_n315), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n288), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT68), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT68), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n322), .B(new_n288), .C1(new_n317), .C2(new_n319), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n314), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n312), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n233), .B1(new_n328), .B2(new_n289), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n232), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT32), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n330), .A2(KEYINPUT69), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT69), .B1(new_n330), .B2(new_n331), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(KEYINPUT32), .B(new_n232), .C1(new_n324), .C2(new_n329), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n280), .B1(new_n260), .B2(new_n272), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT28), .B1(new_n282), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n288), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n318), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n281), .B1(new_n309), .B2(new_n313), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(new_n288), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n188), .B1(new_n339), .B2(new_n340), .ZN(new_n344));
  OAI21_X1  g158(.A(G472), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n335), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n231), .B1(new_n334), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n330), .A2(new_n331), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n330), .A2(KEYINPUT69), .A3(new_n331), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n346), .A3(new_n231), .A4(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n230), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G469), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n257), .A2(new_n258), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT1), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n291), .B2(new_n196), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n359), .B2(new_n202), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(KEYINPUT75), .B(new_n357), .C1(new_n359), .C2(new_n202), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n301), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G104), .ZN(new_n369));
  INV_X1    g183(.A(G101), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(G107), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n366), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n365), .A2(G107), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n368), .A2(G104), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT76), .B1(new_n364), .B2(new_n377), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n356), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n298), .A2(new_n301), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n382), .A2(new_n356), .A3(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT74), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G101), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n387), .B2(new_n372), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT4), .B1(new_n386), .B2(G101), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n384), .B1(new_n390), .B2(new_n294), .ZN(new_n391));
  INV_X1    g205(.A(new_n294), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n392), .B(KEYINPUT74), .C1(new_n388), .C2(new_n389), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n383), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n380), .A2(new_n290), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G110), .B(G140), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n215), .A2(G227), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n381), .A2(new_n377), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n378), .B2(new_n379), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT12), .A3(new_n244), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT12), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n300), .B1(G128), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n301), .B1(new_n407), .B2(KEYINPUT75), .ZN(new_n408));
  INV_X1    g222(.A(new_n363), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n377), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n377), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n401), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n405), .B1(new_n414), .B2(new_n290), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n400), .B1(new_n404), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n380), .A2(new_n394), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n244), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n399), .B1(new_n418), .B2(new_n395), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n355), .B(new_n188), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n395), .A3(new_n399), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n391), .A2(new_n393), .ZN(new_n422));
  INV_X1    g236(.A(new_n383), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n413), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(new_n356), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n415), .A2(new_n404), .B1(new_n426), .B2(new_n290), .ZN(new_n427));
  OAI211_X1 g241(.A(G469), .B(new_n421), .C1(new_n427), .C2(new_n399), .ZN(new_n428));
  INV_X1    g242(.A(G902), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n355), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n420), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT9), .B(G234), .ZN(new_n433));
  OAI21_X1  g247(.A(G221), .B1(new_n433), .B2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(G475), .A2(G902), .ZN(new_n436));
  XNOR2_X1  g250(.A(G113), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(new_n365), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n284), .A2(new_n215), .A3(G214), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n254), .A3(new_n256), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n284), .A2(new_n215), .A3(G143), .A4(G214), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G131), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n242), .B1(new_n440), .B2(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n198), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n191), .B(KEYINPUT19), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n196), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(KEYINPUT88), .A3(new_n196), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n191), .B(new_n196), .ZN(new_n453));
  NAND2_X1  g267(.A1(KEYINPUT18), .A2(G131), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT84), .B1(new_n442), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n457));
  AOI211_X1 g271(.A(new_n457), .B(new_n454), .C1(new_n440), .C2(new_n441), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n453), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(KEYINPUT85), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n440), .A2(new_n441), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT86), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n452), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n456), .A2(new_n458), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT86), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n463), .B(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT87), .A4(new_n453), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n451), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT89), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n438), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n465), .A2(new_n469), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT89), .B1(new_n473), .B2(new_n451), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n465), .A2(new_n469), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n199), .B1(KEYINPUT17), .B2(new_n444), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n443), .A2(new_n444), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(KEYINPUT17), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n438), .B(KEYINPUT90), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n436), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT91), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n472), .B2(new_n474), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT20), .B1(new_n436), .B2(KEYINPUT92), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(KEYINPUT92), .B2(new_n436), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n490), .B(KEYINPUT20), .C1(new_n486), .C2(new_n436), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n476), .A2(new_n479), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(new_n438), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n429), .B1(new_n494), .B2(new_n481), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G475), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n215), .A2(G952), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(G234), .B2(G237), .ZN(new_n498));
  AOI211_X1 g312(.A(new_n215), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT21), .B(G898), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n274), .A2(G122), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n368), .B1(new_n503), .B2(KEYINPUT14), .ZN(new_n504));
  XNOR2_X1  g318(.A(G116), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n247), .A2(G128), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n202), .A2(G143), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n235), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n235), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n505), .B(new_n368), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n507), .A2(KEYINPUT13), .A3(new_n508), .ZN(new_n514));
  OAI21_X1  g328(.A(G134), .B1(new_n507), .B2(KEYINPUT13), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n509), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n433), .A2(new_n187), .A3(G953), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n518), .B(KEYINPUT93), .Z(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n519), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n516), .A3(new_n512), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(KEYINPUT94), .A3(new_n522), .ZN(new_n523));
  OR3_X1    g337(.A1(new_n517), .A2(KEYINPUT94), .A3(new_n519), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n188), .ZN(new_n525));
  INV_X1    g339(.A(G478), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n525), .B(new_n527), .Z(new_n528));
  NAND4_X1  g342(.A1(new_n492), .A2(new_n496), .A3(new_n502), .A4(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n435), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G210), .B1(G237), .B2(G902), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT80), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n273), .A2(new_n275), .A3(KEYINPUT5), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G113), .B1(new_n273), .B2(KEYINPUT5), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(KEYINPUT77), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n538));
  INV_X1    g352(.A(new_n536), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(new_n534), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n276), .A2(new_n279), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n533), .B(new_n376), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT77), .B1(new_n535), .B2(new_n536), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n538), .A3(new_n534), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT80), .B1(new_n546), .B2(new_n377), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n536), .B1(new_n534), .B2(KEYINPUT79), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(KEYINPUT79), .B2(new_n534), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n376), .A2(new_n542), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n550), .B1(new_n537), .B2(new_n540), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT78), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n308), .B1(new_n388), .B2(new_n389), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n550), .B(KEYINPUT78), .C1(new_n537), .C2(new_n540), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n558), .A2(new_n553), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n294), .A2(G125), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(G125), .B2(new_n381), .ZN(new_n563));
  INV_X1    g377(.A(G224), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G953), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(KEYINPUT7), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(KEYINPUT7), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n562), .B(new_n568), .C1(G125), .C2(new_n381), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n555), .A2(new_n561), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT81), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n429), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n574));
  INV_X1    g388(.A(new_n553), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(KEYINPUT6), .A3(new_n561), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT6), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n563), .B(new_n565), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n572), .B1(new_n571), .B2(new_n429), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n532), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n583), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(new_n531), .A3(new_n581), .A4(new_n573), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT82), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(G214), .B1(G237), .B2(G902), .ZN(new_n589));
  INV_X1    g403(.A(new_n582), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n590), .A2(KEYINPUT82), .A3(new_n531), .A4(new_n585), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT83), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT83), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n588), .A2(new_n594), .A3(new_n589), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n530), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n354), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n370), .ZN(G3));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n523), .A2(new_n524), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n520), .A2(KEYINPUT33), .A3(new_n522), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n601), .A2(G478), .A3(new_n188), .A4(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n525), .A2(new_n526), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n603), .B2(new_n604), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n492), .B2(new_n496), .ZN(new_n609));
  INV_X1    g423(.A(new_n589), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n584), .B2(new_n586), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n609), .A2(new_n502), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n435), .ZN(new_n613));
  INV_X1    g427(.A(G472), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n324), .A2(new_n329), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n615), .B2(new_n188), .ZN(new_n616));
  INV_X1    g430(.A(new_n330), .ZN(new_n617));
  INV_X1    g431(.A(new_n230), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  NAND2_X1  g436(.A1(new_n483), .A2(new_n484), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n485), .A2(new_n491), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n496), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n525), .B(new_n527), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n611), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n625), .A2(new_n627), .A3(new_n501), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n613), .A3(new_n619), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n616), .A2(new_n617), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n220), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n214), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n634), .A2(new_n229), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n228), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n530), .A2(new_n596), .A3(new_n632), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT96), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT37), .B(G110), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  NAND3_X1  g455(.A1(new_n350), .A2(new_n346), .A3(new_n351), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT71), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n352), .ZN(new_n644));
  AOI211_X1 g458(.A(new_n610), .B(new_n636), .C1(new_n586), .C2(new_n584), .ZN(new_n645));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n499), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n498), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n624), .A2(new_n496), .A3(new_n626), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n644), .A2(new_n613), .A3(new_n645), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  NAND2_X1  g467(.A1(new_n588), .A2(new_n591), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT38), .Z(new_n655));
  AND2_X1   g469(.A1(new_n492), .A2(new_n496), .ZN(new_n656));
  NOR4_X1   g470(.A1(new_n656), .A2(new_n610), .A3(new_n528), .A4(new_n637), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n342), .A2(new_n338), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n316), .A2(new_n281), .A3(new_n288), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n658), .A2(new_n429), .A3(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n334), .B(new_n335), .C1(new_n614), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n655), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n649), .B(KEYINPUT39), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n613), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT40), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n666), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n247), .B(KEYINPUT98), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G45));
  AND2_X1   g484(.A1(new_n609), .A2(new_n649), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n644), .A2(new_n613), .A3(new_n645), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  OR2_X1    g487(.A1(new_n416), .A2(new_n419), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n355), .B1(new_n674), .B2(new_n188), .ZN(new_n675));
  INV_X1    g489(.A(new_n434), .ZN(new_n676));
  INV_X1    g490(.A(new_n420), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n644), .A2(new_n612), .A3(new_n230), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NAND4_X1  g495(.A1(new_n644), .A2(new_n230), .A3(new_n628), .A4(new_n678), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  NOR2_X1   g497(.A1(new_n416), .A2(new_n419), .ZN(new_n684));
  INV_X1    g498(.A(new_n188), .ZN(new_n685));
  OAI21_X1  g499(.A(G469), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n645), .A2(new_n434), .A3(new_n420), .A4(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n529), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n644), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  NAND2_X1  g504(.A1(new_n492), .A2(new_n496), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n626), .A3(new_n611), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n686), .A2(new_n502), .A3(new_n434), .A4(new_n420), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n615), .A2(new_n188), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G472), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n232), .B(KEYINPUT99), .Z(new_n696));
  INV_X1    g510(.A(new_n329), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n320), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n314), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n698), .B1(new_n697), .B2(new_n320), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n696), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n695), .A2(new_n702), .A3(new_n230), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n692), .A2(new_n693), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(G122), .Z(G24));
  NAND2_X1  g519(.A1(new_n609), .A2(new_n649), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n695), .A2(new_n702), .A3(new_n637), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n686), .A2(new_n434), .A3(new_n420), .A4(new_n611), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n193), .ZN(G27));
  NAND2_X1  g524(.A1(new_n346), .A2(new_n348), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n609), .A2(new_n230), .A3(new_n649), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n428), .A2(KEYINPUT101), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n414), .A2(new_n405), .A3(new_n290), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT12), .B1(new_n403), .B2(new_n244), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n395), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n398), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT101), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n718), .A3(G469), .A4(new_n421), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n713), .A2(new_n420), .A3(new_n719), .A4(new_n431), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n676), .A2(new_n610), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n588), .B2(new_n591), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT42), .B1(new_n712), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n720), .A2(new_n723), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n726), .B(new_n230), .C1(new_n347), .C2(new_n353), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n706), .A2(KEYINPUT42), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(KEYINPUT102), .B(new_n725), .C1(new_n727), .C2(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n242), .ZN(G33));
  NOR2_X1   g548(.A1(new_n727), .A2(new_n650), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n235), .ZN(G36));
  INV_X1    g550(.A(new_n608), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n656), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n632), .A2(new_n636), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(KEYINPUT44), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n654), .A2(new_n589), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n400), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n716), .A2(new_n398), .B1(new_n750), .B2(new_n418), .ZN(new_n751));
  OAI21_X1  g565(.A(G469), .B1(new_n751), .B2(KEYINPUT45), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n717), .A2(KEYINPUT45), .A3(new_n421), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n430), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT103), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n677), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n434), .A3(new_n663), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n749), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n238), .ZN(G39));
  NOR4_X1   g578(.A1(new_n644), .A2(new_n230), .A3(new_n706), .A4(new_n747), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n761), .A2(new_n434), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n434), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(G140), .Z(G42));
  NOR2_X1   g586(.A1(new_n675), .A2(new_n677), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT104), .Z(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT49), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n661), .A2(new_n618), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n776), .A2(new_n655), .A3(new_n722), .A4(new_n738), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n704), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n679), .A2(new_n682), .A3(new_n689), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n707), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n671), .A2(new_n726), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n727), .B2(new_n650), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n528), .A2(KEYINPUT106), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT106), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n626), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n637), .A3(new_n649), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n747), .A2(new_n789), .A3(new_n625), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n644), .A2(new_n790), .A3(new_n613), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT107), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n644), .A2(new_n790), .A3(new_n793), .A4(new_n613), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n780), .A2(new_n784), .A3(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n609), .A2(new_n502), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n596), .A3(new_n613), .A4(new_n619), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n354), .B2(new_n597), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT105), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT105), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n798), .B(new_n801), .C1(new_n354), .C2(new_n597), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n691), .A2(new_n788), .A3(new_n501), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n596), .A2(new_n803), .A3(new_n613), .A4(new_n619), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n638), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n800), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n796), .A2(new_n807), .A3(new_n733), .ZN(new_n808));
  INV_X1    g622(.A(new_n645), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n435), .B(new_n809), .C1(new_n643), .C2(new_n352), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n709), .B1(new_n810), .B2(new_n651), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n649), .B(KEYINPUT108), .Z(new_n813));
  NAND2_X1  g627(.A1(new_n636), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT109), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(new_n434), .ZN(new_n816));
  INV_X1    g630(.A(new_n692), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n661), .A4(new_n720), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n811), .A2(new_n812), .A3(new_n672), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n671), .A2(new_n678), .A3(new_n611), .A4(new_n781), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n652), .A2(new_n672), .A3(new_n820), .A4(new_n818), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n808), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n783), .B1(new_n792), .B2(new_n794), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n805), .B1(new_n799), .B2(KEYINPUT105), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n802), .A3(new_n827), .A4(new_n780), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n652), .A2(new_n820), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT53), .B1(new_n829), .B2(KEYINPUT52), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n828), .A2(new_n823), .A3(new_n733), .A4(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n796), .A2(new_n807), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(KEYINPUT52), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n729), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(new_n824), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n828), .A2(new_n823), .A3(new_n733), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(KEYINPUT53), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(KEYINPUT110), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n843), .B(KEYINPUT54), .C1(new_n825), .C2(new_n831), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n842), .B1(new_n841), .B2(new_n844), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n739), .A2(new_n498), .A3(new_n740), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n703), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n611), .A3(new_n678), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT115), .Z(new_n851));
  NAND2_X1  g665(.A1(new_n678), .A2(new_n748), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n648), .A3(new_n776), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n497), .B1(new_n855), .B2(new_n609), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT48), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n854), .A2(new_n848), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n711), .A2(new_n230), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n857), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n854), .A2(new_n848), .A3(KEYINPUT48), .A4(new_n859), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n847), .B1(new_n851), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n861), .A2(new_n862), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n850), .B(KEYINPUT115), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT116), .A4(new_n856), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n691), .A2(new_n737), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n855), .A2(new_n868), .B1(new_n858), .B2(new_n781), .ZN(new_n869));
  INV_X1    g683(.A(new_n703), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n741), .A2(new_n498), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n773), .A2(new_n434), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n655), .A2(new_n589), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT50), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND4_X1   g689(.A1(KEYINPUT50), .A2(new_n849), .A3(new_n678), .A4(new_n874), .ZN(new_n876));
  OAI211_X1 g690(.A(KEYINPUT51), .B(new_n869), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n774), .A2(KEYINPUT112), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n774), .A2(KEYINPUT112), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n676), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n769), .A2(new_n770), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n871), .A2(new_n747), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n864), .A2(new_n867), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n882), .A2(KEYINPUT113), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT113), .B1(new_n882), .B2(new_n883), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n869), .B1(new_n875), .B2(new_n876), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n885), .B1(new_n889), .B2(KEYINPUT51), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n845), .A2(new_n846), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(G952), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n215), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT117), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n778), .B1(new_n891), .B2(new_n894), .ZN(G75));
  OAI21_X1  g709(.A(new_n837), .B1(new_n839), .B2(KEYINPUT53), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n896), .A2(new_n685), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n532), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n577), .A2(new_n579), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT118), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n580), .B(KEYINPUT55), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n898), .B2(new_n899), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n215), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  NAND2_X1  g721(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n840), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n430), .B(KEYINPUT57), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n684), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n896), .A2(new_n685), .A3(new_n755), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT120), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n896), .A2(new_n916), .A3(new_n685), .A4(new_n755), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n911), .B2(new_n912), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n906), .B1(new_n913), .B2(new_n919), .ZN(G54));
  NAND3_X1  g734(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n486), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT121), .B1(new_n921), .B2(new_n486), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n906), .B1(new_n921), .B2(new_n486), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(G60));
  AND2_X1   g739(.A1(new_n601), .A2(new_n602), .ZN(new_n926));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n909), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(G952), .B2(new_n215), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n845), .B2(new_n846), .ZN(new_n932));
  INV_X1    g746(.A(new_n926), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT60), .Z(new_n936));
  AOI21_X1  g750(.A(new_n223), .B1(new_n896), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n906), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT61), .B1(new_n938), .B2(KEYINPUT122), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n896), .A2(new_n634), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G66));
  OAI21_X1  g756(.A(G953), .B1(new_n500), .B2(new_n564), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n827), .A2(new_n802), .A3(new_n780), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n901), .B1(G898), .B2(new_n215), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT123), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G69));
  XNOR2_X1  g762(.A(new_n306), .B(new_n446), .ZN(new_n949));
  NAND2_X1  g763(.A1(G900), .A2(G953), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n811), .A2(new_n672), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT124), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n771), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n733), .A2(new_n735), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n762), .A2(new_n692), .A3(new_n859), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n763), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n949), .B(new_n950), .C1(new_n957), .C2(G953), .ZN(new_n958));
  INV_X1    g772(.A(new_n952), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n668), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n788), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n609), .B1(new_n656), .B2(new_n963), .ZN(new_n964));
  OR4_X1    g778(.A1(new_n354), .A2(new_n664), .A3(new_n747), .A4(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n749), .B2(new_n762), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(KEYINPUT125), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(KEYINPUT125), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n771), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(G953), .B1(new_n962), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n958), .B1(new_n970), .B2(new_n949), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n215), .B1(G227), .B2(G900), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n972), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n974), .B(new_n958), .C1(new_n970), .C2(new_n949), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(G72));
  NAND3_X1  g790(.A1(new_n962), .A2(new_n969), .A3(new_n944), .ZN(new_n977));
  XNOR2_X1  g791(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n614), .A2(new_n429), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n978), .B(new_n979), .Z(new_n980));
  NAND2_X1  g794(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n658), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n342), .A2(new_n338), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n953), .A2(new_n944), .A3(new_n956), .A4(new_n954), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n985), .A2(new_n986), .A3(new_n980), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n985), .B2(new_n980), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n825), .A2(new_n831), .ZN(new_n990));
  INV_X1    g804(.A(new_n980), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n342), .A2(new_n288), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n328), .A2(new_n289), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n906), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n983), .A2(new_n989), .A3(new_n995), .ZN(G57));
endmodule


