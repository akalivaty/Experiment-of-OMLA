//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT64), .B(G238), .Z(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n226), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT67), .Z(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G68), .Z(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NOR2_X1   g0046(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT69), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(KEYINPUT69), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(new_n260), .B2(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  OAI211_X1 g0066(.A(G1), .B(G13), .C1(new_n253), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G274), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G41), .A2(G45), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT68), .B1(new_n274), .B2(G1), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n267), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n271), .B1(new_n277), .B2(G226), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n265), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G190), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT74), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n203), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n253), .A2(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n285), .B1(new_n286), .B2(new_n288), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n213), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n207), .A3(G1), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(new_n294), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n207), .A2(G1), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n202), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n300), .A2(new_n302), .B1(new_n202), .B2(new_n299), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n296), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n284), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n305), .B2(new_n304), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n279), .A2(G200), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n247), .B1(new_n283), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n281), .B(KEYINPUT74), .ZN(new_n311));
  INV_X1    g0111(.A(new_n247), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n308), .A4(new_n307), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n279), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n304), .C1(G179), .C2(new_n279), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n310), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n289), .A2(new_n301), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n300), .B1(new_n299), .B2(new_n289), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT7), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n254), .A2(new_n255), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(G20), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n249), .A2(new_n250), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G68), .ZN(new_n327));
  XNOR2_X1  g0127(.A(G58), .B(G68), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n294), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n325), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n251), .A2(new_n256), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n207), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n334), .B1(new_n336), .B2(new_n321), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n329), .B1(new_n337), .B2(new_n218), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n331), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n320), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G232), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G223), .A2(G1698), .ZN(new_n342));
  INV_X1    g0142(.A(G226), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(G1698), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n322), .B1(G33), .B2(G87), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n270), .B1(new_n276), .B2(new_n341), .C1(new_n267), .C2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n280), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(G200), .B2(new_n346), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n340), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT17), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n345), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n271), .B1(new_n354), .B2(new_n264), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n277), .A2(G232), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n314), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT81), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n346), .A2(G169), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(G179), .A3(new_n356), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT81), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT18), .B1(new_n363), .B2(new_n340), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n338), .A2(new_n331), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n319), .B1(new_n365), .B2(new_n332), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n358), .A4(new_n362), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n340), .A2(KEYINPUT17), .A3(new_n348), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n351), .A2(new_n364), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT71), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n291), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n289), .A2(new_n288), .B1(new_n207), .B2(new_n260), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n294), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n301), .A2(new_n260), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n300), .A2(new_n378), .B1(new_n260), .B2(new_n299), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G244), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n270), .B1(new_n276), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n384));
  INV_X1    g0184(.A(G107), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n384), .B1(new_n385), .B2(new_n257), .C1(new_n261), .C2(new_n217), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n264), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT72), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(G190), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n380), .B1(new_n387), .B2(G169), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n387), .A2(new_n352), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT73), .B(new_n380), .C1(new_n387), .C2(G169), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  OR3_X1    g0201(.A1(new_n317), .A2(new_n370), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n343), .A2(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n251), .A2(new_n256), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT76), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n251), .A2(new_n256), .A3(KEYINPUT76), .A4(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n251), .A2(new_n256), .A3(G232), .A4(G1698), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT77), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT77), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n264), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT13), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n271), .B1(new_n277), .B2(G238), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n416), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g0220(.A(G200), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT79), .B1(new_n299), .B2(new_n218), .ZN(new_n422));
  XOR2_X1   g0222(.A(new_n422), .B(KEYINPUT12), .Z(new_n423));
  INV_X1    g0223(.A(KEYINPUT11), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n290), .A2(G77), .B1(G20), .B2(new_n218), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n202), .B2(new_n288), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n294), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n423), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(KEYINPUT11), .A3(new_n294), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n300), .B(G68), .C1(G1), .C2(new_n207), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT77), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT77), .B1(new_n408), .B2(new_n411), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n434), .A2(new_n435), .A3(new_n267), .ZN(new_n436));
  INV_X1    g0236(.A(new_n418), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT13), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n433), .B1(new_n440), .B2(new_n280), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n438), .A2(KEYINPUT78), .A3(G190), .A4(new_n439), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n432), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(G179), .A3(new_n439), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT80), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n438), .A2(new_n439), .A3(new_n446), .A4(G179), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(G169), .B1(new_n419), .B2(new_n420), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT14), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n440), .A2(new_n451), .A3(G169), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n431), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n443), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n402), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  INV_X1    g0258(.A(G87), .ZN(new_n459));
  OR2_X1    g0259(.A1(KEYINPUT89), .A2(KEYINPUT22), .ZN(new_n460));
  NAND2_X1  g0260(.A1(KEYINPUT89), .A2(KEYINPUT22), .ZN(new_n461));
  AOI211_X1 g0261(.A(G20), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n257), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n322), .A2(new_n207), .A3(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT22), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n207), .B2(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n385), .A2(KEYINPUT23), .A3(G20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G116), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n468), .A2(new_n469), .B1(new_n471), .B2(new_n207), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n458), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n472), .ZN(new_n474));
  AOI211_X1 g0274(.A(KEYINPUT24), .B(new_n474), .C1(new_n463), .C2(new_n465), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n294), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n206), .A2(G33), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n300), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n385), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT25), .B1(new_n299), .B2(new_n385), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n478), .A2(new_n385), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n268), .A2(G1), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(G264), .A3(new_n267), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G250), .A2(G1698), .ZN(new_n488));
  INV_X1    g0288(.A(G257), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(G1698), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(new_n322), .B1(G33), .B2(G294), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n491), .B2(new_n267), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n267), .A2(G274), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(G190), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n487), .C1(new_n267), .C2(new_n491), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G200), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n476), .A2(new_n483), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n485), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n500), .A2(G250), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n267), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n494), .B2(new_n500), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n322), .A2(G244), .A3(G1698), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT85), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT85), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n322), .A2(new_n507), .A3(G244), .A4(G1698), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n324), .A2(G1698), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n471), .B1(new_n510), .B2(G238), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n352), .B(new_n504), .C1(new_n512), .C2(new_n267), .ZN(new_n513));
  INV_X1    g0313(.A(new_n299), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n372), .B2(new_n373), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n322), .A2(new_n207), .A3(G68), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n291), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n207), .B1(new_n410), .B2(new_n517), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n459), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT86), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT86), .B1(new_n520), .B2(new_n522), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n516), .B(new_n519), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n515), .B1(new_n527), .B2(new_n294), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n478), .B2(new_n374), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n509), .A2(new_n511), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n503), .B1(new_n530), .B2(new_n264), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n513), .B(new_n529), .C1(G169), .C2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G190), .B(new_n504), .C1(new_n512), .C2(new_n267), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n478), .A2(new_n459), .ZN(new_n534));
  AOI211_X1 g0334(.A(new_n515), .B(new_n534), .C1(new_n527), .C2(new_n294), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n533), .B(new_n535), .C1(new_n388), .C2(new_n531), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n499), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n337), .A2(new_n385), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n518), .A2(new_n385), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(new_n521), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n385), .A2(KEYINPUT6), .A3(G97), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n543), .A2(new_n207), .B1(new_n260), .B2(new_n288), .ZN(new_n544));
  OAI211_X1 g0344(.A(KEYINPUT82), .B(new_n294), .C1(new_n538), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n478), .A2(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n514), .A2(new_n518), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT83), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT82), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n336), .A2(new_n321), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n325), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n544), .B1(new_n553), .B2(G107), .ZN(new_n554));
  INV_X1    g0354(.A(new_n294), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n382), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n257), .A2(new_n258), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n322), .A2(G244), .A3(new_n258), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n558), .B1(G33), .B2(G283), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n264), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n486), .A2(new_n267), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n489), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n486), .A2(new_n494), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT84), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT84), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G200), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n564), .A2(new_n568), .A3(G190), .A4(new_n569), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n550), .A2(new_n556), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n556), .A2(new_n549), .A3(new_n545), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n314), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n564), .A2(new_n568), .A3(new_n352), .A4(new_n569), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n537), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n497), .A2(G179), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n314), .B2(new_n497), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n466), .A2(new_n472), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT24), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n466), .A2(new_n458), .A3(new_n472), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n555), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n580), .B1(new_n584), .B2(new_n482), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G283), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n587), .B(new_n207), .C1(G33), .C2(new_n518), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n294), .C1(new_n207), .C2(G116), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n589), .B(KEYINPUT20), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n514), .A2(G116), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G116), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n478), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT88), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n478), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n591), .B1(new_n596), .B2(G116), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT20), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n589), .B(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT88), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n322), .A2(G257), .A3(new_n258), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n322), .A2(KEYINPUT87), .A3(G257), .A4(new_n258), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(G264), .A2(G1698), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n335), .A2(G303), .B1(new_n322), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n267), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G270), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n495), .B1(new_n611), .B2(new_n565), .ZN(new_n612));
  OAI21_X1  g0412(.A(G169), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n586), .B1(new_n602), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n595), .A2(new_n601), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n610), .A2(new_n352), .A3(new_n612), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n610), .A2(new_n612), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n615), .A2(new_n619), .A3(KEYINPUT21), .A4(G169), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n585), .A2(new_n614), .A3(new_n617), .A4(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n615), .B1(G190), .B2(new_n618), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n388), .B2(new_n618), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n578), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n457), .A2(new_n625), .ZN(G372));
  OAI21_X1  g0426(.A(new_n366), .B1(new_n357), .B2(new_n353), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(new_n367), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n451), .B1(new_n440), .B2(G169), .ZN(new_n629));
  AOI211_X1 g0429(.A(KEYINPUT14), .B(new_n314), .C1(new_n438), .C2(new_n439), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n431), .B1(new_n631), .B2(new_n448), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n441), .A2(new_n442), .ZN(new_n633));
  INV_X1    g0433(.A(new_n432), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n400), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n351), .A2(new_n369), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n628), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT90), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n310), .A2(new_n313), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n642), .B(new_n628), .C1(new_n637), .C2(new_n638), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n316), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n621), .A2(new_n537), .A3(new_n573), .A4(new_n577), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n556), .A2(new_n549), .A3(new_n545), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n575), .A2(new_n576), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n532), .A2(new_n536), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT26), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n577), .A2(new_n653), .A3(new_n650), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n646), .B(new_n532), .C1(new_n652), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n457), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n645), .A2(new_n656), .ZN(G369));
  NAND3_X1  g0457(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n615), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n614), .A2(new_n617), .A3(new_n620), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n624), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n585), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n663), .B1(new_n584), .B2(new_n482), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n499), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n585), .A2(new_n663), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n663), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n676), .A2(new_n665), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT91), .ZN(new_n682));
  INV_X1    g0482(.A(new_n675), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n681), .B2(new_n683), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n679), .B1(new_n685), .B2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n210), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n206), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n521), .A2(new_n459), .A3(new_n593), .ZN(new_n692));
  INV_X1    g0492(.A(new_n689), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n691), .A2(new_n692), .B1(new_n216), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT94), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n655), .A2(new_n696), .A3(new_n680), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n655), .B2(new_n680), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT29), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n655), .A2(new_n680), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(KEYINPUT29), .B2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n618), .A2(new_n531), .A3(G179), .A4(new_n493), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT30), .B1(new_n702), .B2(new_n570), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n492), .B(new_n503), .C1(new_n530), .C2(new_n264), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n616), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT92), .ZN(new_n709));
  INV_X1    g0509(.A(new_n531), .ZN(new_n710));
  AOI21_X1  g0510(.A(G179), .B1(new_n493), .B2(new_n495), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n570), .A2(new_n619), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n709), .B1(new_n708), .B2(new_n712), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n713), .A2(new_n714), .A3(new_n680), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT93), .B1(new_n715), .B2(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n708), .A2(new_n712), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n680), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n625), .A2(new_n680), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(KEYINPUT92), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(new_n663), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n718), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n716), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n701), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n695), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n298), .A2(G20), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G45), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n690), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n670), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n668), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(G330), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n213), .B1(G20), .B2(new_n314), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n688), .A2(new_n335), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT96), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n746), .A2(G355), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n688), .A2(new_n322), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G45), .B2(new_n216), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n245), .A2(new_n268), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n749), .A2(new_n750), .B1(G116), .B2(new_n210), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n744), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n207), .A2(new_n352), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n754), .A2(new_n280), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n280), .A2(new_n388), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n207), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n755), .A2(G58), .B1(G87), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n280), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n207), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n760), .B(new_n257), .C1(new_n518), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G159), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT32), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n753), .A2(new_n756), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n388), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n753), .A2(new_n770), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n769), .A2(new_n202), .B1(new_n771), .B2(new_n218), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n753), .A2(new_n764), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n757), .A2(new_n770), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n773), .A2(new_n260), .B1(new_n774), .B2(new_n385), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n763), .A2(new_n768), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n755), .A2(G322), .B1(G329), .B2(new_n766), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n778), .B2(new_n774), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n758), .B1(new_n773), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT97), .B(G326), .Z(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  OAI22_X1  g0584(.A1(new_n783), .A2(new_n769), .B1(new_n784), .B2(new_n771), .ZN(new_n785));
  INV_X1    g0585(.A(G294), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n335), .B1(new_n786), .B2(new_n762), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n779), .A2(new_n782), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n743), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n752), .A2(new_n789), .A3(new_n734), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n737), .B1(new_n742), .B2(new_n790), .ZN(G396));
  INV_X1    g0591(.A(new_n727), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n400), .A2(KEYINPUT98), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n381), .A2(new_n680), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n400), .A2(KEYINPUT98), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n793), .A2(new_n394), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n636), .A2(new_n794), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(new_n700), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n792), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n734), .B1(new_n792), .B2(new_n801), .ZN(new_n804));
  INV_X1    g0604(.A(new_n799), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n738), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n743), .A2(new_n738), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n734), .B1(G77), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n771), .ZN(new_n810));
  INV_X1    g0610(.A(new_n773), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G150), .A2(new_n810), .B1(new_n811), .B2(G159), .ZN(new_n812));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  INV_X1    g0614(.A(new_n755), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n812), .B1(new_n813), .B2(new_n769), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n758), .A2(new_n202), .B1(new_n765), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G58), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n762), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n774), .A2(new_n218), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n821), .A2(new_n823), .A3(new_n324), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n818), .A2(new_n819), .A3(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n758), .A2(new_n385), .B1(new_n765), .B2(new_n781), .ZN(new_n827));
  INV_X1    g0627(.A(new_n769), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(G303), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n762), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n257), .B1(G97), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n774), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n755), .A2(G294), .B1(G87), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G116), .A2(new_n811), .B1(new_n810), .B2(G283), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n829), .A2(new_n831), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n826), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n809), .B1(new_n836), .B2(new_n743), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n803), .A2(new_n804), .B1(new_n806), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  OAI21_X1  g0639(.A(G77), .B1(new_n822), .B2(new_n218), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n840), .A2(new_n216), .B1(G50), .B2(new_n218), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(G1), .A3(new_n298), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT100), .ZN(new_n843));
  INV_X1    g0643(.A(new_n543), .ZN(new_n844));
  OAI211_X1 g0644(.A(G116), .B(new_n214), .C1(new_n844), .C2(KEYINPUT35), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n845), .A2(KEYINPUT99), .B1(KEYINPUT35), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(KEYINPUT99), .B2(new_n845), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT36), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n445), .A2(new_n447), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n450), .A2(new_n452), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n454), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n431), .A2(new_n680), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n635), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT101), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n455), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n854), .B1(new_n453), .B2(new_n443), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT102), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n862), .B(new_n854), .C1(new_n453), .C2(new_n443), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n858), .A2(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n723), .A2(new_n718), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n625), .A2(new_n680), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n721), .A2(new_n722), .A3(new_n719), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT105), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n721), .A2(new_n722), .A3(KEYINPUT105), .A4(new_n719), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n799), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT106), .B1(new_n864), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT101), .B1(new_n455), .B2(new_n855), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n632), .A2(new_n857), .A3(new_n443), .A4(new_n854), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n635), .A2(new_n448), .A3(new_n631), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n862), .B1(new_n877), .B2(new_n854), .ZN(new_n878));
  INV_X1    g0678(.A(new_n863), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n875), .A2(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n873), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT106), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n366), .A2(new_n358), .A3(new_n362), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n661), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n366), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n349), .B(new_n891), .C1(new_n885), .C2(new_n886), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n627), .A2(new_n891), .A3(new_n349), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(KEYINPUT37), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n638), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n891), .B1(new_n628), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n884), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT16), .B1(new_n327), .B2(new_n329), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n319), .B1(new_n332), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n359), .A2(new_n360), .A3(new_n661), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n340), .A2(new_n348), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n889), .A2(new_n892), .B1(new_n888), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n900), .A2(new_n890), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n370), .A2(KEYINPUT103), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT103), .B1(new_n370), .B2(new_n904), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n903), .B(KEYINPUT38), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT40), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n874), .A2(new_n883), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT107), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT107), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n874), .A2(new_n883), .A3(new_n913), .A4(new_n910), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n370), .A2(new_n904), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n370), .A2(KEYINPUT103), .A3(new_n904), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n920), .B2(new_n903), .ZN(new_n921));
  INV_X1    g0721(.A(new_n907), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n864), .A2(new_n923), .A3(new_n873), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n912), .A2(new_n914), .B1(new_n915), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n867), .ZN(new_n927));
  INV_X1    g0727(.A(new_n872), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n457), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n926), .A2(new_n930), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n931), .A2(new_n932), .A3(new_n669), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT108), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n628), .A2(new_n890), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n908), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n920), .A2(new_n903), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n884), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(KEYINPUT39), .A3(new_n907), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n853), .A2(new_n663), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n936), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n793), .A2(new_n796), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n663), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n655), .A2(new_n680), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n947), .B2(new_n799), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n864), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n922), .B2(new_n921), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n701), .A2(new_n457), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n645), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n935), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n954), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n934), .A2(new_n956), .B1(new_n206), .B2(new_n731), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n850), .B1(new_n955), .B2(new_n957), .ZN(G367));
  OAI211_X1 g0758(.A(new_n573), .B(new_n577), .C1(new_n647), .C2(new_n680), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n649), .A2(new_n663), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n678), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n535), .A2(new_n680), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n651), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n532), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n962), .B(new_n966), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n968));
  INV_X1    g0768(.A(new_n961), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT42), .B1(new_n681), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n577), .B1(new_n959), .B2(new_n585), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n680), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n681), .A2(KEYINPUT42), .A3(new_n969), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n968), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT109), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n967), .B(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT110), .ZN(new_n978));
  INV_X1    g0778(.A(new_n686), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n684), .A3(new_n969), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n961), .B1(new_n685), .B2(new_n686), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(KEYINPUT45), .B(new_n961), .C1(new_n685), .C2(new_n686), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n982), .A2(new_n679), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n679), .B1(new_n982), .B2(new_n987), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n681), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n676), .B1(new_n665), .B2(new_n680), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n671), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n728), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n728), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n689), .B(KEYINPUT41), .Z(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n978), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n988), .A2(new_n989), .A3(new_n995), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n728), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n978), .B(new_n998), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n732), .A2(G1), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n977), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n233), .A2(new_n748), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n744), .B1(new_n374), .B2(new_n210), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n734), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G77), .A2(new_n832), .B1(new_n766), .B2(G137), .ZN(new_n1010));
  INV_X1    g0810(.A(G159), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n822), .B2(new_n758), .C1(new_n1011), .C2(new_n771), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n755), .A2(G150), .B1(G50), .B2(new_n811), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n814), .B2(new_n769), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n762), .A2(new_n218), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1012), .A2(new_n1014), .A3(new_n335), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G294), .A2(new_n810), .B1(new_n766), .B2(G317), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n781), .B2(new_n769), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n815), .A2(new_n780), .B1(new_n518), .B2(new_n774), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n759), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT46), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n758), .B2(new_n593), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(new_n385), .C2(new_n762), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n324), .B1(new_n773), .B2(new_n778), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1018), .A2(new_n1019), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1016), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT47), .Z(new_n1027));
  AOI21_X1  g0827(.A(new_n1009), .B1(new_n1027), .B2(new_n743), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n741), .B2(new_n965), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1006), .A2(new_n1029), .ZN(G387));
  AOI22_X1  g0830(.A1(new_n746), .A2(new_n692), .B1(new_n385), .B2(new_n688), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n289), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  AOI211_X1 g0833(.A(G45), .B(new_n692), .C1(G68), .C2(G77), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n748), .B(new_n1035), .C1(new_n238), .C2(new_n268), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT111), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n744), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1037), .A2(KEYINPUT111), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n734), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n322), .B1(new_n832), .B2(G116), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n762), .A2(new_n778), .B1(new_n758), .B2(new_n786), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n755), .A2(G317), .B1(new_n828), .B2(G322), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n780), .B2(new_n773), .C1(new_n781), .C2(new_n771), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1043), .B1(new_n765), .B2(new_n783), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n769), .A2(new_n1011), .B1(new_n765), .B2(new_n286), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n324), .B(new_n1053), .C1(G97), .C2(new_n832), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n372), .A2(new_n830), .A3(new_n373), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n758), .A2(new_n260), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G68), .B2(new_n811), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n289), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n755), .A2(G50), .B1(new_n1058), .B2(new_n810), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT113), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n743), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1042), .B(new_n1064), .C1(new_n677), .C2(new_n740), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n994), .B2(new_n1003), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n995), .A2(new_n689), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n728), .A2(new_n994), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(G393));
  NOR2_X1   g0869(.A1(new_n1000), .A2(new_n693), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n990), .A2(new_n995), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n748), .A2(new_n242), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1073), .B(new_n744), .C1(new_n518), .C2(new_n210), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT114), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT114), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n734), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G303), .A2(new_n810), .B1(new_n832), .B2(G107), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n830), .A2(G116), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1078), .A2(new_n335), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G294), .A2(new_n811), .B1(new_n766), .B2(G322), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n778), .C2(new_n758), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n755), .A2(G311), .B1(new_n828), .B2(G317), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n755), .A2(G159), .B1(new_n828), .B2(G150), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G50), .A2(new_n810), .B1(new_n759), .B2(G68), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1058), .A2(new_n811), .B1(new_n766), .B2(G143), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n830), .A2(G77), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n324), .B1(new_n832), .B2(G87), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1082), .A2(new_n1084), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1077), .B1(new_n743), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n961), .B2(new_n741), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n990), .B2(new_n1004), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1072), .A2(new_n1095), .ZN(G390));
  INV_X1    g0896(.A(KEYINPUT115), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n943), .B(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n697), .A2(new_n698), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n946), .B1(new_n1099), .B2(new_n799), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n908), .B(new_n1098), .C1(new_n1100), .C2(new_n864), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n948), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n943), .B1(new_n880), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n942), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n873), .A2(new_n669), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n880), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n726), .A2(G330), .A3(new_n799), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT116), .B1(new_n864), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n726), .A2(G330), .A3(new_n799), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n880), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1114), .B(new_n1101), .C1(new_n942), .C2(new_n1103), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n457), .A2(new_n929), .A3(G330), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n644), .A2(new_n952), .A3(new_n316), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1100), .B1(new_n1105), .B2(new_n880), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1113), .B2(new_n1110), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n864), .A2(new_n1109), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n948), .B1(new_n1106), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1119), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT117), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n697), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n698), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n799), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n946), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n881), .A2(G330), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n864), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1114), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1106), .A2(new_n1122), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1102), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1118), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT117), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n1115), .A4(new_n1108), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n693), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT118), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1116), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1108), .A2(new_n1115), .A3(KEYINPUT118), .ZN(new_n1142));
  AND4_X1   g0942(.A1(KEYINPUT119), .A2(new_n1141), .A3(new_n1142), .A4(new_n1124), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1136), .B1(new_n1116), .B2(new_n1140), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT119), .B1(new_n1144), .B2(new_n1142), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1139), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n734), .B1(new_n1058), .B2(new_n808), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n815), .A2(new_n593), .B1(new_n769), .B2(new_n778), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G107), .B2(new_n810), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n773), .A2(new_n518), .B1(new_n765), .B2(new_n786), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n824), .B(new_n1150), .C1(G87), .C2(new_n759), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1149), .A2(new_n335), .A3(new_n1089), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n815), .A2(new_n820), .B1(new_n765), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G137), .B2(new_n810), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT53), .B1(new_n758), .B2(new_n286), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G128), .A2(new_n828), .B1(new_n811), .B2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n758), .A2(KEYINPUT53), .A3(new_n286), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G159), .B2(new_n830), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1155), .A2(new_n1156), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n257), .B1(new_n202), .B2(new_n774), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT120), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1152), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1147), .B1(new_n1165), .B2(new_n743), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n942), .B2(new_n739), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1116), .B2(new_n1004), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1146), .A2(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(new_n951), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n304), .A2(new_n890), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n317), .B(new_n1172), .Z(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n912), .A2(new_n914), .ZN(new_n1176));
  OAI21_X1  g0976(.A(G330), .B1(new_n924), .B2(KEYINPUT40), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1175), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1175), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1180), .B(new_n1177), .C1(new_n912), .C2(new_n914), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1171), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n858), .A2(new_n859), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n861), .A2(new_n863), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n873), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n909), .B1(new_n1185), .B2(new_n882), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n913), .B1(new_n1186), .B2(new_n874), .ZN(new_n1187));
  AND4_X1   g0987(.A1(new_n913), .A2(new_n874), .A3(new_n883), .A4(new_n910), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1178), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1180), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1176), .A2(new_n1178), .A3(new_n1175), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n951), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1182), .A2(new_n1192), .A3(KEYINPUT121), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1119), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT121), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1190), .A2(new_n1196), .A3(new_n951), .A4(new_n1191), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1194), .B2(new_n1119), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1182), .A2(new_n1192), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n693), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1193), .A2(new_n1003), .A3(new_n1197), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n820), .A2(new_n771), .B1(new_n758), .B2(new_n1157), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n755), .A2(G128), .B1(new_n828), .B2(G125), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n813), .B2(new_n773), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1206), .B(new_n1208), .C1(G150), .C2(new_n830), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n253), .B(new_n266), .C1(new_n774), .C2(new_n1011), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G124), .B2(new_n766), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n774), .A2(new_n822), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G116), .B2(new_n828), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n518), .B2(new_n771), .C1(new_n374), .C2(new_n773), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n324), .A2(new_n266), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1056), .A2(new_n1219), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n815), .A2(new_n385), .B1(new_n765), .B2(new_n778), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1218), .A2(new_n1015), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1219), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1215), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n743), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n733), .B1(new_n202), .B2(new_n807), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n1180), .C2(new_n739), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1205), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1204), .A2(new_n1231), .ZN(G375));
  NOR2_X1   g1032(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1233));
  OR3_X1    g1033(.A1(new_n1233), .A2(KEYINPUT122), .A3(new_n1004), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n733), .B1(new_n218), .B2(new_n807), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n755), .A2(G137), .B1(new_n810), .B2(new_n1158), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n820), .B2(new_n769), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT123), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(KEYINPUT123), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n286), .A2(new_n773), .B1(new_n758), .B2(new_n1011), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G128), .B2(new_n766), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n324), .B(new_n1216), .C1(G50), .C2(new_n830), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n769), .A2(new_n786), .B1(new_n774), .B2(new_n260), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n771), .A2(new_n593), .B1(new_n765), .B2(new_n780), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n257), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n518), .A2(new_n758), .B1(new_n773), .B2(new_n385), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G283), .B2(new_n755), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1248), .A3(new_n1055), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1243), .A2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(KEYINPUT124), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n743), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1235), .B1(new_n1251), .B2(new_n1253), .C1(new_n880), .C2(new_n739), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT122), .B1(new_n1233), .B2(new_n1004), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1234), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1233), .A2(new_n1118), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n998), .A3(new_n1124), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(G381));
  NOR2_X1   g1060(.A1(G375), .A2(G378), .ZN(new_n1261));
  OR2_X1    g1061(.A1(G390), .A2(G384), .ZN(new_n1262));
  OR2_X1    g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(new_n1262), .A2(G387), .A3(G381), .A4(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(G407));
  OAI21_X1  g1065(.A(new_n1261), .B1(new_n1264), .B2(new_n662), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(G213), .ZN(G409));
  AND3_X1   g1067(.A1(G390), .A2(new_n1006), .A3(new_n1029), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G390), .B1(new_n1006), .B2(new_n1029), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT126), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  XOR2_X1   g1070(.A(G393), .B(G396), .Z(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1271), .ZN(new_n1273));
  OAI211_X1 g1073(.A(KEYINPUT126), .B(new_n1273), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1258), .B1(new_n1276), .B2(new_n1136), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1233), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n689), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n838), .B1(new_n1280), .B2(new_n1256), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1257), .A2(new_n1279), .A3(G384), .ZN(new_n1282));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G343), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT125), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1282), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(G2897), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1286), .B(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1193), .A2(new_n1195), .A3(new_n998), .A4(new_n1197), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1229), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1202), .B2(new_n1003), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G378), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1230), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(G378), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1288), .B1(new_n1294), .B2(new_n1284), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1204), .A2(G378), .A3(new_n1231), .ZN(new_n1298));
  INV_X1    g1098(.A(G378), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1284), .B(new_n1297), .C1(new_n1298), .C2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1295), .B(new_n1296), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1297), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1284), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1298), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1305), .B(new_n1306), .C1(new_n1307), .C2(new_n1292), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1275), .B1(new_n1304), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1275), .B1(new_n1308), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1302), .A2(KEYINPUT63), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1312), .A2(new_n1296), .A3(new_n1313), .A4(new_n1295), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(new_n1314), .ZN(G405));
  OAI21_X1  g1115(.A(new_n1297), .B1(new_n1293), .B2(G378), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(G375), .A2(new_n1299), .A3(new_n1305), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1275), .A2(new_n1317), .A3(new_n1316), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1307), .A2(KEYINPUT127), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1307), .A2(KEYINPUT127), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(new_n1320), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(G402));
endmodule


