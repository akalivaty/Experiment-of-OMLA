//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT65), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n208), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n213), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  INV_X1    g0042(.A(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT66), .B(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G107), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G97), .ZN(new_n248));
  INV_X1    g0048(.A(G97), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G107), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n246), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G274), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n255), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n256), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(KEYINPUT67), .A3(new_n261), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n263), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G97), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n234), .A2(G1698), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G226), .B2(G1698), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n272), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n261), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n278), .A2(new_n279), .B1(new_n280), .B2(G238), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n269), .A2(new_n271), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT13), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT13), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n269), .A2(new_n284), .A3(new_n271), .A4(new_n281), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT71), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n282), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n290), .A2(G179), .A3(new_n291), .A4(new_n285), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT14), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n286), .A2(new_n293), .A3(G169), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G68), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT12), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n296), .A2(new_n227), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n207), .A2(G20), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(G68), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n227), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G20), .A2(G33), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n310), .A2(new_n202), .B1(new_n208), .B2(G68), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n208), .A2(G33), .ZN(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT11), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT72), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n300), .A2(new_n317), .A3(new_n305), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n307), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n295), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n286), .B2(G200), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n290), .A2(G190), .A3(new_n291), .A4(new_n285), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  XOR2_X1   g0125(.A(KEYINPUT8), .B(G58), .Z(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n304), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n327), .A2(new_n302), .B1(new_n296), .B2(new_n326), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT76), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT76), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n330), .B1(new_n296), .B2(new_n326), .C1(new_n327), .C2(new_n302), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n308), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT7), .B1(new_n277), .B2(new_n208), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  INV_X1    g0135(.A(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(G68), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT75), .ZN(new_n342));
  INV_X1    g0142(.A(G159), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n310), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n309), .A2(KEYINPUT75), .A3(G159), .ZN(new_n345));
  XNOR2_X1  g0145(.A(G58), .B(G68), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n344), .A2(new_n345), .B1(new_n346), .B2(G20), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n333), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT74), .B1(new_n275), .B2(new_n276), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT74), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n337), .A2(new_n352), .A3(new_n338), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n353), .A3(new_n208), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n340), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT16), .B(new_n347), .C1(new_n356), .C2(new_n298), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n332), .B1(new_n350), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n215), .A2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G223), .B2(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G87), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n361), .A2(new_n277), .B1(new_n336), .B2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n279), .B1(G232), .B2(new_n280), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n359), .B1(new_n364), .B2(new_n268), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n280), .A2(G232), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n215), .B2(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n337), .A2(new_n338), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(new_n369), .B1(G33), .B2(G87), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n366), .B1(new_n370), .B2(new_n257), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n266), .A2(KEYINPUT67), .A3(new_n261), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT67), .B1(new_n266), .B2(new_n261), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n365), .B1(G179), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT18), .B1(new_n358), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n344), .A2(new_n345), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n346), .A2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n337), .A2(new_n208), .A3(new_n338), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n355), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n298), .B1(new_n382), .B2(new_n339), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n349), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n357), .A2(new_n308), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n332), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n375), .A2(G179), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n375), .B2(new_n359), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G200), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n371), .B2(new_n374), .ZN(new_n393));
  INV_X1    g0193(.A(G190), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n364), .A2(new_n394), .A3(new_n268), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT77), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(KEYINPUT77), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n358), .A2(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AND4_X1   g0201(.A1(new_n385), .A2(new_n396), .A3(new_n386), .A4(new_n400), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n377), .B(new_n391), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n303), .A2(G77), .A3(new_n304), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT68), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n297), .A2(new_n313), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n326), .A2(new_n309), .B1(G20), .B2(G77), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT15), .B(G87), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n312), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n308), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G1698), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n277), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(G238), .B1(new_n277), .B2(G107), .ZN(new_n416));
  AOI21_X1  g0216(.A(G1698), .B1(new_n337), .B2(new_n338), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G232), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n257), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n280), .A2(G244), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n268), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(G200), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  OR3_X1    g0222(.A1(new_n419), .A2(new_n421), .A3(new_n394), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n413), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OR3_X1    g0224(.A1(new_n419), .A2(new_n421), .A3(G179), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n359), .B1(new_n419), .B2(new_n421), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n412), .A3(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n374), .B1(G226), .B2(new_n280), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n415), .A2(G223), .B1(new_n277), .B2(G77), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n417), .A2(G222), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n279), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n392), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT10), .B1(new_n434), .B2(KEYINPUT69), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(new_n433), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G200), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n429), .A2(new_n433), .A3(G190), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n303), .A2(G50), .A3(new_n304), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(G50), .B2(new_n296), .ZN(new_n441));
  INV_X1    g0241(.A(new_n312), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n326), .A2(new_n442), .B1(G150), .B2(new_n309), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n203), .A2(G20), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n333), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT9), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT9), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n441), .B2(new_n445), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n438), .A2(new_n439), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n436), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n447), .A2(new_n449), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n435), .A2(new_n452), .A3(new_n438), .A4(new_n439), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n446), .B1(new_n437), .B2(new_n359), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(G179), .B2(new_n437), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n325), .A2(new_n404), .A3(new_n428), .A4(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n302), .B1(new_n207), .B2(G33), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT25), .B1(new_n297), .B2(new_n247), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n247), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n462), .A2(G107), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT86), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n208), .B2(G107), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT23), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n468), .B(new_n471), .C1(new_n208), .C2(G107), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n470), .A2(new_n472), .B1(G116), .B2(new_n442), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n208), .B1(new_n275), .B2(new_n276), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT85), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT22), .ZN(new_n477));
  OAI21_X1  g0277(.A(G87), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n474), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n362), .B1(KEYINPUT85), .B2(KEYINPUT22), .ZN(new_n480));
  INV_X1    g0280(.A(new_n474), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n369), .A2(new_n480), .A3(new_n208), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT24), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n473), .A2(new_n479), .A3(new_n485), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n467), .B1(new_n487), .B2(new_n308), .ZN(new_n488));
  AOI211_X1 g0288(.A(KEYINPUT87), .B(new_n333), .C1(new_n484), .C2(new_n486), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n466), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n207), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n493));
  OAI211_X1 g0293(.A(G264), .B(new_n257), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n260), .A2(G1), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT80), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(KEYINPUT5), .C2(new_n259), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(KEYINPUT80), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(new_n498), .A3(new_n266), .A4(new_n491), .ZN(new_n499));
  OAI211_X1 g0299(.A(G257), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G294), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n417), .A2(KEYINPUT88), .A3(G250), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(new_n414), .C1(new_n275), .C2(new_n276), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT88), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n502), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n494), .B(new_n499), .C1(new_n507), .C2(new_n257), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G169), .ZN(new_n509));
  INV_X1    g0309(.A(G179), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n508), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n490), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT89), .ZN(new_n513));
  INV_X1    g0313(.A(new_n502), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT88), .B1(new_n417), .B2(G250), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n504), .A2(new_n505), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n279), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(new_n394), .A3(new_n494), .A4(new_n499), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n508), .A2(new_n392), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n466), .C1(new_n489), .C2(new_n488), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n512), .A2(new_n513), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n513), .B1(new_n512), .B2(new_n522), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n277), .A2(G303), .ZN(new_n526));
  OAI211_X1 g0326(.A(G264), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n527));
  OAI211_X1 g0327(.A(G257), .B(new_n414), .C1(new_n275), .C2(new_n276), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n526), .A2(KEYINPUT84), .A3(new_n527), .A4(new_n528), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n257), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n257), .B1(new_n492), .B2(new_n493), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n499), .B1(new_n217), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n208), .C1(G33), .C2(new_n249), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n538), .B(new_n308), .C1(new_n208), .C2(G116), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n539), .B(KEYINPUT20), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n296), .A2(G116), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n303), .B1(G1), .B2(new_n336), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n216), .ZN(new_n544));
  OAI21_X1  g0344(.A(G169), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT21), .B1(new_n536), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT20), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n539), .B(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n541), .B1(new_n462), .B2(G116), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n359), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n551), .C1(new_n535), .C2(new_n533), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n540), .A2(new_n544), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n499), .B(G179), .C1(new_n217), .C2(new_n534), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n531), .A2(new_n532), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n279), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n546), .A2(new_n552), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n536), .A2(G190), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n559), .B(new_n553), .C1(new_n392), .C2(new_n536), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR4_X1   g0361(.A1(new_n313), .A2(KEYINPUT78), .A3(G20), .A4(G33), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT78), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n309), .B2(G77), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n247), .A2(KEYINPUT6), .A3(G97), .ZN(new_n566));
  XNOR2_X1  g0366(.A(G97), .B(G107), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT6), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n565), .B1(new_n569), .B2(new_n208), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n247), .B1(new_n382), .B2(new_n339), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n308), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n296), .A2(G97), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n462), .B2(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G257), .B(new_n257), .C1(new_n492), .C2(new_n493), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n499), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(new_n414), .C1(new_n275), .C2(new_n276), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT79), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n579), .B2(new_n580), .ZN(new_n583));
  OAI211_X1 g0383(.A(G250), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n537), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n578), .B1(new_n586), .B2(new_n257), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n575), .B1(G200), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n579), .A2(new_n580), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT4), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n591));
  INV_X1    g0391(.A(new_n585), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n577), .B1(new_n593), .B2(new_n279), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G190), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n588), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n510), .B(new_n578), .C1(new_n586), .C2(new_n257), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n575), .C1(G169), .C2(new_n594), .ZN(new_n598));
  INV_X1    g0398(.A(new_n409), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n296), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n208), .B1(new_n272), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  AND2_X1   g0403(.A1(KEYINPUT82), .A2(G87), .ZN(new_n604));
  NOR2_X1   g0404(.A1(KEYINPUT82), .A2(G87), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(G97), .A2(G107), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OR2_X1    g0408(.A1(KEYINPUT82), .A2(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(KEYINPUT82), .A2(G87), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n603), .A2(new_n609), .A3(new_n607), .A4(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n602), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n601), .B1(new_n312), .B2(new_n249), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n475), .B2(new_n298), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n600), .B1(new_n616), .B2(new_n308), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n462), .A2(G87), .ZN(new_n618));
  OAI211_X1 g0418(.A(G238), .B(new_n414), .C1(new_n275), .C2(new_n276), .ZN(new_n619));
  OAI211_X1 g0419(.A(G244), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n620));
  NAND2_X1  g0420(.A1(G33), .A2(G116), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n279), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n495), .A2(new_n264), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n257), .C1(G250), .C2(new_n495), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(G190), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G200), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n617), .A2(new_n618), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n600), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n462), .A2(new_n599), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n609), .A2(new_n607), .A3(new_n610), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT83), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n606), .A2(new_n603), .A3(new_n607), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n614), .B1(new_n635), .B2(new_n602), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n630), .B(new_n631), .C1(new_n636), .C2(new_n333), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n623), .A2(new_n510), .A3(new_n625), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT81), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n627), .A2(new_n359), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n623), .A2(KEYINPUT81), .A3(new_n510), .A4(new_n625), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n637), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n596), .A2(new_n598), .A3(new_n629), .A4(new_n643), .ZN(new_n644));
  NOR4_X1   g0444(.A1(new_n461), .A2(new_n525), .A3(new_n561), .A4(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n323), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n320), .B1(new_n646), .B2(new_n427), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n401), .A2(new_n402), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n391), .A2(new_n377), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n454), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n456), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n596), .A2(new_n598), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n637), .A2(new_n641), .A3(new_n638), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n629), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n522), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT90), .B1(new_n512), .B2(new_n558), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n512), .A2(KEYINPUT90), .A3(new_n558), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n643), .A2(new_n629), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT26), .B1(new_n661), .B2(new_n598), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n575), .B1(new_n594), .B2(G169), .ZN(new_n663));
  INV_X1    g0463(.A(new_n597), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n629), .A4(new_n655), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n662), .A2(new_n667), .A3(new_n655), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT91), .ZN(new_n669));
  INV_X1    g0469(.A(new_n655), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n587), .A2(new_n359), .B1(new_n572), .B2(new_n574), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n643), .A3(new_n629), .A4(new_n597), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n670), .B1(new_n672), .B2(KEYINPUT26), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT91), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n667), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n659), .A2(new_n660), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n653), .B1(new_n461), .B2(new_n676), .ZN(G369));
  INV_X1    g0477(.A(new_n466), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n487), .A2(new_n308), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT87), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n487), .A2(new_n467), .A3(new_n308), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G213), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n523), .B2(new_n524), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n490), .A2(new_n511), .A3(new_n688), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n688), .B1(new_n540), .B2(new_n544), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n558), .A2(new_n560), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n558), .B2(new_n697), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT93), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n512), .A2(new_n688), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n558), .A2(new_n688), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n696), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n211), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n635), .A2(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n225), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT95), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n669), .A2(new_n675), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n512), .A2(new_n558), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT90), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND4_X1   g0520(.A1(new_n522), .A2(new_n656), .A3(new_n598), .A4(new_n596), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n660), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n688), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n716), .B1(new_n723), .B2(KEYINPUT29), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  OAI211_X1 g0525(.A(KEYINPUT95), .B(new_n725), .C1(new_n676), .C2(new_n688), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT96), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n718), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n656), .A2(new_n665), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT26), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n672), .A2(KEYINPUT26), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(new_n655), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n688), .A2(new_n725), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n724), .A2(new_n726), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n561), .A2(new_n644), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n738), .B(new_n689), .C1(new_n523), .C2(new_n524), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n627), .A2(new_n554), .ZN(new_n740));
  INV_X1    g0540(.A(new_n494), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n517), .B2(new_n279), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n740), .A2(new_n594), .A3(new_n557), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT94), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT30), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(KEYINPUT94), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n583), .A2(new_n585), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n257), .B1(new_n748), .B2(new_n591), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n749), .A2(new_n577), .B1(new_n533), .B2(new_n535), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n508), .A2(new_n510), .A3(new_n627), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n745), .A2(new_n747), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n688), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n739), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n737), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n715), .B1(new_n762), .B2(G1), .ZN(G364));
  AND2_X1   g0563(.A1(new_n208), .A2(G13), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n207), .B1(new_n764), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n710), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT97), .Z(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n227), .B1(G20), .B2(new_n359), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n246), .A2(G45), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n351), .A2(new_n353), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n709), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n774), .B(new_n776), .C1(G45), .C2(new_n226), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n709), .A2(new_n277), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G355), .B1(new_n216), .B2(new_n709), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n772), .B(new_n773), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n208), .A2(new_n394), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n510), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n208), .A2(G190), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G179), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G322), .A2(new_n784), .B1(new_n788), .B2(G329), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n392), .A2(G179), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n781), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G303), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n782), .A2(new_n785), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n277), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G190), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n208), .B1(new_n786), .B2(G190), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n798), .A2(new_n394), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(G294), .B1(G326), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n785), .A2(new_n790), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT99), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G283), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n794), .A2(new_n801), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(G107), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n788), .A2(G159), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT32), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n791), .A2(new_n606), .ZN(new_n813));
  AND4_X1   g0613(.A1(new_n369), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n802), .A2(new_n249), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n811), .B2(KEYINPUT32), .ZN(new_n816));
  INV_X1    g0616(.A(new_n799), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n814), .B(new_n816), .C1(new_n298), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n795), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G58), .A2(new_n784), .B1(new_n819), .B2(G77), .ZN(new_n820));
  INV_X1    g0620(.A(new_n804), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n202), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT98), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n809), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n769), .B(new_n780), .C1(new_n773), .C2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT100), .Z(new_n826));
  INV_X1    g0626(.A(new_n772), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n699), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n700), .A2(new_n767), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(G330), .B2(new_n699), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n412), .A2(new_n688), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n424), .A2(new_n427), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(KEYINPUT101), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT101), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n424), .A2(new_n427), .A3(new_n836), .A4(new_n833), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n689), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n673), .A2(new_n674), .A3(new_n667), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n674), .B1(new_n673), .B2(new_n667), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n660), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n844), .A2(new_n657), .A3(new_n658), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n840), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n427), .A2(new_n689), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n835), .A2(new_n837), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n846), .B1(new_n723), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n767), .B1(new_n849), .B2(new_n760), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n760), .B2(new_n849), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n773), .A2(new_n770), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n768), .B1(G77), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n369), .B(new_n815), .C1(G116), .C2(new_n819), .ZN(new_n854));
  INV_X1    g0654(.A(G294), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n247), .A2(new_n791), .B1(new_n783), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G311), .B2(new_n788), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G283), .A2(new_n799), .B1(new_n804), .B2(G303), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n807), .A2(G87), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n854), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G143), .A2(new_n784), .B1(new_n819), .B2(G159), .ZN(new_n861));
  INV_X1    g0661(.A(G137), .ZN(new_n862));
  INV_X1    g0662(.A(G150), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n861), .B1(new_n821), .B2(new_n862), .C1(new_n863), .C2(new_n817), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT34), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n807), .A2(G68), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n791), .A2(new_n202), .B1(new_n787), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n775), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n869), .B(new_n870), .C1(G58), .C2(new_n803), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n866), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n864), .A2(new_n865), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n860), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n853), .B1(new_n874), .B2(new_n773), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n848), .B2(new_n771), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n851), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(G384));
  INV_X1    g0678(.A(new_n569), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n216), .B(new_n229), .C1(new_n879), .C2(KEYINPUT35), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(KEYINPUT35), .B2(new_n879), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT36), .Z(new_n882));
  INV_X1    g0682(.A(new_n225), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n883), .B(G77), .C1(new_n243), .C2(new_n298), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n202), .A2(G68), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n207), .B(G13), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n888));
  INV_X1    g0688(.A(new_n686), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n403), .A2(new_n387), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n376), .A2(new_n686), .B1(new_n385), .B2(new_n386), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT106), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n387), .B1(new_n389), .B2(new_n889), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n358), .A2(new_n396), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n895), .A2(new_n893), .A3(new_n896), .A4(new_n891), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n888), .B1(new_n890), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT107), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n347), .B1(new_n356), .B2(new_n298), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(new_n349), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n357), .A2(new_n308), .ZN(new_n907));
  OAI211_X1 g0707(.A(KEYINPUT103), .B(new_n386), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n349), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n308), .A3(new_n357), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT103), .B1(new_n911), .B2(new_n386), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n403), .A2(new_n889), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n386), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n376), .A2(new_n686), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n919), .A3(new_n908), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n915), .B1(new_n920), .B2(new_n896), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n897), .A2(new_n891), .ZN(new_n922));
  OAI211_X1 g0722(.A(KEYINPUT38), .B(new_n914), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT107), .B(new_n888), .C1(new_n890), .C2(new_n900), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n903), .A2(new_n904), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n922), .ZN(new_n926));
  INV_X1    g0726(.A(new_n896), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n913), .B2(new_n919), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n928), .B2(new_n915), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n929), .B2(new_n914), .ZN(new_n930));
  INV_X1    g0730(.A(new_n923), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT39), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n925), .A2(new_n932), .A3(KEYINPUT108), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n320), .A2(new_n688), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n924), .A2(new_n923), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT108), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n904), .A4(new_n903), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n319), .A2(new_n688), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n320), .A2(new_n323), .A3(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n319), .B(new_n688), .C1(new_n646), .C2(new_n295), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT102), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n839), .B1(new_n717), .B2(new_n722), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n427), .A2(new_n688), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n946), .ZN(new_n948));
  OAI211_X1 g0748(.A(KEYINPUT102), .B(new_n948), .C1(new_n676), .C2(new_n839), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n943), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n930), .A2(new_n931), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n651), .A2(new_n686), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n938), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n735), .A2(new_n736), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n689), .B1(new_n843), .B2(new_n845), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT95), .B1(new_n956), .B2(new_n725), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n723), .A2(new_n716), .A3(KEYINPUT29), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n460), .B(new_n955), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n653), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n954), .B(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT40), .ZN(new_n962));
  INV_X1    g0762(.A(new_n848), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n940), .B2(new_n941), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n759), .B(new_n964), .C1(new_n930), .C2(new_n931), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n964), .A2(new_n759), .A3(KEYINPUT40), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n903), .A2(new_n923), .A3(new_n924), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n962), .A2(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n460), .A3(new_n759), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(G330), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n968), .B1(new_n460), .B2(new_n759), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n961), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n207), .B2(new_n764), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n961), .A2(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n887), .B1(new_n974), .B2(new_n975), .ZN(G367));
  NOR2_X1   g0776(.A1(new_n772), .A2(new_n773), .ZN(new_n977));
  INV_X1    g0777(.A(new_n776), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n977), .B1(new_n211), .B2(new_n409), .C1(new_n978), .C2(new_n240), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n768), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n792), .A2(G116), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  INV_X1    g0782(.A(new_n806), .ZN(new_n983));
  XOR2_X1   g0783(.A(KEYINPUT111), .B(G317), .Z(new_n984));
  AOI22_X1  g0784(.A1(G97), .A2(new_n983), .B1(new_n788), .B2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G303), .A2(new_n784), .B1(new_n819), .B2(G283), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n982), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n803), .A2(G107), .B1(G311), .B2(new_n804), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n988), .B(new_n870), .C1(new_n855), .C2(new_n817), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G50), .A2(new_n819), .B1(new_n788), .B2(G137), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n313), .B2(new_n806), .C1(new_n863), .C2(new_n783), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n802), .A2(new_n298), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n804), .B2(G143), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n277), .B1(new_n792), .B2(G58), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n343), .C2(new_n817), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n987), .A2(new_n989), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n980), .B1(new_n997), .B2(new_n773), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n617), .A2(new_n618), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n688), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n656), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n670), .A2(new_n999), .A3(new_n688), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n998), .B1(new_n827), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT112), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n511), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n522), .B1(new_n682), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT89), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n512), .A2(new_n513), .A3(new_n522), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n690), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n693), .B(KEYINPUT92), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n706), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n706), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n692), .A2(new_n695), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT110), .B1(new_n699), .B2(G330), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n737), .A2(new_n1018), .A3(new_n761), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n575), .A2(new_n688), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n654), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n665), .A2(new_n688), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1020), .B1(new_n707), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n705), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1012), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1024), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(KEYINPUT44), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1012), .A2(new_n1026), .A3(new_n1024), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1012), .A2(KEYINPUT45), .A3(new_n1026), .A4(new_n1024), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT109), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1019), .B1(new_n1036), .B2(new_n703), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1025), .A2(new_n1029), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1038), .A2(KEYINPUT109), .A3(new_n704), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n762), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n710), .B(KEYINPUT41), .Z(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n766), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1013), .B1(new_n692), .B2(new_n695), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1024), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT42), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n598), .B1(new_n1022), .B2(new_n512), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1045), .A2(KEYINPUT42), .B1(new_n689), .B2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1046), .A2(new_n1048), .B1(KEYINPUT43), .B2(new_n1003), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1003), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT43), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1046), .A2(new_n1048), .A3(new_n1051), .A4(new_n1050), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n704), .A2(new_n1028), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1055), .B(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1005), .B1(new_n1043), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1055), .B(new_n1056), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1036), .A2(new_n703), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n704), .B1(new_n1038), .B2(KEYINPUT109), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n1063), .A3(new_n1019), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1041), .B1(new_n1064), .B2(new_n762), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1061), .B1(new_n1065), .B2(new_n766), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT113), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n1005), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1060), .A2(new_n1068), .ZN(G387));
  NOR2_X1   g0869(.A1(new_n1019), .A2(new_n711), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n762), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n778), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1073), .A2(new_n712), .B1(G107), .B2(new_n211), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n237), .A2(G45), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT114), .Z(new_n1076));
  OAI21_X1  g0876(.A(new_n260), .B1(new_n298), .B2(new_n313), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n326), .A2(new_n202), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT50), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(KEYINPUT50), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n978), .B1(new_n1081), .B2(new_n712), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1074), .B1(new_n1076), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n977), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n768), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n696), .A2(new_n827), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G68), .A2(new_n819), .B1(new_n788), .B2(G150), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n202), .B2(new_n783), .C1(new_n313), .C2(new_n791), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n870), .B1(new_n326), .B2(new_n799), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n343), .B2(new_n821), .C1(new_n409), .C2(new_n802), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(G97), .C2(new_n807), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT115), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n784), .A2(new_n984), .B1(new_n819), .B2(G303), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT116), .B(G322), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1093), .B1(new_n821), .B2(new_n1094), .C1(new_n796), .C2(new_n817), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT48), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(G283), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n791), .A2(new_n855), .B1(new_n802), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT49), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1097), .A2(KEYINPUT49), .A3(new_n1100), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G116), .A2(new_n983), .B1(new_n788), .B2(G326), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n870), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1092), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1085), .B(new_n1086), .C1(new_n773), .C2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n766), .B2(new_n1071), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1072), .A2(new_n1107), .ZN(G393));
  AOI21_X1  g0908(.A(KEYINPUT44), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1020), .B(new_n1024), .C1(new_n1012), .C2(new_n1026), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT45), .B1(new_n707), .B2(new_n1024), .ZN(new_n1111));
  NOR4_X1   g0911(.A1(new_n1044), .A2(new_n1032), .A3(new_n705), .A4(new_n1028), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1109), .A2(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n704), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n1071), .A3(new_n760), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1030), .A2(new_n1035), .A3(new_n703), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n710), .C1(new_n1037), .C2(new_n1039), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n977), .B1(new_n249), .B2(new_n211), .C1(new_n978), .C2(new_n253), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n768), .A2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n784), .A2(G159), .B1(G150), .B2(new_n804), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT51), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n870), .B1(G50), .B2(new_n799), .ZN(new_n1124));
  INV_X1    g0924(.A(G143), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n791), .A2(new_n298), .B1(new_n787), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n326), .B2(new_n819), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n803), .A2(G77), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1124), .A2(new_n859), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n369), .B1(new_n819), .B2(G294), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1094), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G283), .A2(new_n792), .B1(new_n788), .B2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n803), .A2(G116), .B1(G303), .B2(new_n799), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n810), .A2(new_n1130), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n784), .A2(G311), .B1(G317), .B2(new_n804), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT52), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1123), .A2(new_n1129), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1121), .B1(new_n1137), .B2(new_n773), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1024), .B2(new_n827), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT117), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1030), .A2(new_n1035), .A3(new_n703), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n703), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1114), .A2(KEYINPUT117), .A3(new_n1117), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n1144), .A3(new_n766), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1119), .A2(new_n1139), .A3(new_n1145), .ZN(G390));
  NAND4_X1  g0946(.A1(new_n759), .A2(G330), .A3(new_n848), .A4(new_n942), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT102), .B1(new_n846), .B2(new_n948), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n945), .A2(new_n944), .A3(new_n946), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n942), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n934), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1151), .A2(new_n1152), .B1(new_n933), .B2(new_n937), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n733), .B1(new_n728), .B2(new_n721), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n948), .B1(new_n1154), .B2(new_n839), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n942), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n1152), .A3(new_n967), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1148), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n933), .A2(new_n937), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n950), .A2(new_n934), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1147), .B(new_n1157), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n759), .A2(G330), .A3(new_n848), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n943), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n946), .B1(new_n735), .B2(new_n840), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1147), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1165), .A2(new_n1147), .B1(new_n947), .B2(new_n949), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n460), .A2(new_n761), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n959), .A2(new_n653), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1163), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1159), .A2(new_n1176), .A3(new_n1162), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n710), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1159), .A2(new_n766), .A3(new_n1162), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n768), .B1(new_n326), .B2(new_n852), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n791), .A2(new_n863), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT53), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G132), .A2(new_n784), .B1(new_n788), .B2(G125), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT54), .B(G143), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1182), .B(new_n1183), .C1(new_n795), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n277), .B1(new_n983), .B2(G50), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G128), .A2(new_n804), .B1(new_n799), .B2(G137), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n343), .C2(new_n802), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n369), .B1(new_n784), .B2(G116), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G87), .A2(new_n792), .B1(new_n788), .B2(G294), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n803), .A2(G77), .B1(G283), .B2(new_n804), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n867), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n817), .A2(new_n247), .B1(new_n795), .B2(new_n249), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT118), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n1185), .A2(new_n1188), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1180), .B1(new_n1195), .B2(new_n773), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1160), .B2(new_n771), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1179), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1178), .A2(new_n1199), .ZN(G378));
  NOR2_X1   g1000(.A1(new_n775), .A2(G41), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G50), .B(new_n1201), .C1(new_n336), .C2(new_n259), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n806), .A2(new_n243), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G283), .B2(new_n788), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n1201), .C1(new_n409), .C2(new_n795), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n817), .A2(new_n249), .B1(new_n821), .B2(new_n216), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n313), .A2(new_n791), .B1(new_n783), .B2(new_n247), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n992), .A4(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1202), .B1(new_n1208), .B2(KEYINPUT58), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n817), .A2(new_n868), .B1(new_n802), .B2(new_n863), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1184), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G128), .A2(new_n784), .B1(new_n792), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n862), .B2(new_n795), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1210), .B(new_n1213), .C1(G125), .C2(new_n804), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n336), .B(new_n259), .C1(new_n806), .C2(new_n343), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G124), .B2(new_n788), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT59), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1218), .B1(new_n1214), .B2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1209), .B1(KEYINPUT58), .B2(new_n1208), .C1(new_n1216), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n773), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n767), .C1(G50), .C2(new_n852), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n457), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n457), .A2(new_n1224), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n446), .A2(new_n686), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT119), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OR3_X1    g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1223), .B1(new_n1232), .B2(new_n770), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT120), .Z(new_n1234));
  AOI21_X1  g1034(.A(new_n1232), .B1(new_n968), .B2(G330), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n965), .A2(new_n962), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n966), .A2(new_n967), .ZN(new_n1237));
  AND4_X1   g1037(.A1(G330), .A2(new_n1236), .A3(new_n1237), .A4(new_n1232), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n954), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(G330), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1232), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n950), .A2(new_n951), .B1(new_n651), .B2(new_n686), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1236), .A2(new_n1237), .A3(new_n1232), .A4(G330), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1242), .A2(new_n938), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1239), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1234), .B1(new_n1246), .B2(new_n765), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1177), .A2(new_n1173), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1239), .A2(KEYINPUT57), .A3(new_n1245), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n710), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1246), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1248), .B1(new_n1252), .B2(new_n1254), .ZN(G375));
  NAND2_X1  g1055(.A1(new_n943), .A2(new_n770), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n768), .B1(G68), .B2(new_n852), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G159), .A2(new_n792), .B1(new_n788), .B2(G128), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT122), .Z(new_n1259));
  AOI21_X1  g1059(.A(new_n870), .B1(G132), .B2(new_n804), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n819), .A2(G150), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1203), .B1(G137), .B2(new_n784), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G50), .A2(new_n803), .B1(new_n1211), .B2(new_n799), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n819), .A2(G107), .B1(G116), .B2(new_n799), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT121), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n807), .A2(G77), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n369), .B1(new_n784), .B2(G283), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G97), .A2(new_n792), .B1(new_n788), .B2(G303), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n803), .A2(new_n599), .B1(G294), .B2(new_n804), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1259), .A2(new_n1264), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1257), .B1(new_n1272), .B2(new_n773), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1170), .A2(new_n766), .B1(new_n1256), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1176), .A2(new_n1041), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(G381));
  NAND3_X1  g1079(.A1(new_n1072), .A2(new_n831), .A3(new_n1107), .ZN(new_n1280));
  OR4_X1    g1080(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1280), .ZN(new_n1281));
  OR4_X1    g1081(.A1(G387), .A2(new_n1281), .A3(G378), .A4(G375), .ZN(G407));
  AOI21_X1  g1082(.A(new_n711), .B1(new_n1163), .B2(new_n1174), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1198), .B1(new_n1283), .B2(new_n1177), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n687), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G407), .B(G213), .C1(G375), .C2(new_n1285), .ZN(G409));
  OAI211_X1 g1086(.A(G390), .B(new_n1005), .C1(new_n1043), .C2(new_n1058), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G390), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1059), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1066), .A2(KEYINPUT124), .A3(new_n1005), .A4(G390), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1289), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1280), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1060), .A2(new_n1068), .A3(new_n1290), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1287), .A2(new_n1295), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G378), .B(new_n1248), .C1(new_n1252), .C2(new_n1254), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1249), .A2(new_n1042), .A3(new_n1253), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1248), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1284), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(G213), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1308), .A2(G343), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1277), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT60), .B1(new_n1277), .B2(KEYINPUT123), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n710), .B(new_n1174), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(G384), .A3(new_n1274), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1174), .A2(new_n710), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1277), .A2(KEYINPUT123), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1320), .B2(new_n1312), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n877), .B1(new_n1321), .B2(new_n1275), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1309), .A2(G2897), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1316), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1316), .B2(new_n1322), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1311), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1302), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1316), .A2(new_n1322), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1307), .A2(new_n1310), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(KEYINPUT62), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1309), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT62), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1335), .A3(new_n1331), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1333), .A2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1301), .B1(new_n1329), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT63), .B1(new_n1334), .B2(new_n1331), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1339), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1297), .A2(KEYINPUT125), .A3(new_n1300), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1323), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1330), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1316), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1328), .B1(new_n1347), .B2(new_n1334), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1343), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1342), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1338), .A2(new_n1350), .ZN(G405));
  NAND2_X1  g1151(.A1(new_n1301), .A2(KEYINPUT126), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1284), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1303), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1331), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1353), .A2(new_n1303), .A3(new_n1330), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT126), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1339), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1352), .A2(new_n1357), .A3(new_n1359), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1360), .B1(new_n1359), .B2(new_n1357), .ZN(G402));
endmodule


