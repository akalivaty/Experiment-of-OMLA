//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n212, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT65), .B(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G87), .ZN(G355));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n214), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT66), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n223), .B1(new_n214), .B2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G13), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n225), .A2(KEYINPUT66), .A3(G1), .A4(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G50), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n206), .A2(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n222), .B(new_n229), .C1(new_n232), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G244), .A3(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(G238), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G116), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n252), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n266), .B(new_n260), .C1(G250), .C2(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G190), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(G200), .B2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n251), .A2(new_n231), .A3(G68), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n255), .A2(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G97), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT19), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G97), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n231), .B1(new_n277), .B2(new_n275), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G87), .B2(new_n212), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n272), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n280), .A2(KEYINPUT88), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(new_n230), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n280), .B2(KEYINPUT88), .ZN(new_n284));
  XOR2_X1   g0084(.A(KEYINPUT15), .B(G87), .Z(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n225), .A2(new_n231), .A3(G1), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n281), .A2(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT67), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(new_n289), .A3(new_n230), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n282), .B2(new_n230), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n291), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT79), .ZN(new_n294));
  INV_X1    g0094(.A(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G33), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n292), .ZN(new_n298));
  INV_X1    g0098(.A(new_n287), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(new_n290), .A4(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT79), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G87), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n288), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n285), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n262), .A2(new_n267), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n288), .A2(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n268), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n271), .A2(new_n304), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT84), .ZN(new_n313));
  INV_X1    g0113(.A(G41), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n295), .B(G45), .C1(new_n314), .C2(KEYINPUT5), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT83), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT5), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G41), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT83), .B1(new_n264), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n313), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n295), .A2(G45), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n316), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n264), .A2(KEYINPUT83), .A3(new_n319), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(KEYINPUT84), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n318), .A2(KEYINPUT85), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT85), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT5), .ZN(new_n329));
  AOI21_X1  g0129(.A(G41), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n259), .ZN(new_n331));
  OAI21_X1  g0131(.A(G274), .B1(new_n331), .B2(new_n230), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n321), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n327), .A2(new_n329), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n324), .B(new_n325), .C1(new_n335), .C2(G41), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G257), .A3(new_n260), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(new_n253), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT4), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G250), .A2(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(KEYINPUT4), .A2(G244), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G283), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT81), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT81), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(G33), .A3(G283), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n251), .A2(new_n347), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT82), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n344), .A2(new_n352), .A3(KEYINPUT82), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n261), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n338), .A2(G179), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n309), .B1(new_n338), .B2(new_n357), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n210), .B1(new_n297), .B2(new_n301), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n282), .A2(new_n230), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT6), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n363), .A2(new_n210), .A3(G107), .ZN(new_n364));
  XNOR2_X1  g0164(.A(G97), .B(G107), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n363), .ZN(new_n366));
  INV_X1    g0166(.A(G77), .ZN(new_n367));
  NOR2_X1   g0167(.A1(G20), .A2(G33), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n366), .A2(new_n231), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n251), .B2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n339), .A2(new_n341), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n211), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n362), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n287), .A2(new_n210), .ZN(new_n377));
  XOR2_X1   g0177(.A(new_n377), .B(KEYINPUT78), .Z(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n359), .A2(new_n360), .B1(new_n361), .B2(new_n379), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n355), .A2(new_n261), .A3(new_n356), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n334), .A2(new_n337), .ZN(new_n382));
  OAI21_X1  g0182(.A(G200), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n383), .A2(KEYINPUT86), .B1(new_n384), .B2(G190), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT80), .B1(new_n379), .B2(new_n361), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n302), .A2(G97), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT80), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(new_n376), .A4(new_n378), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n338), .A2(new_n357), .A3(KEYINPUT86), .A4(G190), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n380), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT87), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT87), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n380), .B(new_n394), .C1(new_n385), .C2(new_n391), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n312), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n295), .A2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n293), .A2(G50), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(G50), .B2(new_n299), .ZN(new_n399));
  AND2_X1   g0199(.A1(KEYINPUT69), .A2(G58), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT8), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(KEYINPUT68), .A2(KEYINPUT69), .A3(G58), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT8), .B1(KEYINPUT68), .B2(G58), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n273), .B1(G150), .B2(new_n368), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n208), .A2(G20), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n406), .A2(new_n407), .B1(new_n298), .B2(new_n290), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n399), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n339), .A2(new_n341), .A3(G1698), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(G223), .B1(G77), .B2(new_n373), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n251), .A2(G222), .A3(new_n253), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n261), .ZN(new_n414));
  AOI21_X1  g0214(.A(G1), .B1(new_n314), .B2(new_n263), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n260), .A2(G274), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n314), .A2(new_n263), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n295), .A2(new_n418), .B1(new_n258), .B2(new_n259), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(G226), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n409), .B1(new_n309), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n414), .A2(new_n307), .A3(new_n420), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n409), .A2(KEYINPUT9), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT71), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n414), .A2(G190), .A3(new_n420), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT72), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n409), .A2(KEYINPUT9), .B1(new_n421), .B2(G200), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(KEYINPUT10), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(KEYINPUT10), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n424), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n410), .A2(G238), .B1(G107), .B2(new_n373), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n251), .A2(G232), .A3(new_n253), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n261), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT70), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n417), .B1(G244), .B2(new_n419), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n437), .B2(new_n439), .ZN(new_n442));
  OAI21_X1  g0242(.A(G190), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n442), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(G200), .A3(new_n440), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n285), .A2(new_n273), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT8), .B(G58), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n446), .B1(new_n231), .B2(new_n367), .C1(new_n369), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n362), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n287), .A2(new_n362), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n367), .B1(new_n295), .B2(G20), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n450), .A2(new_n451), .B1(new_n367), .B2(new_n287), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n443), .A2(new_n445), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n307), .B1(new_n441), .B2(new_n442), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n444), .A2(new_n309), .A3(new_n440), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(new_n453), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n273), .A2(G77), .ZN(new_n460));
  OAI221_X1 g0260(.A(new_n460), .B1(new_n231), .B2(G68), .C1(new_n233), .C2(new_n369), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n298), .A2(new_n290), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT74), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT11), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT74), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n466), .B1(new_n465), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n287), .A2(new_n202), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT12), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n450), .A2(G68), .A3(new_n397), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OR3_X1    g0273(.A1(new_n468), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT14), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n339), .A2(new_n341), .A3(G226), .A4(new_n253), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n277), .A3(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n478), .A2(new_n261), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT73), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n416), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n260), .A2(new_n415), .A3(KEYINPUT73), .A4(G274), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n419), .A2(G238), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n479), .A2(KEYINPUT13), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT13), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n478), .A2(new_n261), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n475), .B(G169), .C1(new_n485), .C2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT13), .B1(new_n479), .B2(new_n484), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(new_n486), .A3(new_n488), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(G179), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n475), .B1(new_n495), .B2(G169), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n474), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n468), .A2(new_n469), .A3(new_n473), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(G200), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n498), .B(new_n499), .C1(new_n269), .C2(new_n495), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n405), .A2(new_n397), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT76), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT76), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n405), .A2(new_n504), .A3(new_n397), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n293), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n405), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n287), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(KEYINPUT68), .A2(G58), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT68), .A2(G58), .ZN(new_n511));
  OAI21_X1  g0311(.A(G68), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT75), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n206), .ZN(new_n515));
  OAI211_X1 g0315(.A(KEYINPUT75), .B(G68), .C1(new_n510), .C2(new_n511), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n368), .A2(G159), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT7), .B1(new_n373), .B2(new_n231), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n371), .B(G20), .C1(new_n339), .C2(new_n341), .ZN(new_n521));
  OAI21_X1  g0321(.A(G68), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT16), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n517), .A2(G20), .B1(G159), .B2(new_n368), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n372), .A2(new_n374), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n527), .B2(G68), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n283), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n509), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT77), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n339), .A2(new_n341), .A3(G223), .A4(new_n253), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n339), .A2(new_n341), .A3(G226), .A4(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G87), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n261), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n295), .B1(G41), .B2(G45), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n260), .A2(G232), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n416), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n536), .A2(new_n269), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(G200), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n531), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n536), .A2(new_n539), .A3(new_n269), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n416), .A2(new_n538), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n261), .B2(new_n535), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n543), .B(KEYINPUT77), .C1(new_n545), .C2(G200), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n530), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT17), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(G179), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n309), .B2(new_n545), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT18), .B1(new_n530), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n509), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n518), .A2(KEYINPUT16), .A3(new_n522), .A4(new_n519), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n362), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT16), .B1(new_n526), .B2(new_n522), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT18), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n552), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n530), .A2(new_n547), .A3(KEYINPUT17), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n550), .A2(new_n554), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n433), .A2(new_n459), .A3(new_n501), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n324), .A2(new_n325), .ZN(new_n567));
  OAI211_X1 g0367(.A(G264), .B(new_n260), .C1(new_n567), .C2(new_n330), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT92), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n336), .A2(KEYINPUT92), .A3(G264), .A4(new_n260), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n253), .A2(G257), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(G250), .B2(G1698), .ZN(new_n573));
  INV_X1    g0373(.A(G294), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n573), .A2(new_n373), .B1(new_n255), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n570), .A2(new_n571), .B1(new_n261), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(G179), .A3(new_n334), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n261), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n334), .A2(new_n578), .A3(new_n568), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G169), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n339), .A2(new_n341), .A3(new_n231), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT22), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT22), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n251), .A2(new_n583), .A3(new_n231), .A4(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT23), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n211), .A3(G20), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT23), .B1(new_n231), .B2(G107), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT91), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n586), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT24), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n585), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n585), .B2(new_n593), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n362), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n287), .A2(new_n211), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT25), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n302), .B2(G107), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n577), .A2(new_n580), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT93), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n579), .A2(G190), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n570), .A2(new_n571), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n334), .A3(new_n578), .ZN(new_n605));
  INV_X1    g0405(.A(G200), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n600), .A2(new_n597), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n602), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n600), .A2(new_n597), .ZN(new_n610));
  AOI21_X1  g0410(.A(G200), .B1(new_n576), .B2(new_n334), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n610), .B(KEYINPUT93), .C1(new_n611), .C2(new_n603), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n601), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n336), .A2(G270), .A3(new_n260), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n334), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT90), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n339), .A2(new_n341), .A3(G264), .A4(G1698), .ZN(new_n617));
  INV_X1    g0417(.A(G303), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n251), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT89), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n251), .A2(new_n620), .A3(G257), .A4(new_n253), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n339), .A2(new_n341), .A3(G257), .A4(new_n253), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT89), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n619), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n616), .B1(new_n624), .B2(new_n260), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n621), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n410), .A2(G264), .B1(G303), .B2(new_n373), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(KEYINPUT90), .A3(new_n261), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n615), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n231), .A2(G116), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n283), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n349), .A2(new_n351), .ZN(new_n633));
  AOI21_X1  g0433(.A(G20), .B1(new_n255), .B2(G97), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n632), .A2(new_n635), .A3(KEYINPUT20), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n256), .B1(new_n295), .B2(G33), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n225), .A2(G1), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n450), .A2(new_n641), .B1(new_n642), .B2(new_n631), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G169), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT21), .B1(new_n630), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n615), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT90), .B1(new_n628), .B2(new_n261), .ZN(new_n648));
  AOI211_X1 g0448(.A(new_n616), .B(new_n260), .C1(new_n626), .C2(new_n627), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT21), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n309), .B1(new_n640), .B2(new_n643), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n630), .A2(G179), .A3(new_n644), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n647), .B(G190), .C1(new_n648), .C2(new_n649), .ZN(new_n656));
  INV_X1    g0456(.A(new_n644), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n656), .B(new_n657), .C1(new_n606), .C2(new_n630), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n654), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n396), .A2(new_n566), .A3(new_n613), .A4(new_n659), .ZN(G372));
  NAND2_X1  g0460(.A1(new_n431), .A2(new_n432), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n550), .A2(new_n562), .ZN(new_n662));
  INV_X1    g0462(.A(new_n458), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n500), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(new_n497), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n554), .A2(new_n561), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n424), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n288), .A2(new_n305), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n306), .A2(new_n307), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n267), .B(KEYINPUT94), .Z(new_n672));
  INV_X1    g0472(.A(new_n262), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n309), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n386), .A2(new_n389), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n338), .A2(new_n357), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G169), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n358), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n306), .A2(G190), .ZN(new_n680));
  OAI21_X1  g0480(.A(G200), .B1(new_n672), .B2(new_n673), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n288), .A4(new_n303), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n675), .A2(new_n676), .A3(new_n679), .A4(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(KEYINPUT95), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n379), .A2(new_n361), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n678), .B2(new_n358), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n311), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n685), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT95), .B1(new_n683), .B2(new_n684), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n675), .A2(new_n682), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n609), .B2(new_n612), .ZN(new_n693));
  INV_X1    g0493(.A(new_n601), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n654), .A3(new_n655), .ZN(new_n695));
  INV_X1    g0495(.A(new_n391), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n338), .A2(G190), .A3(new_n357), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n606), .B1(new_n338), .B2(new_n357), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT86), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n687), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n693), .A2(new_n695), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n675), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n691), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n669), .B1(new_n566), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT96), .Z(G369));
  NAND2_X1  g0506(.A1(new_n642), .A2(new_n231), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G213), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G343), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n654), .B2(new_n655), .ZN(new_n713));
  INV_X1    g0513(.A(new_n712), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n613), .A2(new_n713), .B1(new_n601), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n654), .A2(new_n655), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n657), .A2(new_n714), .ZN(new_n717));
  MUX2_X1   g0517(.A(new_n659), .B(new_n716), .S(new_n717), .Z(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n608), .A2(new_n712), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n613), .A2(new_n720), .B1(new_n601), .B2(new_n712), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n715), .B1(new_n719), .B2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n227), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(G87), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n210), .A3(new_n211), .A4(new_n256), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n724), .A2(new_n295), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n234), .B2(new_n724), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT28), .Z(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n704), .A2(new_n730), .A3(new_n714), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n683), .A2(KEYINPUT26), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n311), .A2(new_n684), .A3(new_n687), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n702), .A2(new_n675), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n714), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G330), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n613), .A2(new_n659), .A3(new_n714), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n396), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n630), .A2(new_n306), .A3(new_n576), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n742), .B2(new_n358), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n576), .A2(new_n306), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n359), .A3(KEYINPUT30), .A4(new_n630), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n672), .A2(new_n673), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G179), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n650), .A3(new_n605), .A4(new_n677), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n743), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n749), .B2(new_n712), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n738), .B1(new_n740), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n737), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n729), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(new_n225), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n295), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n724), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n227), .A2(G355), .A3(new_n251), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G116), .B2(new_n227), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n249), .A2(G45), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n227), .A2(new_n373), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n263), .B2(new_n234), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n230), .B1(G20), .B2(new_n309), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n761), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n231), .A2(new_n269), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G179), .A3(new_n606), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n606), .A2(G179), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n776), .A2(new_n777), .B1(new_n779), .B2(new_n618), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n231), .A2(new_n307), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(new_n269), .A3(new_n606), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n251), .B(new_n780), .C1(G311), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT100), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n231), .B2(G190), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n269), .A2(KEYINPUT100), .A3(G20), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G329), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n786), .A2(new_n788), .A3(new_n778), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n784), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n781), .A2(G200), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n269), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n231), .B1(new_n787), .B2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n799), .A2(G326), .B1(G294), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT102), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n798), .A2(G190), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n796), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT103), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(KEYINPUT103), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G50), .A2(new_n799), .B1(new_n804), .B2(G68), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n792), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n813), .A2(G77), .B1(G107), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n789), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n510), .A2(new_n511), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n251), .B1(new_n779), .B2(new_n725), .C1(new_n820), .C2(new_n776), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G97), .B2(new_n801), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n809), .A2(new_n815), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n807), .A2(new_n808), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n774), .B1(new_n824), .B2(new_n771), .ZN(new_n825));
  INV_X1    g0625(.A(new_n770), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n718), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n718), .A2(G330), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT97), .Z(new_n829));
  INV_X1    g0629(.A(new_n761), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n719), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT104), .Z(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n704), .A2(new_n714), .ZN(new_n835));
  AND4_X1   g0635(.A1(new_n453), .A2(new_n456), .A3(new_n457), .A4(new_n714), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n453), .A2(new_n712), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n455), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n836), .B1(new_n458), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n714), .B(new_n839), .C1(new_n691), .C2(new_n703), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n761), .B1(new_n843), .B2(new_n754), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n753), .A3(new_n842), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n771), .A2(new_n768), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n814), .A2(G87), .ZN(new_n849));
  INV_X1    g0649(.A(G311), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n850), .B2(new_n789), .C1(new_n812), .C2(new_n256), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n373), .B1(new_n779), .B2(new_n211), .C1(new_n574), .C2(new_n776), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G97), .B2(new_n801), .ZN(new_n853));
  INV_X1    g0653(.A(new_n804), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n793), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n851), .B(new_n855), .C1(G303), .C2(new_n799), .ZN(new_n856));
  INV_X1    g0656(.A(new_n776), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n813), .A2(G159), .B1(G143), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  INV_X1    g0659(.A(new_n799), .ZN(new_n860));
  INV_X1    g0660(.A(G150), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n858), .B1(new_n859), .B2(new_n860), .C1(new_n861), .C2(new_n854), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT34), .Z(new_n863));
  INV_X1    g0663(.A(KEYINPUT105), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n792), .A2(new_n202), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n251), .B1(new_n800), .B2(new_n820), .C1(new_n233), .C2(new_n779), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n866), .B(new_n867), .C1(G132), .C2(new_n790), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n863), .B2(new_n864), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n856), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n771), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n761), .B1(G77), .B2(new_n848), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n768), .B2(new_n840), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n846), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  INV_X1    g0676(.A(new_n366), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n232), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n234), .A2(G77), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n514), .A2(new_n516), .ZN(new_n883));
  INV_X1    g0683(.A(new_n207), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n882), .A2(new_n883), .B1(new_n202), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n295), .A2(G13), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n559), .A2(new_n552), .ZN(new_n888));
  INV_X1    g0688(.A(new_n710), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n559), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n890), .A3(new_n548), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n888), .A2(new_n890), .A3(new_n548), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n890), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n895), .A2(KEYINPUT109), .B1(new_n563), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT109), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n892), .A2(new_n898), .A3(new_n894), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n556), .A2(new_n462), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n555), .B1(new_n902), .B2(new_n558), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n552), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n548), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n903), .A2(new_n889), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n894), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n563), .A2(KEYINPUT108), .A3(new_n906), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT108), .B1(new_n563), .B2(new_n906), .ZN(new_n910));
  OAI211_X1 g0710(.A(KEYINPUT38), .B(new_n908), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT39), .B1(new_n901), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n497), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n714), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n497), .A2(KEYINPUT107), .A3(new_n500), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n474), .A2(new_n712), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT107), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n497), .A2(new_n926), .A3(new_n500), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n924), .A2(new_n494), .A3(new_n496), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n836), .B(KEYINPUT106), .Z(new_n931));
  AOI21_X1  g0731(.A(new_n930), .B1(new_n842), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n915), .A2(new_n911), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n666), .A2(new_n710), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n922), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n565), .B1(new_n731), .B2(new_n736), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(new_n669), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n936), .B(new_n938), .Z(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT110), .ZN(new_n941));
  INV_X1    g0741(.A(new_n751), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n943));
  INV_X1    g0743(.A(new_n395), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n700), .A2(new_n386), .A3(new_n389), .A4(new_n390), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n394), .B1(new_n945), .B2(new_n380), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n311), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n613), .A2(new_n659), .A3(new_n714), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n942), .B(new_n943), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n925), .A2(new_n929), .A3(new_n839), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n911), .B2(new_n915), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n941), .B1(new_n953), .B2(KEYINPUT40), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n950), .B1(new_n740), .B2(new_n752), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n933), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(KEYINPUT110), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n911), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n955), .B(KEYINPUT40), .C1(new_n959), .C2(new_n900), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT111), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n895), .A2(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n563), .A2(new_n896), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n962), .A2(new_n899), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n911), .B1(new_n964), .B2(KEYINPUT38), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT111), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT40), .A4(new_n955), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n954), .A2(new_n958), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n565), .B1(new_n740), .B2(new_n752), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n970), .A2(new_n971), .A3(new_n738), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n940), .A2(new_n972), .B1(new_n295), .B2(new_n758), .ZN(new_n973));
  INV_X1    g0773(.A(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n939), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n887), .B1(new_n973), .B2(new_n975), .ZN(G367));
  NAND2_X1  g0776(.A1(new_n676), .A2(new_n712), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n701), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n676), .A2(new_n679), .A3(new_n712), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n613), .A3(new_n713), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT42), .Z(new_n982));
  INV_X1    g0782(.A(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n380), .B1(new_n983), .B2(new_n694), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n714), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n304), .A2(new_n714), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(new_n308), .A3(new_n674), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n692), .B2(new_n986), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n982), .A2(new_n985), .B1(KEYINPUT43), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n719), .A2(new_n721), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n980), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n991), .B(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n724), .B(KEYINPUT41), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n980), .A2(new_n715), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n992), .A2(KEYINPUT114), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n980), .A2(new_n715), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n992), .A2(KEYINPUT114), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  MUX2_X1   g0804(.A(new_n721), .B(new_n613), .S(new_n713), .Z(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(new_n719), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n756), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1004), .B1(new_n1008), .B2(KEYINPUT113), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(KEYINPUT113), .B2(new_n1008), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n995), .B1(new_n1010), .B2(new_n756), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n994), .B1(new_n1011), .B2(new_n760), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n242), .A2(new_n765), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n772), .B1(new_n227), .B2(new_n286), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n761), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n792), .A2(new_n367), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n251), .B1(new_n800), .B2(new_n202), .C1(new_n776), .C2(new_n861), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n813), .C2(new_n884), .ZN(new_n1018));
  INV_X1    g0818(.A(G143), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n860), .C1(new_n816), .C2(new_n854), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n789), .A2(new_n859), .B1(new_n779), .B2(new_n820), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT115), .Z(new_n1022));
  OAI221_X1 g0822(.A(new_n373), .B1(new_n800), .B2(new_n211), .C1(new_n776), .C2(new_n618), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n779), .A2(new_n256), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT46), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(G311), .C2(new_n799), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n574), .B2(new_n854), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n813), .A2(G283), .B1(G97), .B2(new_n814), .ZN(new_n1028));
  INV_X1    g0828(.A(G317), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n789), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1020), .A2(new_n1022), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT47), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1015), .B1(new_n1032), .B2(new_n771), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n826), .B2(new_n988), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1012), .A2(new_n1034), .ZN(G387));
  NAND2_X1  g0835(.A1(new_n755), .A2(new_n1006), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1008), .A2(new_n724), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n210), .A2(new_n792), .B1(new_n789), .B2(new_n861), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n286), .A2(new_n800), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n776), .A2(new_n233), .B1(new_n779), .B2(new_n367), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n251), .B1(new_n782), .B2(new_n202), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n860), .B2(new_n816), .C1(new_n507), .C2(new_n854), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n813), .A2(G303), .B1(G317), .B2(new_n857), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n850), .B2(new_n854), .C1(new_n777), .C2(new_n860), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n779), .A2(new_n574), .B1(new_n800), .B2(new_n793), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n251), .B1(new_n790), .B2(G326), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n256), .C2(new_n792), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1050), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n771), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n239), .A2(new_n263), .A3(new_n251), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n447), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1058));
  OAI21_X1  g0858(.A(KEYINPUT50), .B1(new_n447), .B2(G50), .ZN(new_n1059));
  AOI21_X1  g0859(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n726), .B1(new_n1061), .B2(new_n373), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n227), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n773), .B1(new_n723), .B2(G107), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n830), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n721), .B2(new_n770), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n1007), .B2(new_n760), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1037), .A2(new_n1068), .ZN(G393));
  INV_X1    g0869(.A(new_n1004), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n759), .B1(new_n1070), .B2(KEYINPUT117), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(KEYINPUT117), .B2(new_n1070), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n983), .A2(new_n770), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT118), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n246), .A2(new_n227), .A3(new_n373), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n773), .B1(new_n723), .B2(G97), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n830), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n779), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n373), .B1(new_n1078), .B2(G68), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1079), .B(new_n849), .C1(new_n367), .C2(new_n800), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n812), .A2(new_n447), .B1(new_n1019), .B2(new_n789), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n884), .C2(new_n804), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n799), .A2(G150), .B1(G159), .B2(new_n857), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n799), .A2(G317), .B1(G311), .B2(new_n857), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n211), .A2(new_n792), .B1(new_n789), .B2(new_n777), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n251), .B1(new_n783), .B2(G294), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n256), .B2(new_n800), .C1(new_n793), .C2(new_n779), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(G303), .C2(new_n804), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1082), .A2(new_n1085), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1074), .B(new_n1077), .C1(new_n872), .C2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1072), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n724), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1008), .B2(new_n1004), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1010), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1098), .ZN(G390));
  NAND2_X1  g0899(.A1(new_n842), .A2(new_n931), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n930), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n753), .B2(new_n839), .ZN(new_n1102));
  AND4_X1   g0902(.A1(G330), .A2(new_n949), .A3(new_n839), .A4(new_n1101), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT119), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n838), .A2(new_n458), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n734), .A2(new_n714), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n836), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OR3_X1    g0910(.A1(new_n1102), .A2(new_n1103), .A3(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(KEYINPUT119), .B(new_n1100), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1106), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n754), .A2(new_n565), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n937), .A2(new_n669), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT39), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n959), .B2(new_n900), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1117), .A2(new_n920), .B1(new_n1119), .B2(new_n916), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n965), .A2(new_n920), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n930), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1103), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n912), .A2(new_n917), .B1(new_n932), .B2(new_n921), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1103), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1113), .A2(new_n1124), .A3(new_n1128), .A4(new_n1115), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n724), .A3(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(KEYINPUT120), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(KEYINPUT120), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n813), .A2(G97), .B1(new_n799), .B2(G283), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n211), .B2(new_n854), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT121), .Z(new_n1138));
  NOR2_X1   g0938(.A1(new_n800), .A2(new_n367), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n373), .B1(new_n779), .B2(new_n725), .C1(new_n256), .C2(new_n776), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n202), .A2(new_n792), .B1(new_n789), .B2(new_n574), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(G125), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1143), .A2(new_n789), .B1(new_n792), .B2(new_n207), .ZN(new_n1144));
  INV_X1    g0944(.A(G132), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n251), .B1(new_n776), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1078), .A2(G150), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(G159), .C2(new_n801), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n860), .C1(new_n859), .C2(new_n854), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  AOI211_X1 g0952(.A(new_n1144), .B(new_n1151), .C1(new_n813), .C2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n771), .B1(new_n1142), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n830), .B1(new_n507), .B2(new_n847), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n918), .C2(new_n769), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1129), .B2(new_n759), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1135), .A2(new_n1158), .ZN(G378));
  OAI21_X1  g0959(.A(new_n889), .B1(new_n399), .B2(new_n408), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n433), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n433), .B1(new_n409), .B2(new_n710), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1163), .B(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n968), .B2(G330), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n961), .A2(new_n967), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT110), .B1(new_n956), .B2(new_n957), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n941), .B(KEYINPUT40), .C1(new_n933), .C2(new_n955), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(G330), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1166), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n936), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT123), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n936), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n954), .A2(new_n958), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(new_n1166), .A3(G330), .A4(new_n1168), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1174), .A2(new_n1175), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1131), .A2(new_n1115), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT123), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1131), .B2(new_n1115), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1177), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n724), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1181), .A2(new_n760), .A3(new_n1184), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1172), .A2(new_n768), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n761), .B1(new_n884), .B2(new_n848), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(G33), .A2(G41), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G50), .B(new_n1197), .C1(new_n373), .C2(new_n314), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G97), .A2(new_n804), .B1(new_n799), .B2(G116), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n314), .B(new_n373), .C1(new_n779), .C2(new_n367), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n286), .A2(new_n782), .B1(new_n211), .B2(new_n776), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G68), .C2(new_n801), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n820), .A2(new_n792), .B1(new_n789), .B2(new_n793), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1199), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT58), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1198), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1150), .A2(new_n776), .B1(new_n782), .B2(new_n859), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1078), .A2(new_n1152), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT122), .Z(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G150), .C2(new_n801), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n1143), .B2(new_n860), .C1(new_n1145), .C2(new_n854), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1197), .B1(new_n792), .B2(new_n816), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G124), .B2(new_n790), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1207), .B1(new_n1206), .B2(new_n1205), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1196), .B1(new_n1218), .B2(new_n771), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1195), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1194), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1193), .A2(new_n1222), .ZN(G375));
  NOR2_X1   g1023(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n995), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1226), .A3(new_n1116), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n367), .A2(new_n792), .B1(new_n789), .B2(new_n618), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n860), .A2(new_n574), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n854), .A2(new_n256), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n373), .B1(new_n779), .B2(new_n210), .C1(new_n793), .C2(new_n776), .ZN(new_n1231));
  OR4_X1    g1031(.A1(new_n1039), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1228), .B(new_n1232), .C1(G107), .C2(new_n813), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n820), .A2(new_n792), .B1(new_n789), .B2(new_n1150), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n251), .B1(new_n779), .B2(new_n816), .C1(new_n861), .C2(new_n782), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(G50), .C2(new_n801), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT124), .Z(new_n1237));
  AOI22_X1  g1037(.A1(new_n804), .A2(new_n1152), .B1(G137), .B2(new_n857), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1145), .B2(new_n860), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n771), .B1(new_n1233), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n761), .C1(G68), .C2(new_n848), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n930), .B2(new_n768), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1113), .B2(new_n760), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1227), .A2(new_n1244), .ZN(G381));
  NAND4_X1  g1045(.A1(new_n1012), .A2(new_n1034), .A3(new_n1098), .A4(new_n1095), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1132), .A2(new_n1158), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n833), .A2(new_n1037), .A3(new_n1068), .ZN(new_n1248));
  OR3_X1    g1048(.A1(G381), .A2(G384), .A3(new_n1248), .ZN(new_n1249));
  OR4_X1    g1049(.A1(G375), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(G407));
  INV_X1    g1050(.A(new_n1247), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n711), .A2(G213), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT125), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G407), .B(G213), .C1(G375), .C2(new_n1254), .ZN(G409));
  NAND2_X1  g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1248), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G387), .A2(G390), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1260), .B1(new_n1261), .B2(new_n1246), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1246), .A3(new_n1260), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1224), .A2(KEYINPUT60), .A3(new_n1116), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n724), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1224), .B1(KEYINPUT60), .B2(new_n1116), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1244), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n875), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G384), .B(new_n1244), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1191), .B1(new_n1186), .B2(new_n1185), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1157), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1221), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n759), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(new_n1195), .B2(new_n1219), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1181), .A2(new_n1226), .A3(new_n1182), .A4(new_n1184), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1247), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1252), .B(new_n1274), .C1(new_n1277), .C2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1193), .A2(G378), .A3(new_n1222), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1281), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1253), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1273), .A2(new_n1283), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1282), .A2(new_n1283), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  INV_X1    g1089(.A(G2897), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1273), .A2(new_n1290), .A3(new_n1252), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1271), .A2(new_n1272), .B1(G2897), .B2(new_n1253), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1286), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1266), .B1(new_n1288), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1252), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1292), .B2(new_n1291), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1282), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1286), .A2(KEYINPUT63), .A3(new_n1274), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1296), .A2(new_n1298), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1302), .ZN(G405));
  NAND2_X1  g1103(.A1(G375), .A2(new_n1251), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1284), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1274), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1273), .A3(new_n1284), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT127), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1263), .A2(new_n1309), .A3(new_n1264), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1264), .ZN(new_n1311));
  OAI21_X1  g1111(.A(KEYINPUT127), .B1(new_n1311), .B2(new_n1262), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1308), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1306), .A2(new_n1265), .A3(KEYINPUT127), .A4(new_n1307), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(G402));
endmodule


