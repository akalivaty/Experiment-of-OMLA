//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g030(.A(G2105), .ZN(new_n456));
  NAND3_X1  g031(.A1(new_n456), .A2(G101), .A3(G2104), .ZN(new_n457));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(G137), .A3(new_n456), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n456), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n462), .A2(new_n465), .ZN(G160));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n467), .A2(KEYINPUT68), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT68), .B1(new_n467), .B2(new_n468), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n456), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n456), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n471), .A2(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(G136), .B2(new_n477), .ZN(G162));
  INV_X1    g053(.A(G114), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n481));
  AND2_X1   g056(.A1(G126), .A2(G2105), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n483), .B2(new_n484), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n488), .B(new_n491), .C1(new_n484), .C2(new_n483), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n486), .B1(new_n490), .B2(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(G543), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n498), .A2(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT69), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n506), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G166));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  INV_X1    g090(.A(G51), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n502), .B2(new_n516), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT5), .B(G543), .Z(new_n518));
  NAND2_X1  g093(.A1(new_n499), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(G168));
  INV_X1    g097(.A(G90), .ZN(new_n523));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n500), .A2(new_n523), .B1(new_n502), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n525), .B(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n498), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n506), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  NAND2_X1  g106(.A1(G68), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G56), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n518), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n506), .B1(new_n534), .B2(KEYINPUT71), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n535), .B1(KEYINPUT71), .B2(new_n534), .ZN(new_n536));
  AND2_X1   g111(.A1(KEYINPUT6), .A2(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(KEYINPUT6), .A2(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n518), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n495), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(G81), .B1(new_n541), .B2(G43), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  AOI22_X1  g123(.A1(new_n498), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n506), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(KEYINPUT9), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n541), .B(new_n553), .C1(new_n552), .C2(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n540), .A2(G91), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT72), .B(new_n556), .C1(new_n502), .C2(new_n551), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n550), .A2(new_n554), .A3(new_n555), .A4(new_n557), .ZN(G299));
  INV_X1    g133(.A(G168), .ZN(G286));
  OR3_X1    g134(.A1(new_n504), .A2(new_n510), .A3(KEYINPUT73), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT73), .B1(new_n504), .B2(new_n510), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(G303));
  OAI21_X1  g137(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n563));
  INV_X1    g138(.A(G49), .ZN(new_n564));
  INV_X1    g139(.A(G87), .ZN(new_n565));
  OAI221_X1 g140(.A(new_n563), .B1(new_n502), .B2(new_n564), .C1(new_n565), .C2(new_n500), .ZN(G288));
  INV_X1    g141(.A(G61), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n496), .B2(new_n497), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT74), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(G73), .A3(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n498), .A2(new_n499), .A3(G86), .ZN(new_n575));
  OAI211_X1 g150(.A(G48), .B(G543), .C1(new_n537), .C2(new_n538), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n499), .A2(new_n578), .A3(G48), .A4(G543), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n574), .A2(new_n575), .A3(new_n577), .A4(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(G72), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G60), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n518), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n506), .B1(new_n583), .B2(KEYINPUT76), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(KEYINPUT76), .B2(new_n583), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n540), .A2(G85), .B1(new_n541), .B2(G47), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n500), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n518), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n541), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n591), .B1(G868), .B2(new_n601), .ZN(G284));
  OAI21_X1  g177(.A(new_n591), .B1(G868), .B2(new_n601), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n536), .A2(new_n542), .ZN(new_n610));
  INV_X1    g185(.A(new_n601), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT78), .B1(new_n611), .B2(G559), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n601), .A2(new_n613), .A3(new_n608), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n610), .B(new_n615), .S(G868), .Z(G323));
  XOR2_X1   g191(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n617));
  XNOR2_X1  g192(.A(G323), .B(new_n617), .ZN(G282));
  NAND2_X1  g193(.A1(new_n477), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n472), .A2(G123), .ZN(new_n620));
  OR2_X1    g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n621), .B(G2104), .C1(G111), .C2(new_n456), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT80), .B(G2100), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n456), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n624), .A2(new_n625), .A3(new_n630), .ZN(G156));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n635), .B(new_n641), .Z(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n645), .A3(G14), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2072), .B(G2078), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(KEYINPUT17), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT81), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n650), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n655), .A2(new_n648), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n649), .A2(new_n648), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n654), .B(new_n657), .C1(new_n652), .C2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT82), .B(G2100), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n662), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  MUX2_X1   g247(.A(new_n670), .B(new_n668), .S(new_n672), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n667), .A3(KEYINPUT83), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n673), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT85), .B(KEYINPUT86), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G4), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n601), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1348), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(G20), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT23), .Z(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G299), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1956), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n543), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G16), .B2(G19), .ZN(new_n700));
  INV_X1    g275(.A(G1341), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI211_X1 g277(.A(new_n694), .B(new_n702), .C1(new_n701), .C2(new_n700), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G26), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n477), .A2(G140), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n472), .A2(G128), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n456), .A2(G116), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n710), .B1(new_n715), .B2(G29), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2067), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n707), .A2(G35), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G162), .B2(new_n707), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT29), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n703), .B(new_n717), .C1(G2090), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(G2090), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT99), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n477), .A2(G141), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n472), .A2(G129), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n456), .A2(G105), .A3(G2104), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT26), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n728), .A2(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n724), .A2(new_n725), .A3(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G32), .B(new_n735), .S(G29), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT27), .ZN(new_n737));
  INV_X1    g312(.A(G1996), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G160), .A2(G29), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G34), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n708), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n691), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n691), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT94), .B(G1966), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n745), .A2(new_n746), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n748), .A2(new_n750), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT30), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n755));
  OR2_X1    g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  NAND2_X1  g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n623), .A2(new_n708), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT95), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n752), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n751), .B(new_n761), .C1(new_n746), .C2(new_n745), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n691), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n691), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n456), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n456), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n477), .B2(G139), .ZN(new_n773));
  MUX2_X1   g348(.A(new_n768), .B(new_n773), .S(G29), .Z(new_n774));
  INV_X1    g349(.A(G2072), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n774), .A2(new_n775), .B1(new_n760), .B2(new_n759), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n707), .A2(G27), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G164), .B2(new_n707), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT96), .B(G2078), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT97), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n780), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n739), .A2(new_n767), .A3(new_n777), .A4(new_n784), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n721), .B(new_n723), .C1(KEYINPUT98), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n691), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n691), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1971), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G23), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT90), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G288), .B2(new_n691), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT32), .B(G1981), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n789), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT34), .ZN(new_n799));
  AND2_X1   g374(.A1(G290), .A2(KEYINPUT89), .ZN(new_n800));
  NOR2_X1   g375(.A1(G290), .A2(KEYINPUT89), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n800), .A2(new_n801), .A3(new_n691), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n691), .A2(G24), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n802), .A2(G1986), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(G1986), .B1(new_n802), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n477), .A2(G131), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n456), .A2(G107), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n472), .A2(KEYINPUT88), .A3(G119), .ZN(new_n809));
  AOI21_X1  g384(.A(KEYINPUT88), .B1(new_n472), .B2(G119), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n806), .B1(new_n807), .B2(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G25), .B(new_n811), .S(new_n707), .Z(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT35), .B(G1991), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n812), .B(new_n813), .Z(new_n814));
  NAND4_X1  g389(.A1(new_n799), .A2(new_n804), .A3(new_n805), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n785), .A2(KEYINPUT98), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n786), .A2(new_n817), .A3(new_n819), .A4(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  NAND2_X1  g397(.A1(new_n601), .A2(G559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT38), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n498), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n506), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n500), .A2(new_n827), .B1(new_n502), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n543), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n610), .B1(new_n826), .B2(new_n829), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n824), .B(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n830), .A2(new_n836), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(G145));
  XNOR2_X1  g417(.A(G162), .B(new_n623), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n811), .B(new_n629), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  INV_X1    g421(.A(G118), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(G2105), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n477), .A2(G142), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT102), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n848), .B(new_n850), .C1(G130), .C2(new_n472), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT103), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n486), .A2(KEYINPUT101), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n490), .A2(new_n492), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n481), .A2(new_n485), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n715), .B(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n860), .A2(new_n773), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n773), .ZN(new_n862));
  OR3_X1    g437(.A1(new_n861), .A2(new_n862), .A3(new_n735), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n735), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n852), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n854), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n865), .B1(new_n854), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n844), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n865), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n844), .B1(new_n872), .B2(new_n853), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g451(.A1(new_n601), .A2(G299), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT105), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n601), .A2(G299), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n879), .B(KEYINPUT104), .Z(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(KEYINPUT41), .A3(new_n878), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n878), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n831), .A2(new_n832), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n615), .B(new_n887), .ZN(new_n888));
  MUX2_X1   g463(.A(new_n885), .B(new_n886), .S(new_n888), .Z(new_n889));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n889), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G290), .B(G305), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n512), .B(G288), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n890), .B2(KEYINPUT42), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n893), .A2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(G868), .B2(new_n830), .ZN(G295));
  OAI21_X1  g476(.A(new_n900), .B1(G868), .B2(new_n830), .ZN(G331));
  INV_X1    g477(.A(new_n896), .ZN(new_n903));
  XNOR2_X1  g478(.A(G301), .B(G168), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n833), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n904), .A2(new_n833), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n833), .A3(KEYINPUT108), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n907), .A2(new_n886), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n882), .A2(new_n884), .B1(new_n908), .B2(new_n905), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(KEYINPUT109), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n908), .A2(new_n905), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n885), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n896), .B1(new_n918), .B2(new_n910), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n919), .B2(G37), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n896), .A3(new_n910), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n918), .A2(KEYINPUT110), .A3(new_n896), .A4(new_n910), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT43), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n925), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n886), .A2(new_n908), .A3(new_n905), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(KEYINPUT41), .B2(new_n886), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n933), .B2(new_n903), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n927), .B(KEYINPUT44), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n921), .B2(new_n928), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n926), .A2(new_n934), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n942));
  OAI21_X1  g517(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(G397));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  INV_X1    g519(.A(new_n492), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n491), .B1(new_n460), .B2(new_n488), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n858), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n460), .A2(new_n482), .B1(new_n949), .B2(new_n480), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(new_n857), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n944), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G125), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n467), .B2(new_n468), .ZN(new_n957));
  INV_X1    g532(.A(new_n464), .ZN(new_n958));
  OAI21_X1  g533(.A(G2105), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(new_n459), .A3(G40), .A4(new_n461), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n811), .A2(new_n813), .ZN(new_n962));
  INV_X1    g537(.A(G2067), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n715), .B(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n735), .B(new_n738), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n811), .A2(new_n813), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(G290), .B(G1986), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n960), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n950), .B1(new_n945), .B2(new_n946), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n944), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n972), .B2(new_n954), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT45), .B1(new_n859), .B2(new_n944), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n749), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n960), .B1(new_n972), .B2(KEYINPUT50), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n977));
  NAND3_X1  g552(.A1(new_n859), .A2(new_n944), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n746), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G8), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  NOR2_X1   g557(.A1(G168), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(KEYINPUT51), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT124), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n975), .A2(new_n979), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n975), .B2(new_n979), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n987), .A2(new_n988), .A3(G286), .ZN(new_n989));
  NAND2_X1  g564(.A1(KEYINPUT51), .A2(G8), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n970), .A2(new_n944), .A3(new_n859), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  OR2_X1    g573(.A1(G288), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n999), .A3(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT52), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT113), .B(G1981), .Z(new_n1006));
  NOR2_X1   g581(.A1(G305), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G305), .A2(G1981), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1012), .A2(new_n1013), .A3(KEYINPUT49), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1007), .ZN(new_n1015));
  AND3_X1   g590(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT114), .B1(G305), .B2(G1981), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT115), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n997), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1015), .B(KEYINPUT49), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT116), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1005), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT45), .B(new_n944), .C1(new_n947), .C2(new_n951), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n954), .B1(G164), .B2(G1384), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n970), .ZN(new_n1027));
  INV_X1    g602(.A(G1971), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n976), .A2(new_n978), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(G2090), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n560), .A2(G8), .A3(new_n561), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n560), .A2(KEYINPUT55), .A3(new_n561), .A4(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1031), .A2(new_n1036), .A3(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n970), .B1(new_n972), .B2(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n977), .B1(new_n859), .B2(new_n944), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  INV_X1    g616(.A(new_n977), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n952), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1384), .B1(new_n856), .B2(new_n950), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n960), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1040), .A2(new_n1041), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n982), .B1(new_n1049), .B2(new_n1029), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1037), .B1(new_n1050), .B2(new_n1036), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1024), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1027), .B2(G2078), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1030), .A2(new_n765), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n973), .A2(new_n974), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1053), .A2(G2078), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1054), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1052), .A2(G171), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n994), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1062));
  INV_X1    g637(.A(G1956), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT56), .B(G2072), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1025), .A2(new_n1026), .A3(new_n970), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n1068));
  XNOR2_X1  g643(.A(G299), .B(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1064), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1348), .B1(new_n976), .B2(new_n978), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n995), .A2(G2067), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n601), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1071), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n543), .A2(KEYINPUT120), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1025), .A2(new_n1026), .A3(new_n738), .A4(new_n970), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  NAND2_X1  g656(.A1(new_n995), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1077), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1069), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1072), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1348), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1030), .A2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n995), .A2(G2067), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n596), .A2(KEYINPUT123), .A3(new_n600), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT123), .B1(new_n596), .B2(new_n600), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n1093), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1073), .A2(new_n1074), .A3(new_n1098), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1095), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1097), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1086), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1103), .B(new_n1077), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1104));
  AND4_X1   g679(.A1(new_n1087), .A2(new_n1090), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1064), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1071), .A2(KEYINPUT61), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1071), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n1106), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1076), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G301), .B(KEYINPUT54), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1025), .A2(new_n970), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1057), .B(new_n1114), .C1(new_n952), .C2(new_n954), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1055), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1117), .A2(new_n1054), .B1(new_n1113), .B2(new_n1058), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n993), .A2(new_n1052), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1013), .B1(new_n1012), .B2(KEYINPUT49), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1018), .A2(KEYINPUT115), .A3(new_n1019), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n996), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1022), .B(new_n1124), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n1004), .B(new_n1037), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n1015), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1126), .B1(new_n1130), .B2(new_n997), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n981), .A2(G286), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT63), .B1(new_n1052), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1037), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1036), .B1(new_n1031), .B2(G8), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n980), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1004), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1131), .B(KEYINPUT118), .C1(new_n1133), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1036), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1143));
  AOI21_X1  g718(.A(G2090), .B1(new_n1062), .B2(KEYINPUT117), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1048), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1145), .B2(new_n982), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1138), .A2(new_n1037), .A3(new_n1146), .A4(new_n1132), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1147), .A2(new_n1148), .B1(new_n1138), .B2(new_n1137), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1007), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1150), .A2(new_n996), .B1(new_n1024), .B2(new_n1037), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1141), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1120), .B1(new_n1140), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1061), .B1(new_n1153), .B2(KEYINPUT125), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1155), .B(new_n1120), .C1(new_n1140), .C2(new_n1152), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n969), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n961), .ZN(new_n1158));
  INV_X1    g733(.A(new_n735), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n964), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT46), .B1(new_n1158), .B2(G1996), .ZN(new_n1161));
  OR3_X1    g736(.A1(new_n1158), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT47), .ZN(new_n1164));
  OR3_X1    g739(.A1(G290), .A2(new_n1158), .A3(G1986), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(KEYINPUT48), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1166), .A2(KEYINPUT48), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1167), .B(new_n1168), .C1(new_n961), .C2(new_n967), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n964), .A2(new_n965), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1170), .A2(new_n962), .B1(G2067), .B2(new_n715), .ZN(new_n1171));
  AOI211_X1 g746(.A(new_n1164), .B(new_n1169), .C1(new_n961), .C2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1157), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n663), .A2(new_n664), .A3(G319), .ZN(new_n1176));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n1177));
  XNOR2_X1  g751(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  INV_X1    g752(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n689), .A2(new_n646), .ZN(new_n1180));
  INV_X1    g754(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n1175), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g756(.A1(new_n1178), .A2(new_n1180), .A3(KEYINPUT127), .ZN(new_n1183));
  OAI21_X1  g757(.A(new_n875), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g758(.A1(new_n1184), .A2(new_n941), .ZN(G308));
  OAI221_X1 g759(.A(new_n875), .B1(new_n1182), .B2(new_n1183), .C1(new_n940), .C2(new_n938), .ZN(G225));
endmodule


