

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U552 ( .A(KEYINPUT1), .B(n560), .Z(n657) );
  NOR2_X2 U553 ( .A1(n769), .A2(n768), .ZN(n825) );
  BUF_X1 U554 ( .A(n689), .Z(n548) );
  NOR2_X2 U555 ( .A1(G2105), .A2(n528), .ZN(n895) );
  NOR2_X2 U556 ( .A1(n658), .A2(n559), .ZN(n650) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n701) );
  XNOR2_X1 U558 ( .A(n763), .B(KEYINPUT65), .ZN(n765) );
  XNOR2_X1 U559 ( .A(n524), .B(n523), .ZN(n689) );
  XNOR2_X1 U560 ( .A(n522), .B(KEYINPUT17), .ZN(n523) );
  NAND2_X1 U561 ( .A1(G101), .A2(n895), .ZN(n525) );
  AND2_X1 U562 ( .A1(n694), .A2(n693), .ZN(G164) );
  XNOR2_X1 U563 ( .A(KEYINPUT86), .B(n687), .ZN(n519) );
  XOR2_X1 U564 ( .A(n739), .B(KEYINPUT31), .Z(n520) );
  OR2_X1 U565 ( .A1(n729), .A2(n728), .ZN(n521) );
  INV_X1 U566 ( .A(G2104), .ZN(n528) );
  INV_X1 U567 ( .A(n708), .ZN(n724) );
  NOR2_X1 U568 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n740) );
  INV_X1 U570 ( .A(KEYINPUT105), .ZN(n741) );
  XNOR2_X1 U571 ( .A(n740), .B(KEYINPUT104), .ZN(n752) );
  INV_X1 U572 ( .A(n931), .ZN(n760) );
  NOR2_X1 U573 ( .A1(n833), .A2(n760), .ZN(n761) );
  AND2_X1 U574 ( .A1(n762), .A2(n761), .ZN(n763) );
  INV_X1 U575 ( .A(KEYINPUT33), .ZN(n764) );
  INV_X1 U576 ( .A(KEYINPUT66), .ZN(n522) );
  AND2_X1 U577 ( .A1(n765), .A2(n764), .ZN(n769) );
  XNOR2_X1 U578 ( .A(n596), .B(KEYINPUT15), .ZN(n597) );
  XOR2_X1 U579 ( .A(KEYINPUT74), .B(n597), .Z(n716) );
  NOR2_X1 U580 ( .A1(G651), .A2(n658), .ZN(n653) );
  NOR2_X2 U581 ( .A1(n529), .A2(G2104), .ZN(n900) );
  NOR2_X1 U582 ( .A1(n587), .A2(n586), .ZN(n923) );
  NOR2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  NAND2_X1 U584 ( .A1(G137), .A2(n689), .ZN(n527) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n525), .Z(n526) );
  NAND2_X1 U586 ( .A1(n527), .A2(n526), .ZN(n533) );
  INV_X1 U587 ( .A(G2105), .ZN(n529) );
  NOR2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n686) );
  NAND2_X1 U589 ( .A1(G113), .A2(n686), .ZN(n531) );
  NAND2_X1 U590 ( .A1(G125), .A2(n900), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X2 U592 ( .A1(n533), .A2(n532), .ZN(G160) );
  XOR2_X1 U593 ( .A(G2438), .B(G2454), .Z(n535) );
  XNOR2_X1 U594 ( .A(G2435), .B(G2430), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U596 ( .A(n536), .B(G2427), .Z(n538) );
  XNOR2_X1 U597 ( .A(G1348), .B(G1341), .ZN(n537) );
  XNOR2_X1 U598 ( .A(n538), .B(n537), .ZN(n542) );
  XOR2_X1 U599 ( .A(G2443), .B(G2446), .Z(n540) );
  XNOR2_X1 U600 ( .A(KEYINPUT108), .B(G2451), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U602 ( .A(n542), .B(n541), .Z(n543) );
  AND2_X1 U603 ( .A1(G14), .A2(n543), .ZN(G401) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U605 ( .A1(G123), .A2(n900), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n544), .B(KEYINPUT76), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n545), .B(KEYINPUT18), .ZN(n547) );
  NAND2_X1 U608 ( .A1(G99), .A2(n895), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n552) );
  BUF_X1 U610 ( .A(n686), .Z(n899) );
  NAND2_X1 U611 ( .A1(n899), .A2(G111), .ZN(n550) );
  NAND2_X1 U612 ( .A1(G135), .A2(n548), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n999) );
  XNOR2_X1 U615 ( .A(n999), .B(G2096), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n553), .B(KEYINPUT77), .ZN(n554) );
  OR2_X1 U617 ( .A1(G2100), .A2(n554), .ZN(G156) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  NOR2_X1 U621 ( .A1(G651), .A2(G543), .ZN(n646) );
  NAND2_X1 U622 ( .A1(n646), .A2(G90), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT69), .B(n555), .Z(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT0), .B(G543), .Z(n658) );
  INV_X1 U625 ( .A(G651), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n650), .A2(G77), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n558), .B(KEYINPUT9), .ZN(n562) );
  NOR2_X1 U629 ( .A1(G543), .A2(n559), .ZN(n560) );
  NAND2_X1 U630 ( .A1(G64), .A2(n657), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n653), .A2(G52), .ZN(n563) );
  XOR2_X1 U633 ( .A(KEYINPUT68), .B(n563), .Z(n564) );
  NOR2_X1 U634 ( .A1(n565), .A2(n564), .ZN(G171) );
  NAND2_X1 U635 ( .A1(G50), .A2(n653), .ZN(n566) );
  XNOR2_X1 U636 ( .A(n566), .B(KEYINPUT82), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G62), .A2(n657), .ZN(n567) );
  XOR2_X1 U638 ( .A(KEYINPUT81), .B(n567), .Z(n568) );
  NAND2_X1 U639 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G88), .A2(n646), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G75), .A2(n650), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U643 ( .A(KEYINPUT83), .B(n572), .Z(n573) );
  NOR2_X1 U644 ( .A1(n574), .A2(n573), .ZN(G166) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U646 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U647 ( .A(G223), .ZN(n844) );
  NAND2_X1 U648 ( .A1(n844), .A2(G567), .ZN(n576) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U650 ( .A1(n657), .A2(G56), .ZN(n577) );
  XNOR2_X1 U651 ( .A(n577), .B(KEYINPUT14), .ZN(n579) );
  NAND2_X1 U652 ( .A1(G43), .A2(n653), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n646), .A2(G81), .ZN(n580) );
  XOR2_X1 U655 ( .A(KEYINPUT12), .B(n580), .Z(n583) );
  NAND2_X1 U656 ( .A1(n650), .A2(G68), .ZN(n581) );
  XOR2_X1 U657 ( .A(n581), .B(KEYINPUT70), .Z(n582) );
  NOR2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U659 ( .A(KEYINPUT71), .B(n584), .Z(n585) );
  XNOR2_X1 U660 ( .A(n585), .B(KEYINPUT13), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n923), .A2(G860), .ZN(G153) );
  INV_X1 U662 ( .A(G171), .ZN(G301) );
  NAND2_X1 U663 ( .A1(G301), .A2(G868), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n588), .B(KEYINPUT72), .ZN(n599) );
  INV_X1 U665 ( .A(G868), .ZN(n669) );
  NAND2_X1 U666 ( .A1(G79), .A2(n650), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G92), .A2(n646), .ZN(n590) );
  NAND2_X1 U668 ( .A1(G54), .A2(n653), .ZN(n589) );
  NAND2_X1 U669 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U670 ( .A1(G66), .A2(n657), .ZN(n591) );
  XNOR2_X1 U671 ( .A(KEYINPUT73), .B(n591), .ZN(n592) );
  NOR2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U674 ( .A(n716), .ZN(n625) );
  INV_X1 U675 ( .A(n625), .ZN(n933) );
  NAND2_X1 U676 ( .A1(n669), .A2(n933), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U678 ( .A1(n646), .A2(G89), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n600), .B(KEYINPUT4), .ZN(n602) );
  NAND2_X1 U680 ( .A1(G76), .A2(n650), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U682 ( .A(KEYINPUT5), .B(n603), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n653), .A2(G51), .ZN(n604) );
  XOR2_X1 U684 ( .A(KEYINPUT75), .B(n604), .Z(n606) );
  NAND2_X1 U685 ( .A1(n657), .A2(G63), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U687 ( .A(KEYINPUT6), .B(n607), .Z(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U689 ( .A(KEYINPUT7), .B(n610), .ZN(G168) );
  XOR2_X1 U690 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U691 ( .A1(G65), .A2(n657), .ZN(n612) );
  NAND2_X1 U692 ( .A1(G53), .A2(n653), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G91), .A2(n646), .ZN(n614) );
  NAND2_X1 U695 ( .A1(G78), .A2(n650), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n930) );
  INV_X1 U698 ( .A(n930), .ZN(G299) );
  NOR2_X1 U699 ( .A1(G286), .A2(n669), .ZN(n618) );
  NOR2_X1 U700 ( .A1(G868), .A2(G299), .ZN(n617) );
  NOR2_X1 U701 ( .A1(n618), .A2(n617), .ZN(G297) );
  INV_X1 U702 ( .A(G860), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n619), .A2(G559), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n620), .A2(n625), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U706 ( .A1(G868), .A2(n625), .ZN(n622) );
  NOR2_X1 U707 ( .A1(G559), .A2(n622), .ZN(n624) );
  AND2_X1 U708 ( .A1(n669), .A2(n923), .ZN(n623) );
  NOR2_X1 U709 ( .A1(n624), .A2(n623), .ZN(G282) );
  XOR2_X1 U710 ( .A(n923), .B(KEYINPUT78), .Z(n627) );
  NAND2_X1 U711 ( .A1(G559), .A2(n625), .ZN(n626) );
  XNOR2_X1 U712 ( .A(n627), .B(n626), .ZN(n666) );
  NOR2_X1 U713 ( .A1(G860), .A2(n666), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G67), .A2(n657), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G55), .A2(n653), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G93), .A2(n646), .ZN(n631) );
  NAND2_X1 U718 ( .A1(G80), .A2(n650), .ZN(n630) );
  NAND2_X1 U719 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U720 ( .A(KEYINPUT79), .B(n632), .Z(n633) );
  OR2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n668) );
  XOR2_X1 U722 ( .A(n635), .B(n668), .Z(G145) );
  NAND2_X1 U723 ( .A1(G48), .A2(n653), .ZN(n642) );
  NAND2_X1 U724 ( .A1(G86), .A2(n646), .ZN(n637) );
  NAND2_X1 U725 ( .A1(G61), .A2(n657), .ZN(n636) );
  NAND2_X1 U726 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n650), .A2(G73), .ZN(n638) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n638), .Z(n639) );
  NOR2_X1 U729 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U731 ( .A(n643), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U732 ( .A1(G60), .A2(n657), .ZN(n645) );
  NAND2_X1 U733 ( .A1(G47), .A2(n653), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G85), .A2(n646), .ZN(n647) );
  XNOR2_X1 U736 ( .A(KEYINPUT67), .B(n647), .ZN(n648) );
  NOR2_X1 U737 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n650), .A2(G72), .ZN(n651) );
  NAND2_X1 U739 ( .A1(n652), .A2(n651), .ZN(G290) );
  NAND2_X1 U740 ( .A1(G49), .A2(n653), .ZN(n655) );
  NAND2_X1 U741 ( .A1(G74), .A2(G651), .ZN(n654) );
  NAND2_X1 U742 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U743 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n658), .A2(G87), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n660), .A2(n659), .ZN(G288) );
  XNOR2_X1 U746 ( .A(G305), .B(G166), .ZN(n665) );
  XOR2_X1 U747 ( .A(n668), .B(G290), .Z(n663) );
  XNOR2_X1 U748 ( .A(n930), .B(KEYINPUT19), .ZN(n661) );
  XNOR2_X1 U749 ( .A(n661), .B(G288), .ZN(n662) );
  XNOR2_X1 U750 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U751 ( .A(n665), .B(n664), .ZN(n911) );
  XNOR2_X1 U752 ( .A(n666), .B(n911), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n673), .ZN(n675) );
  XNOR2_X1 U759 ( .A(KEYINPUT84), .B(KEYINPUT21), .ZN(n674) );
  XNOR2_X1 U760 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G2072), .A2(n676), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n677) );
  XNOR2_X1 U764 ( .A(KEYINPUT22), .B(n677), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n678), .A2(G96), .ZN(n679) );
  NOR2_X1 U766 ( .A1(n679), .A2(G218), .ZN(n680) );
  XNOR2_X1 U767 ( .A(n680), .B(KEYINPUT85), .ZN(n848) );
  NAND2_X1 U768 ( .A1(n848), .A2(G2106), .ZN(n684) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n681) );
  NOR2_X1 U770 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U771 ( .A1(G108), .A2(n682), .ZN(n849) );
  NAND2_X1 U772 ( .A1(n849), .A2(G567), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n684), .A2(n683), .ZN(n850) );
  NAND2_X1 U774 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U775 ( .A1(n850), .A2(n685), .ZN(n847) );
  NAND2_X1 U776 ( .A1(n847), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  NAND2_X1 U778 ( .A1(G126), .A2(n900), .ZN(n688) );
  NAND2_X1 U779 ( .A1(G114), .A2(n686), .ZN(n687) );
  AND2_X1 U780 ( .A1(n688), .A2(n519), .ZN(n694) );
  NAND2_X1 U781 ( .A1(G138), .A2(n689), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n895), .A2(G102), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U784 ( .A(n692), .B(KEYINPUT87), .ZN(n693) );
  NOR2_X1 U785 ( .A1(G164), .A2(G1384), .ZN(n778) );
  NAND2_X1 U786 ( .A1(G160), .A2(G40), .ZN(n779) );
  INV_X1 U787 ( .A(n779), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n778), .A2(n695), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n696), .B(KEYINPUT64), .ZN(n708) );
  NAND2_X1 U790 ( .A1(n724), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U791 ( .A(KEYINPUT100), .B(KEYINPUT27), .ZN(n697) );
  XNOR2_X1 U792 ( .A(n698), .B(n697), .ZN(n700) );
  INV_X1 U793 ( .A(G1956), .ZN(n949) );
  NOR2_X1 U794 ( .A1(n724), .A2(n949), .ZN(n699) );
  NOR2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n703) );
  NOR2_X1 U796 ( .A1(n703), .A2(n930), .ZN(n702) );
  XNOR2_X1 U797 ( .A(n702), .B(n701), .ZN(n722) );
  NAND2_X1 U798 ( .A1(n703), .A2(n930), .ZN(n720) );
  XOR2_X1 U799 ( .A(KEYINPUT26), .B(KEYINPUT101), .Z(n705) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n724), .ZN(n704) );
  XNOR2_X1 U801 ( .A(n705), .B(n704), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n706), .A2(n923), .ZN(n714) );
  NAND2_X1 U803 ( .A1(G1341), .A2(n730), .ZN(n707) );
  XNOR2_X1 U804 ( .A(n707), .B(KEYINPUT102), .ZN(n712) );
  NAND2_X1 U805 ( .A1(G2067), .A2(n724), .ZN(n710) );
  BUF_X1 U806 ( .A(n708), .Z(n730) );
  NAND2_X1 U807 ( .A1(n730), .A2(G1348), .ZN(n709) );
  NAND2_X1 U808 ( .A1(n710), .A2(n709), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n711) );
  NAND2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U811 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U815 ( .A(n723), .B(KEYINPUT29), .ZN(n729) );
  NOR2_X1 U816 ( .A1(G1961), .A2(n724), .ZN(n725) );
  XOR2_X1 U817 ( .A(KEYINPUT99), .B(n725), .Z(n727) );
  XOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .Z(n981) );
  NOR2_X1 U819 ( .A1(n730), .A2(n981), .ZN(n726) );
  NOR2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n736) );
  NOR2_X1 U821 ( .A1(G301), .A2(n736), .ZN(n728) );
  NAND2_X1 U822 ( .A1(n708), .A2(G8), .ZN(n833) );
  NOR2_X1 U823 ( .A1(G1966), .A2(n833), .ZN(n754) );
  NOR2_X1 U824 ( .A1(n730), .A2(G2084), .ZN(n751) );
  NOR2_X1 U825 ( .A1(n754), .A2(n751), .ZN(n732) );
  INV_X1 U826 ( .A(KEYINPUT103), .ZN(n731) );
  XNOR2_X1 U827 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U828 ( .A1(n733), .A2(G8), .ZN(n734) );
  XNOR2_X1 U829 ( .A(n734), .B(KEYINPUT30), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n735), .A2(G168), .ZN(n738) );
  AND2_X1 U831 ( .A1(G301), .A2(n736), .ZN(n737) );
  NOR2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n752), .A2(G286), .ZN(n742) );
  XNOR2_X1 U834 ( .A(n742), .B(n741), .ZN(n748) );
  NOR2_X1 U835 ( .A1(n730), .A2(G2090), .ZN(n743) );
  XNOR2_X1 U836 ( .A(n743), .B(KEYINPUT106), .ZN(n745) );
  NOR2_X1 U837 ( .A1(n833), .A2(G1971), .ZN(n744) );
  NOR2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U839 ( .A1(G303), .A2(n746), .ZN(n747) );
  NAND2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U841 ( .A1(n749), .A2(G8), .ZN(n750) );
  XNOR2_X1 U842 ( .A(n750), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X1 U843 ( .A1(G8), .A2(n751), .ZN(n756) );
  INV_X1 U844 ( .A(n752), .ZN(n753) );
  NOR2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n829) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n759) );
  NOR2_X1 U850 ( .A1(n766), .A2(n759), .ZN(n924) );
  NAND2_X1 U851 ( .A1(n829), .A2(n924), .ZN(n762) );
  NAND2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n931) );
  NAND2_X1 U853 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n767), .A2(n833), .ZN(n768) );
  XOR2_X1 U855 ( .A(G305), .B(G1981), .Z(n926) );
  NAND2_X1 U856 ( .A1(G129), .A2(n900), .ZN(n776) );
  NAND2_X1 U857 ( .A1(n899), .A2(G117), .ZN(n771) );
  NAND2_X1 U858 ( .A1(G141), .A2(n548), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n895), .A2(G105), .ZN(n772) );
  XOR2_X1 U861 ( .A(KEYINPUT38), .B(n772), .Z(n773) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n777), .B(KEYINPUT94), .ZN(n878) );
  NOR2_X1 U865 ( .A1(G1996), .A2(n878), .ZN(n1005) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n780), .B(KEYINPUT88), .ZN(n819) );
  INV_X1 U868 ( .A(n819), .ZN(n791) );
  NAND2_X1 U869 ( .A1(G1996), .A2(n878), .ZN(n789) );
  NAND2_X1 U870 ( .A1(n900), .A2(G119), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G131), .A2(n548), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G107), .A2(n899), .ZN(n783) );
  XNOR2_X1 U874 ( .A(KEYINPUT93), .B(n783), .ZN(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n895), .A2(G95), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n888) );
  NAND2_X1 U878 ( .A1(G1991), .A2(n888), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U880 ( .A(KEYINPUT95), .B(n790), .ZN(n1011) );
  NOR2_X1 U881 ( .A1(n791), .A2(n1011), .ZN(n815) );
  NOR2_X1 U882 ( .A1(G1991), .A2(n888), .ZN(n1000) );
  NOR2_X1 U883 ( .A1(G1986), .A2(G290), .ZN(n792) );
  XOR2_X1 U884 ( .A(n792), .B(KEYINPUT107), .Z(n793) );
  NOR2_X1 U885 ( .A1(n1000), .A2(n793), .ZN(n794) );
  NOR2_X1 U886 ( .A1(n815), .A2(n794), .ZN(n795) );
  NOR2_X1 U887 ( .A1(n1005), .A2(n795), .ZN(n796) );
  XNOR2_X1 U888 ( .A(n796), .B(KEYINPUT39), .ZN(n810) );
  XNOR2_X1 U889 ( .A(KEYINPUT36), .B(KEYINPUT92), .ZN(n808) );
  NAND2_X1 U890 ( .A1(G116), .A2(n899), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G128), .A2(n900), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U893 ( .A(KEYINPUT35), .B(n799), .ZN(n806) );
  XNOR2_X1 U894 ( .A(KEYINPUT34), .B(KEYINPUT90), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n895), .A2(G104), .ZN(n802) );
  NAND2_X1 U896 ( .A1(G140), .A2(n548), .ZN(n800) );
  XOR2_X1 U897 ( .A(KEYINPUT89), .B(n800), .Z(n801) );
  NAND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U899 ( .A(n804), .B(n803), .Z(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U902 ( .A(KEYINPUT91), .B(n809), .ZN(n907) );
  XNOR2_X1 U903 ( .A(KEYINPUT37), .B(G2067), .ZN(n811) );
  NOR2_X1 U904 ( .A1(n907), .A2(n811), .ZN(n1021) );
  NAND2_X1 U905 ( .A1(n1021), .A2(n819), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n810), .A2(n814), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n907), .A2(n811), .ZN(n1018) );
  NAND2_X1 U908 ( .A1(n812), .A2(n1018), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n813), .A2(n819), .ZN(n837) );
  INV_X1 U910 ( .A(n837), .ZN(n823) );
  INV_X1 U911 ( .A(n814), .ZN(n817) );
  XNOR2_X1 U912 ( .A(KEYINPUT96), .B(n815), .ZN(n816) );
  NOR2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n818), .B(KEYINPUT97), .ZN(n821) );
  XNOR2_X1 U915 ( .A(G1986), .B(G290), .ZN(n939) );
  AND2_X1 U916 ( .A1(n939), .A2(n819), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  OR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n826) );
  AND2_X1 U919 ( .A1(n926), .A2(n826), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n842) );
  INV_X1 U921 ( .A(n826), .ZN(n840) );
  NOR2_X1 U922 ( .A1(G2090), .A2(G303), .ZN(n827) );
  NAND2_X1 U923 ( .A1(G8), .A2(n827), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  AND2_X1 U925 ( .A1(n830), .A2(n833), .ZN(n836) );
  NOR2_X1 U926 ( .A1(G305), .A2(G1981), .ZN(n831) );
  XOR2_X1 U927 ( .A(n831), .B(KEYINPUT24), .Z(n832) );
  NOR2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n834), .B(KEYINPUT98), .ZN(n835) );
  NOR2_X1 U930 ( .A1(n836), .A2(n835), .ZN(n838) );
  AND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(n839) );
  OR2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U933 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U934 ( .A(n843), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U937 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U939 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  INV_X1 U946 ( .A(n850), .ZN(G319) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n852) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U950 ( .A(KEYINPUT109), .B(G2090), .Z(n854) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U954 ( .A(G2096), .B(G2100), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n860) );
  XOR2_X1 U956 ( .A(G2078), .B(G2084), .Z(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U958 ( .A(G1956), .B(G1966), .Z(n862) );
  XNOR2_X1 U959 ( .A(G1981), .B(G1976), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(n863), .B(G2474), .Z(n865) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U964 ( .A(KEYINPUT41), .B(G1961), .Z(n867) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1971), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U968 ( .A1(G100), .A2(n895), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G112), .A2(n899), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n872), .B(KEYINPUT111), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G136), .A2(n548), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n900), .A2(G124), .ZN(n875) );
  XOR2_X1 U975 ( .A(KEYINPUT44), .B(n875), .Z(n876) );
  NOR2_X1 U976 ( .A1(n877), .A2(n876), .ZN(G162) );
  XNOR2_X1 U977 ( .A(n878), .B(G162), .ZN(n887) );
  NAND2_X1 U978 ( .A1(G118), .A2(n899), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G130), .A2(n900), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U981 ( .A1(n895), .A2(G106), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G142), .A2(n548), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n892) );
  XNOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n888), .B(KEYINPUT112), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U990 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U991 ( .A(G160), .B(n999), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n906) );
  NAND2_X1 U993 ( .A1(n895), .A2(G103), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G139), .A2(n548), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(KEYINPUT113), .B(n898), .Z(n905) );
  NAND2_X1 U997 ( .A1(G115), .A2(n899), .ZN(n902) );
  NAND2_X1 U998 ( .A1(G127), .A2(n900), .ZN(n901) );
  NAND2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n903), .Z(n904) );
  NOR2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(n1012) );
  XOR2_X1 U1002 ( .A(n906), .B(n1012), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G164), .B(n907), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n910), .ZN(G395) );
  XOR2_X1 U1006 ( .A(n911), .B(G286), .Z(n913) );
  XNOR2_X1 U1007 ( .A(G171), .B(n933), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n914), .B(n923), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n915), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(KEYINPUT114), .B(n916), .ZN(G397) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n917), .B(KEYINPUT49), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n918), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(KEYINPUT115), .B(n920), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1021 ( .A(KEYINPUT56), .B(G16), .ZN(n947) );
  XNOR2_X1 U1022 ( .A(n923), .B(G1341), .ZN(n945) );
  XNOR2_X1 U1023 ( .A(G171), .B(G1961), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n943) );
  XNOR2_X1 U1025 ( .A(G1966), .B(G168), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(n928), .B(KEYINPUT57), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(KEYINPUT122), .B(n929), .ZN(n941) );
  XNOR2_X1 U1029 ( .A(G1956), .B(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(G1348), .B(n933), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(G1971), .A2(G303), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n1031) );
  XNOR2_X1 U1040 ( .A(KEYINPUT123), .B(G1961), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(n948), .B(G5), .ZN(n964) );
  XNOR2_X1 U1042 ( .A(G1966), .B(G21), .ZN(n962) );
  XNOR2_X1 U1043 ( .A(n949), .B(G20), .ZN(n958) );
  XOR2_X1 U1044 ( .A(G1341), .B(G19), .Z(n953) );
  XOR2_X1 U1045 ( .A(G1348), .B(KEYINPUT125), .Z(n950) );
  XNOR2_X1 U1046 ( .A(G4), .B(n950), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n951), .B(KEYINPUT59), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT124), .B(G1981), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G6), .B(n954), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(n959), .B(KEYINPUT60), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT126), .B(n960), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n972) );
  XNOR2_X1 U1057 ( .A(G1986), .B(G24), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G23), .B(G1976), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(G1971), .B(KEYINPUT127), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(n967), .B(G22), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT58), .B(n970), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(KEYINPUT61), .B(n973), .ZN(n975) );
  INV_X1 U1066 ( .A(G16), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n976), .A2(G11), .ZN(n1029) );
  XNOR2_X1 U1069 ( .A(G2090), .B(G35), .ZN(n991) );
  XOR2_X1 U1070 ( .A(G1991), .B(G25), .Z(n977) );
  NAND2_X1 U1071 ( .A1(n977), .A2(G28), .ZN(n987) );
  XNOR2_X1 U1072 ( .A(G2067), .B(G26), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G2072), .B(G33), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT118), .B(n980), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G1996), .B(G32), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(G27), .B(n981), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1081 ( .A(KEYINPUT119), .B(n988), .Z(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(KEYINPUT53), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(n992), .B(KEYINPUT120), .ZN(n995) );
  XOR2_X1 U1085 ( .A(G2084), .B(G34), .Z(n993) );
  XNOR2_X1 U1086 ( .A(KEYINPUT54), .B(n993), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT55), .B(n996), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(G29), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(n998), .B(KEYINPUT121), .ZN(n1027) );
  XNOR2_X1 U1091 ( .A(G160), .B(G2084), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n1007) );
  XOR2_X1 U1095 ( .A(G2090), .B(G162), .Z(n1003) );
  XNOR2_X1 U1096 ( .A(KEYINPUT116), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(n1007), .B(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(G2072), .B(n1012), .Z(n1014) );
  XOR2_X1 U1102 ( .A(G164), .B(G2078), .Z(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(KEYINPUT50), .B(n1015), .Z(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(n1022), .B(KEYINPUT52), .ZN(n1024) );
  INV_X1 U1109 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

