//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  AOI21_X1  g000(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT97), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT102), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n208), .B(KEYINPUT89), .Z(new_n209));
  NOR2_X1   g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(KEYINPUT15), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n212), .B(KEYINPUT90), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n209), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n215), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT91), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(KEYINPUT92), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n220), .A2(new_n225), .ZN(new_n231));
  NOR2_X1   g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G99gat), .ZN(new_n236));
  INV_X1    g035(.A(G106gat), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT8), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n235), .B(new_n238), .C1(new_n233), .C2(new_n234), .ZN(new_n239));
  XOR2_X1   g038(.A(G99gat), .B(G106gat), .Z(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n230), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(KEYINPUT99), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT99), .B1(new_n246), .B2(new_n247), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G190gat), .B(G218gat), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT100), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n242), .B1(new_n226), .B2(new_n229), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n247), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT99), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n254), .B1(new_n257), .B2(new_n248), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT100), .ZN(new_n259));
  INV_X1    g058(.A(new_n252), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n207), .B1(new_n253), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT101), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n258), .B2(new_n260), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n251), .A2(KEYINPUT101), .A3(new_n252), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n206), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT102), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n270), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n262), .A2(new_n272), .A3(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT16), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(G1gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(G1gat), .B2(new_n275), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n278), .B(G8gat), .Z(new_n279));
  INV_X1    g078(.A(KEYINPUT21), .ZN(new_n280));
  XNOR2_X1  g079(.A(G57gat), .B(G64gat), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G71gat), .B(G78gat), .Z(new_n284));
  OR2_X1    g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n284), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n279), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(G231gat), .A2(G233gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT96), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  XNOR2_X1  g092(.A(new_n289), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n280), .ZN(new_n295));
  XOR2_X1   g094(.A(G127gat), .B(G155gat), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G211gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n299), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n287), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n245), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n241), .A2(new_n287), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n245), .A2(new_n303), .A3(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G230gat), .A2(G233gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT103), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT103), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n313), .A3(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n304), .A2(new_n306), .ZN(new_n317));
  INV_X1    g116(.A(new_n310), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G120gat), .B(G148gat), .ZN(new_n320));
  INV_X1    g119(.A(G176gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(G204gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n316), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n323), .B1(new_n311), .B2(new_n319), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n274), .A2(new_n302), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT95), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n228), .A2(new_n279), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n231), .A2(new_n279), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n230), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G229gat), .A2(G233gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(KEYINPUT18), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT94), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n228), .B2(new_n279), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(new_n332), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n335), .B(KEYINPUT13), .Z(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n335), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT18), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT93), .ZN(new_n346));
  XNOR2_X1  g145(.A(G113gat), .B(G141gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT11), .ZN(new_n348));
  INV_X1    g147(.A(G169gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G197gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT88), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT12), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n342), .B(new_n345), .C1(new_n346), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n336), .A2(new_n346), .A3(new_n341), .ZN(new_n356));
  INV_X1    g155(.A(new_n354), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n341), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT18), .B1(new_n334), .B2(new_n335), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363));
  AND2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G141gat), .B(G148gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(G155gat), .B2(G162gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n366), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G141gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(G148gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G141gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G155gat), .B(G162gat), .ZN(new_n376));
  INV_X1    g175(.A(G155gat), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT2), .B1(new_n377), .B2(new_n205), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G120gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G113gat), .ZN(new_n382));
  INV_X1    g181(.A(G113gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G120gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G127gat), .B(G134gat), .Z(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(KEYINPUT67), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n381), .A3(G113gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT68), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n383), .ZN(new_n395));
  NAND2_X1  g194(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(G120gat), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT69), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n395), .A2(KEYINPUT69), .A3(G120gat), .A4(new_n396), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n393), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n388), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n380), .B(new_n389), .C1(new_n401), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n393), .ZN(new_n406));
  AND2_X1   g205(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT69), .B1(new_n409), .B2(G120gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n400), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n412), .A2(new_n403), .B1(new_n387), .B2(new_n388), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n376), .B1(new_n378), .B2(new_n375), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT3), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n370), .A2(new_n379), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI22_X1  g218(.A1(new_n363), .A2(new_n405), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n389), .B1(new_n401), .B2(new_n404), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT71), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT71), .B(new_n389), .C1(new_n401), .C2(new_n404), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n380), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n420), .B1(new_n363), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(KEYINPUT5), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n423), .A2(KEYINPUT4), .A3(new_n380), .A4(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n370), .A2(new_n379), .A3(new_n417), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n417), .B1(new_n370), .B2(new_n379), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n405), .A2(new_n431), .B1(new_n434), .B2(new_n421), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT5), .ZN(new_n437));
  INV_X1    g236(.A(new_n380), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n405), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n440), .B2(new_n428), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n426), .A2(new_n429), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n443));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G57gat), .B(G85gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT80), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n436), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n425), .A2(new_n363), .ZN(new_n450));
  INV_X1    g249(.A(new_n420), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n429), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  INV_X1    g253(.A(new_n447), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n449), .A2(new_n452), .A3(new_n447), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT79), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n460), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT79), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n457), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n457), .A2(new_n463), .A3(new_n466), .A4(new_n461), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n453), .A2(new_n455), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(new_n460), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G8gat), .B(G36gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G64gat), .ZN(new_n473));
  INV_X1    g272(.A(G92gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT76), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  XNOR2_X1  g279(.A(G197gat), .B(G204gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G211gat), .B(G218gat), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n479), .A2(new_n483), .A3(new_n480), .A4(new_n481), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G226gat), .ZN(new_n488));
  INV_X1    g287(.A(G233gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G183gat), .A2(G190gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT24), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT24), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(G183gat), .A3(G190gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(G183gat), .A2(G190gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(G169gat), .A2(G176gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(G169gat), .A2(G176gat), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(KEYINPUT23), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT64), .ZN(new_n505));
  OAI22_X1  g304(.A1(new_n496), .A2(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n349), .A2(new_n321), .A3(KEYINPUT23), .ZN(new_n507));
  NAND2_X1  g306(.A1(G169gat), .A2(G176gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI22_X1  g308(.A1(new_n509), .A2(KEYINPUT64), .B1(KEYINPUT23), .B2(new_n503), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT25), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT26), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n508), .B1(new_n503), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n491), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G183gat), .ZN(new_n517));
  INV_X1    g316(.A(G190gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT28), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G183gat), .ZN(new_n522));
  AOI21_X1  g321(.A(G190gat), .B1(new_n522), .B2(KEYINPUT27), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT27), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n524), .A3(G183gat), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT28), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n516), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n528));
  INV_X1    g327(.A(new_n503), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT23), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n504), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n497), .B1(new_n492), .B2(new_n494), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n511), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT29), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n490), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n490), .ZN(new_n539));
  INV_X1    g338(.A(new_n500), .ZN(new_n540));
  NOR3_X1   g339(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n542), .A2(new_n495), .B1(new_n509), .B2(KEYINPUT64), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n504), .A2(new_n505), .B1(new_n530), .B2(new_n529), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n534), .B1(new_n545), .B2(KEYINPUT25), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n539), .B1(new_n546), .B2(new_n527), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n487), .B1(new_n538), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n536), .A2(new_n490), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n485), .A2(new_n486), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT29), .B1(new_n546), .B2(new_n527), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n490), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n548), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n547), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(KEYINPUT77), .A3(new_n550), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n476), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT30), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n554), .A2(new_n556), .A3(new_n476), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n557), .B2(KEYINPUT30), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n471), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G228gat), .A2(G233gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n550), .A2(new_n537), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n380), .B1(new_n565), .B2(new_n417), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n418), .A2(new_n537), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n487), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n564), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT82), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT3), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n571), .B(KEYINPUT29), .C1(new_n485), .C2(new_n486), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n380), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n567), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT83), .B1(new_n576), .B2(new_n550), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT83), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n487), .A2(new_n578), .A3(new_n567), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n577), .A2(new_n579), .A3(G228gat), .A4(G233gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n570), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT84), .B1(new_n581), .B2(G22gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(G78gat), .B(G106gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT31), .B(G50gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n581), .A2(G22gat), .ZN(new_n587));
  INV_X1    g386(.A(G22gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT29), .B1(new_n485), .B2(new_n486), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n417), .B1(new_n589), .B2(KEYINPUT82), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n438), .B1(new_n590), .B2(new_n573), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n564), .B1(new_n568), .B2(KEYINPUT83), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n579), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n588), .B1(new_n593), .B2(new_n570), .ZN(new_n594));
  OAI22_X1  g393(.A1(new_n582), .A2(new_n586), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n588), .A3(new_n570), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n596), .A2(KEYINPUT84), .A3(new_n597), .A4(new_n585), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n563), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n528), .B1(new_n543), .B2(new_n544), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n522), .A2(KEYINPUT27), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n525), .A3(new_n518), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT28), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n515), .B1(new_n605), .B2(new_n519), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n601), .A2(new_n606), .A3(new_n534), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n412), .A2(new_n403), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT71), .B1(new_n608), .B2(new_n389), .ZN(new_n609));
  INV_X1    g408(.A(new_n424), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(G227gat), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(new_n489), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n536), .A2(new_n423), .A3(new_n424), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT32), .ZN(new_n616));
  XNOR2_X1  g415(.A(G15gat), .B(G43gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G71gat), .B(G99gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n620), .B2(KEYINPUT33), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT72), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n616), .A2(KEYINPUT33), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n625), .B2(new_n620), .ZN(new_n626));
  AOI211_X1 g425(.A(KEYINPUT72), .B(new_n619), .C1(new_n615), .C2(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n613), .B1(new_n611), .B2(new_n614), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI211_X1 g431(.A(new_n613), .B(new_n630), .C1(new_n611), .C2(new_n614), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT74), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n634), .B(new_n622), .C1(new_n626), .C2(new_n627), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n639), .A2(KEYINPUT36), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n628), .A2(KEYINPUT74), .A3(new_n635), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT75), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n638), .A2(new_n640), .A3(KEYINPUT75), .A4(new_n641), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n636), .A2(new_n639), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT85), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n427), .B1(new_n450), .B2(new_n451), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT39), .B1(new_n440), .B2(new_n428), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n447), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n651), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n652), .A2(new_n656), .ZN(new_n659));
  INV_X1    g458(.A(new_n651), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n447), .A3(new_n660), .A4(new_n654), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n658), .A2(new_n661), .A3(new_n468), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n557), .A2(KEYINPUT30), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n558), .A3(new_n560), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n599), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n554), .A2(new_n556), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n476), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT37), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT38), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n442), .A2(new_n447), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n462), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n469), .ZN(new_n675));
  INV_X1    g474(.A(new_n557), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n475), .A2(KEYINPUT38), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT86), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n548), .A2(new_n552), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(KEYINPUT37), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT86), .B(new_n670), .C1(new_n548), .C2(new_n552), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n668), .B(new_n677), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n672), .A2(new_n675), .A3(new_n676), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n600), .A2(new_n649), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n628), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n686), .A2(new_n634), .B1(new_n595), .B2(new_n598), .ZN(new_n687));
  AND4_X1   g486(.A1(new_n638), .A2(new_n687), .A3(new_n641), .A4(new_n562), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT35), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n469), .B1(new_n464), .B2(KEYINPUT81), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(new_n467), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n636), .A2(new_n639), .ZN(new_n692));
  INV_X1    g491(.A(new_n675), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n595), .A2(new_n598), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n692), .A2(new_n562), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n688), .A2(new_n691), .B1(new_n695), .B2(new_n689), .ZN(new_n696));
  AOI211_X1 g495(.A(new_n331), .B(new_n362), .C1(new_n685), .C2(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n664), .B1(new_n690), .B2(new_n467), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n684), .B1(new_n699), .B2(new_n694), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n696), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT95), .B1(new_n701), .B2(new_n361), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n330), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n705), .B(new_n330), .C1(new_n697), .C2(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n471), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G1gat), .ZN(G1324gat));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT16), .B(G8gat), .Z(new_n712));
  NAND4_X1  g511(.A1(new_n562), .A2(new_n636), .A3(new_n639), .A4(new_n694), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n689), .B1(new_n713), .B2(new_n675), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n471), .A2(KEYINPUT35), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n687), .A2(new_n638), .A3(new_n641), .A4(new_n562), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n563), .A2(new_n599), .B1(new_n683), .B2(new_n665), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n649), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n331), .B1(new_n719), .B2(new_n362), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n701), .A2(KEYINPUT95), .A3(new_n361), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n705), .B1(new_n722), .B2(new_n330), .ZN(new_n723));
  AOI211_X1 g522(.A(KEYINPUT104), .B(new_n329), .C1(new_n720), .C2(new_n721), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n664), .B(new_n712), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n664), .B1(new_n723), .B2(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G8gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n664), .A2(KEYINPUT42), .A3(new_n712), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n707), .B2(new_n733), .ZN(new_n734));
  AOI211_X1 g533(.A(KEYINPUT105), .B(new_n732), .C1(new_n704), .C2(new_n706), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n711), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n725), .A2(new_n726), .B1(new_n728), .B2(G8gat), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n738), .B(KEYINPUT106), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1325gat));
  INV_X1    g539(.A(new_n707), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n741), .A2(G15gat), .A3(new_n646), .ZN(new_n742));
  OAI21_X1  g541(.A(G15gat), .B1(new_n741), .B2(new_n649), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1326gat));
  NAND2_X1  g543(.A1(new_n707), .A2(new_n599), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT43), .B(G22gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1327gat));
  AND3_X1   g546(.A1(new_n262), .A2(new_n272), .A3(new_n266), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n272), .B1(new_n262), .B2(new_n266), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n327), .A2(new_n302), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n722), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n753), .A2(G29gat), .A3(new_n471), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT45), .Z(new_n755));
  NOR2_X1   g554(.A1(new_n719), .A2(new_n274), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n759));
  NOR3_X1   g558(.A1(new_n719), .A2(new_n274), .A3(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n361), .A2(new_n751), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G29gat), .B1(new_n763), .B2(new_n471), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n755), .A2(new_n764), .ZN(G1328gat));
  OAI21_X1  g564(.A(G36gat), .B1(new_n763), .B2(new_n562), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n562), .A2(G36gat), .ZN(new_n767));
  OR3_X1    g566(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT46), .B1(new_n753), .B2(new_n767), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT108), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n766), .A2(new_n768), .A3(new_n772), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1329gat));
  NAND3_X1  g573(.A1(new_n761), .A2(new_n698), .A3(new_n762), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G43gat), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n753), .A2(G43gat), .A3(new_n646), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT109), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780));
  AOI211_X1 g579(.A(KEYINPUT109), .B(new_n780), .C1(new_n776), .C2(new_n777), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n779), .A2(new_n781), .ZN(G1330gat));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n753), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n722), .A2(KEYINPUT110), .A3(new_n752), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n694), .A2(G50gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT48), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n599), .B(new_n762), .C1(new_n758), .C2(new_n760), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(G50gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT112), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(G50gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n787), .A2(KEYINPUT111), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n788), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n792), .A2(new_n797), .ZN(G1331gat));
  NAND4_X1  g597(.A1(new_n274), .A2(new_n362), .A3(new_n302), .A4(new_n327), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n719), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n708), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g601(.A(new_n562), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT113), .Z(new_n805));
  NOR2_X1   g604(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1333gat));
  NAND2_X1  g606(.A1(new_n800), .A2(new_n698), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n646), .A2(G71gat), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n808), .A2(G71gat), .B1(new_n800), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g610(.A1(new_n800), .A2(new_n599), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g612(.A1(new_n361), .A2(new_n302), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n761), .A2(new_n327), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G85gat), .B1(new_n815), .B2(new_n471), .ZN(new_n816));
  INV_X1    g615(.A(new_n814), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n756), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n820), .B(new_n756), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n327), .A3(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n471), .A2(G85gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n816), .B1(new_n824), .B2(new_n825), .ZN(G1336gat));
  OAI21_X1  g625(.A(G92gat), .B1(new_n815), .B2(new_n562), .ZN(new_n827));
  INV_X1    g626(.A(new_n824), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n474), .A3(new_n664), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(KEYINPUT115), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT52), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n827), .B(new_n829), .C1(KEYINPUT115), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1337gat));
  AOI21_X1  g634(.A(G99gat), .B1(new_n828), .B2(new_n692), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n758), .A2(new_n760), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n328), .A3(new_n817), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n649), .A2(new_n236), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(G1338gat));
  OR2_X1    g639(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n841));
  NAND2_X1  g640(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n842));
  XNOR2_X1  g641(.A(KEYINPUT116), .B(G106gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(new_n838), .B2(new_n599), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n824), .A2(G106gat), .A3(new_n694), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n841), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n843), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n815), .B2(new_n694), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n237), .A3(new_n599), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT117), .A4(KEYINPUT53), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n846), .A2(new_n850), .ZN(G1339gat));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  INV_X1    g651(.A(new_n309), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n318), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n312), .A3(new_n314), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n311), .A2(KEYINPUT54), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n323), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n857), .A3(KEYINPUT55), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n324), .A2(new_n858), .A3(KEYINPUT118), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT118), .B1(new_n324), .B2(new_n858), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n855), .A2(new_n857), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n860), .A2(new_n861), .B1(KEYINPUT55), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n355), .B2(new_n360), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n334), .A2(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n865));
  INV_X1    g664(.A(new_n352), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n345), .A2(new_n341), .A3(new_n336), .A4(new_n354), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n327), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n274), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n863), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n868), .A2(new_n867), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n750), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n302), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n329), .A2(new_n361), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n471), .ZN(new_n878));
  INV_X1    g677(.A(new_n713), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G113gat), .B1(new_n880), .B2(new_n362), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n688), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n361), .A2(new_n409), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(G1340gat));
  NAND3_X1  g683(.A1(new_n878), .A2(new_n879), .A3(new_n327), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(G120gat), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n885), .B2(G120gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n327), .A2(new_n381), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT120), .Z(new_n891));
  OAI22_X1  g690(.A1(new_n888), .A2(new_n889), .B1(new_n882), .B2(new_n891), .ZN(G1341gat));
  INV_X1    g691(.A(new_n302), .ZN(new_n893));
  OAI21_X1  g692(.A(G127gat), .B1(new_n880), .B2(new_n893), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n893), .A2(G127gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n882), .B2(new_n895), .ZN(G1342gat));
  OR2_X1    g695(.A1(new_n274), .A2(G134gat), .ZN(new_n897));
  OR3_X1    g696(.A1(new_n882), .A2(KEYINPUT56), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n880), .B2(new_n274), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT56), .B1(new_n882), .B2(new_n897), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G1343gat));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n862), .A2(KEYINPUT55), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n324), .A2(new_n858), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n361), .A2(new_n905), .B1(new_n869), .B2(KEYINPUT121), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n750), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND4_X1   g707(.A1(new_n271), .A2(new_n872), .A3(new_n273), .A4(new_n873), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n893), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n330), .A2(new_n362), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n902), .B1(new_n912), .B2(new_n599), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n902), .B(new_n599), .C1(new_n875), .C2(new_n876), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n698), .A2(new_n471), .A3(new_n664), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n371), .B1(new_n917), .B2(new_n361), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n599), .B(new_n915), .C1(new_n875), .C2(new_n876), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n362), .A2(G141gat), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT58), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n872), .A2(new_n361), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n750), .B1(new_n924), .B2(new_n869), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n893), .B1(new_n925), .B2(new_n909), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n694), .B1(new_n926), .B2(new_n911), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n927), .A2(KEYINPUT122), .A3(new_n915), .A4(new_n920), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n929), .B1(new_n919), .B2(new_n921), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT58), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n694), .B1(new_n910), .B2(new_n911), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n914), .B(new_n915), .C1(new_n933), .C2(new_n902), .ZN(new_n934));
  OAI21_X1  g733(.A(G141gat), .B1(new_n934), .B2(new_n362), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n932), .A2(new_n935), .A3(KEYINPUT123), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT123), .B1(new_n932), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n923), .B1(new_n936), .B2(new_n937), .ZN(G1344gat));
  NOR3_X1   g737(.A1(new_n919), .A2(G148gat), .A3(new_n328), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT124), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT59), .B(new_n373), .C1(new_n917), .C2(new_n327), .ZN(new_n941));
  XOR2_X1   g740(.A(KEYINPUT125), .B(KEYINPUT59), .Z(new_n942));
  NAND2_X1  g741(.A1(new_n933), .A2(new_n902), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT57), .B1(new_n877), .B2(new_n694), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n943), .A2(new_n944), .A3(new_n327), .A4(new_n915), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n942), .B1(new_n945), .B2(G148gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n940), .B1(new_n941), .B2(new_n946), .ZN(G1345gat));
  OAI21_X1  g746(.A(G155gat), .B1(new_n934), .B2(new_n893), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n302), .A2(new_n377), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n919), .B2(new_n949), .ZN(G1346gat));
  OAI21_X1  g749(.A(G162gat), .B1(new_n934), .B2(new_n274), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n750), .A2(new_n205), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT126), .B1(new_n919), .B2(new_n952), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n919), .A2(KEYINPUT126), .A3(new_n952), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(G1347gat));
  NAND2_X1  g754(.A1(new_n926), .A2(new_n911), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n646), .A2(new_n599), .A3(new_n562), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n471), .A3(new_n957), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n958), .A2(new_n349), .A3(new_n362), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n877), .B2(new_n708), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n956), .A2(KEYINPUT127), .A3(new_n471), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n687), .A2(new_n638), .A3(new_n641), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n961), .A2(new_n962), .A3(new_n664), .A4(new_n963), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n964), .A2(new_n362), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n959), .B1(new_n965), .B2(new_n349), .ZN(G1348gat));
  OAI21_X1  g765(.A(G176gat), .B1(new_n958), .B2(new_n328), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n327), .A2(new_n321), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n964), .B2(new_n968), .ZN(G1349gat));
  OAI21_X1  g768(.A(G183gat), .B1(new_n958), .B2(new_n893), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n302), .A2(new_n517), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n964), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g772(.A(G190gat), .B1(new_n958), .B2(new_n274), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT61), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n974), .A2(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n750), .A2(new_n518), .ZN(new_n978));
  OAI22_X1  g777(.A1(new_n976), .A2(new_n977), .B1(new_n964), .B2(new_n978), .ZN(G1351gat));
  AND2_X1   g778(.A1(new_n943), .A2(new_n944), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n698), .A2(new_n708), .A3(new_n562), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(G197gat), .B1(new_n982), .B2(new_n362), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n698), .A2(new_n694), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n961), .A2(new_n962), .A3(new_n664), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n361), .A2(new_n351), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  NAND3_X1  g786(.A1(new_n980), .A2(new_n327), .A3(new_n981), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G204gat), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n328), .A2(G204gat), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  OR3_X1    g790(.A1(new_n985), .A2(KEYINPUT62), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(KEYINPUT62), .B1(new_n985), .B2(new_n991), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n989), .A2(new_n992), .A3(new_n993), .ZN(G1353gat));
  NAND4_X1  g793(.A1(new_n943), .A2(new_n944), .A3(new_n302), .A4(new_n981), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n302), .A2(new_n298), .ZN(new_n998));
  OAI22_X1  g797(.A1(new_n996), .A2(new_n997), .B1(new_n985), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n982), .B2(new_n274), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n274), .A2(G218gat), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n985), .B2(new_n1001), .ZN(G1355gat));
endmodule


