

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597;

  XNOR2_X1 U327 ( .A(KEYINPUT27), .B(KEYINPUT89), .ZN(n461) );
  NOR2_X1 U328 ( .A1(n473), .A2(n472), .ZN(n484) );
  XNOR2_X1 U329 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U330 ( .A(G50GAT), .B(n500), .Z(n295) );
  INV_X1 U331 ( .A(KEYINPUT9), .ZN(n388) );
  INV_X1 U332 ( .A(KEYINPUT81), .ZN(n336) );
  XNOR2_X1 U333 ( .A(KEYINPUT54), .B(KEYINPUT116), .ZN(n423) );
  XNOR2_X1 U334 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U335 ( .A(n524), .B(n461), .ZN(n468) );
  XNOR2_X1 U336 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U337 ( .A(n424), .B(n423), .ZN(n448) );
  INV_X1 U338 ( .A(KEYINPUT117), .ZN(n449) );
  XNOR2_X1 U339 ( .A(n339), .B(n338), .ZN(n412) );
  XNOR2_X1 U340 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  XNOR2_X1 U341 ( .A(n417), .B(KEYINPUT88), .ZN(n418) );
  XNOR2_X1 U342 ( .A(n572), .B(KEYINPUT36), .ZN(n593) );
  XNOR2_X1 U343 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U344 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U345 ( .A(n400), .B(n399), .ZN(n572) );
  XNOR2_X1 U346 ( .A(KEYINPUT120), .B(G183GAT), .ZN(n453) );
  XNOR2_X1 U347 ( .A(n454), .B(n453), .ZN(G1350GAT) );
  XOR2_X1 U348 ( .A(G155GAT), .B(G127GAT), .Z(n297) );
  XNOR2_X1 U349 ( .A(G15GAT), .B(G22GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U351 ( .A(KEYINPUT13), .B(G57GAT), .Z(n299) );
  XNOR2_X1 U352 ( .A(G211GAT), .B(G78GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n311) );
  XOR2_X1 U355 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n303) );
  XNOR2_X1 U356 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U358 ( .A(KEYINPUT76), .B(G71GAT), .Z(n305) );
  XOR2_X1 U359 ( .A(G1GAT), .B(G8GAT), .Z(n356) );
  XNOR2_X1 U360 ( .A(n356), .B(G183GAT), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U362 ( .A(n307), .B(n306), .Z(n309) );
  NAND2_X1 U363 ( .A1(G231GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U365 ( .A(n311), .B(n310), .Z(n591) );
  XNOR2_X1 U366 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n312), .B(KEYINPUT17), .ZN(n313) );
  XOR2_X1 U368 ( .A(n313), .B(KEYINPUT18), .Z(n315) );
  XNOR2_X1 U369 ( .A(G169GAT), .B(G176GAT), .ZN(n314) );
  XOR2_X1 U370 ( .A(n315), .B(n314), .Z(n420) );
  XOR2_X1 U371 ( .A(G43GAT), .B(G134GAT), .Z(n393) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G71GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n316), .B(G120GAT), .ZN(n369) );
  XOR2_X1 U374 ( .A(n393), .B(n369), .Z(n318) );
  NAND2_X1 U375 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U377 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n320) );
  XNOR2_X1 U378 ( .A(G190GAT), .B(KEYINPUT65), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U380 ( .A(n322), .B(n321), .Z(n324) );
  XOR2_X1 U381 ( .A(G113GAT), .B(G15GAT), .Z(n354) );
  XOR2_X1 U382 ( .A(KEYINPUT0), .B(G127GAT), .Z(n426) );
  XNOR2_X1 U383 ( .A(n354), .B(n426), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U385 ( .A(n420), .B(n325), .Z(n538) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .Z(n357) );
  XOR2_X1 U387 ( .A(G50GAT), .B(G162GAT), .Z(n394) );
  XNOR2_X1 U388 ( .A(n357), .B(n394), .ZN(n328) );
  XOR2_X1 U389 ( .A(G78GAT), .B(G148GAT), .Z(n327) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n368) );
  XNOR2_X1 U392 ( .A(n328), .B(n368), .ZN(n334) );
  XOR2_X1 U393 ( .A(G155GAT), .B(KEYINPUT82), .Z(n330) );
  XNOR2_X1 U394 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n430) );
  XOR2_X1 U396 ( .A(n430), .B(KEYINPUT22), .Z(n332) );
  NAND2_X1 U397 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U398 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U399 ( .A(n334), .B(n333), .Z(n344) );
  XNOR2_X1 U400 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n335), .B(KEYINPUT80), .ZN(n339) );
  XNOR2_X1 U402 ( .A(G197GAT), .B(G218GAT), .ZN(n337) );
  XOR2_X1 U403 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n341) );
  XNOR2_X1 U404 ( .A(G204GAT), .B(KEYINPUT83), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n412), .B(n342), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n467) );
  XOR2_X1 U408 ( .A(KEYINPUT29), .B(G197GAT), .Z(n346) );
  XNOR2_X1 U409 ( .A(G169GAT), .B(G50GAT), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U411 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n348) );
  XNOR2_X1 U412 ( .A(KEYINPUT68), .B(KEYINPUT71), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n363) );
  XNOR2_X1 U415 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n351), .B(KEYINPUT7), .ZN(n391) );
  XOR2_X1 U417 ( .A(n391), .B(KEYINPUT30), .Z(n353) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n361) );
  XOR2_X1 U421 ( .A(G43GAT), .B(G36GAT), .Z(n359) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U425 ( .A(n363), .B(n362), .Z(n506) );
  INV_X1 U426 ( .A(n506), .ZN(n581) );
  XNOR2_X1 U427 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n380) );
  XNOR2_X1 U428 ( .A(G204GAT), .B(G92GAT), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n364), .B(G64GAT), .ZN(n416) );
  XOR2_X1 U430 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n366) );
  NAND2_X1 U431 ( .A1(G230GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U433 ( .A(n367), .B(KEYINPUT31), .Z(n371) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n372), .B(KEYINPUT13), .ZN(n373) );
  XOR2_X1 U437 ( .A(G85GAT), .B(G57GAT), .Z(n425) );
  XOR2_X1 U438 ( .A(G176GAT), .B(n425), .Z(n374) );
  NAND2_X1 U439 ( .A1(n373), .A2(n374), .ZN(n378) );
  INV_X1 U440 ( .A(n373), .ZN(n376) );
  INV_X1 U441 ( .A(n374), .ZN(n375) );
  NAND2_X1 U442 ( .A1(n376), .A2(n375), .ZN(n377) );
  NAND2_X1 U443 ( .A1(n378), .A2(n377), .ZN(n379) );
  XOR2_X1 U444 ( .A(n416), .B(n379), .Z(n587) );
  XOR2_X1 U445 ( .A(n380), .B(n587), .Z(n504) );
  NAND2_X1 U446 ( .A1(n581), .A2(n504), .ZN(n381) );
  XNOR2_X1 U447 ( .A(n381), .B(KEYINPUT46), .ZN(n402) );
  XOR2_X1 U448 ( .A(KEYINPUT74), .B(G92GAT), .Z(n383) );
  XNOR2_X1 U449 ( .A(G85GAT), .B(KEYINPUT11), .ZN(n382) );
  XNOR2_X1 U450 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U451 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n385) );
  XNOR2_X1 U452 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n387), .B(n386), .ZN(n400) );
  NAND2_X1 U455 ( .A1(G232GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U457 ( .A(G36GAT), .B(G190GAT), .Z(n413) );
  XOR2_X1 U458 ( .A(n413), .B(n394), .Z(n396) );
  XNOR2_X1 U459 ( .A(G99GAT), .B(G218GAT), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n399) );
  NOR2_X1 U462 ( .A1(n572), .A2(n591), .ZN(n401) );
  AND2_X1 U463 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n403), .B(KEYINPUT47), .ZN(n410) );
  NAND2_X1 U465 ( .A1(n591), .A2(n593), .ZN(n405) );
  XNOR2_X1 U466 ( .A(KEYINPUT67), .B(KEYINPUT45), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  INV_X1 U468 ( .A(n587), .ZN(n455) );
  NAND2_X1 U469 ( .A1(n406), .A2(n455), .ZN(n407) );
  NOR2_X1 U470 ( .A1(n581), .A2(n407), .ZN(n408) );
  XOR2_X1 U471 ( .A(KEYINPUT106), .B(n408), .Z(n409) );
  AND2_X1 U472 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n411), .B(KEYINPUT48), .ZN(n534) );
  XOR2_X1 U474 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n419) );
  XNOR2_X1 U477 ( .A(G8GAT), .B(n416), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n524) );
  XNOR2_X1 U479 ( .A(KEYINPUT115), .B(n524), .ZN(n422) );
  NOR2_X1 U480 ( .A1(n534), .A2(n422), .ZN(n424) );
  XOR2_X1 U481 ( .A(n425), .B(G162GAT), .Z(n428) );
  XNOR2_X1 U482 ( .A(n426), .B(G134GAT), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U484 ( .A(n429), .B(KEYINPUT75), .Z(n435) );
  XOR2_X1 U485 ( .A(n430), .B(KEYINPUT86), .Z(n432) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(G29GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U490 ( .A(G148GAT), .B(G120GAT), .Z(n437) );
  XNOR2_X1 U491 ( .A(G113GAT), .B(G141GAT), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U493 ( .A(n439), .B(n438), .Z(n447) );
  XOR2_X1 U494 ( .A(KEYINPUT1), .B(KEYINPUT85), .Z(n441) );
  XNOR2_X1 U495 ( .A(KEYINPUT6), .B(KEYINPUT84), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U497 ( .A(KEYINPUT5), .B(KEYINPUT87), .Z(n443) );
  XNOR2_X1 U498 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U501 ( .A(n447), .B(n446), .Z(n521) );
  INV_X1 U502 ( .A(n521), .ZN(n535) );
  NAND2_X1 U503 ( .A1(n448), .A2(n535), .ZN(n579) );
  NOR2_X1 U504 ( .A1(n467), .A2(n579), .ZN(n451) );
  NOR2_X1 U505 ( .A1(n538), .A2(n452), .ZN(n573) );
  NAND2_X1 U506 ( .A1(n591), .A2(n573), .ZN(n454) );
  XNOR2_X1 U507 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n476) );
  NAND2_X1 U508 ( .A1(n455), .A2(n581), .ZN(n456) );
  XOR2_X1 U509 ( .A(KEYINPUT73), .B(n456), .Z(n488) );
  INV_X1 U510 ( .A(n591), .ZN(n457) );
  NOR2_X1 U511 ( .A1(n572), .A2(n457), .ZN(n458) );
  XOR2_X1 U512 ( .A(KEYINPUT16), .B(n458), .Z(n459) );
  XNOR2_X1 U513 ( .A(KEYINPUT77), .B(n459), .ZN(n474) );
  NAND2_X1 U514 ( .A1(n538), .A2(n467), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT26), .ZN(n578) );
  NOR2_X1 U516 ( .A1(n578), .A2(n468), .ZN(n466) );
  INV_X1 U517 ( .A(n524), .ZN(n511) );
  NOR2_X1 U518 ( .A1(n511), .A2(n538), .ZN(n462) );
  NOR2_X1 U519 ( .A1(n467), .A2(n462), .ZN(n463) );
  XNOR2_X1 U520 ( .A(KEYINPUT25), .B(n463), .ZN(n464) );
  NAND2_X1 U521 ( .A1(n464), .A2(n535), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n473) );
  XOR2_X1 U523 ( .A(n467), .B(KEYINPUT28), .Z(n516) );
  INV_X1 U524 ( .A(n516), .ZN(n541) );
  INV_X1 U525 ( .A(n468), .ZN(n537) );
  INV_X1 U526 ( .A(n538), .ZN(n527) );
  XNOR2_X1 U527 ( .A(KEYINPUT79), .B(n527), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n537), .A2(n469), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n541), .A2(n470), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n535), .A2(n471), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n474), .A2(n484), .ZN(n507) );
  NOR2_X1 U532 ( .A1(n488), .A2(n507), .ZN(n481) );
  NAND2_X1 U533 ( .A1(n481), .A2(n521), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U535 ( .A1(n524), .A2(n481), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT90), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U538 ( .A1(n481), .A2(n527), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n480), .ZN(G1326GAT) );
  XOR2_X1 U541 ( .A(G22GAT), .B(KEYINPUT91), .Z(n483) );
  NAND2_X1 U542 ( .A1(n481), .A2(n541), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(G1327GAT) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n492) );
  NAND2_X1 U545 ( .A1(n484), .A2(n593), .ZN(n485) );
  NOR2_X1 U546 ( .A1(n591), .A2(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(KEYINPUT92), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n520) );
  NOR2_X1 U549 ( .A1(n488), .A2(n520), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT93), .ZN(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT38), .B(n490), .ZN(n499) );
  NOR2_X1 U552 ( .A1(n535), .A2(n499), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  INV_X1 U554 ( .A(KEYINPUT94), .ZN(n494) );
  NOR2_X1 U555 ( .A1(n511), .A2(n499), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n495), .ZN(G1329GAT) );
  NOR2_X1 U558 ( .A1(n499), .A2(n538), .ZN(n497) );
  XNOR2_X1 U559 ( .A(KEYINPUT40), .B(KEYINPUT95), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NOR2_X1 U562 ( .A1(n516), .A2(n499), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT96), .B(n295), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n502) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT97), .B(n503), .ZN(n510) );
  INV_X1 U568 ( .A(n504), .ZN(n505) );
  INV_X1 U569 ( .A(n505), .ZN(n567) );
  NAND2_X1 U570 ( .A1(n506), .A2(n567), .ZN(n519) );
  NOR2_X1 U571 ( .A1(n519), .A2(n507), .ZN(n508) );
  XOR2_X1 U572 ( .A(KEYINPUT98), .B(n508), .Z(n515) );
  NOR2_X1 U573 ( .A1(n535), .A2(n515), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n511), .A2(n515), .ZN(n512) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n515), .A2(n538), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(KEYINPUT101), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  NOR2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT102), .ZN(n523) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n530), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(G1336GAT) );
  XOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT103), .Z(n526) );
  NAND2_X1 U588 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n530), .ZN(n528) );
  XNOR2_X1 U591 ( .A(KEYINPUT104), .B(n528), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT105), .B(KEYINPUT44), .Z(n532) );
  NAND2_X1 U594 ( .A1(n530), .A2(n541), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n553) );
  NOR2_X1 U599 ( .A1(n538), .A2(n553), .ZN(n539) );
  XNOR2_X1 U600 ( .A(n539), .B(KEYINPUT107), .ZN(n540) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U602 ( .A(KEYINPUT108), .B(n542), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n581), .A2(n549), .ZN(n543) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT109), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U606 ( .A1(n549), .A2(n567), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n546), .Z(G1341GAT) );
  NAND2_X1 U609 ( .A1(n549), .A2(n591), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT110), .Z(n551) );
  NAND2_X1 U613 ( .A1(n572), .A2(n549), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n552), .ZN(G1343GAT) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT112), .ZN(n556) );
  NOR2_X1 U617 ( .A1(n578), .A2(n553), .ZN(n554) );
  XOR2_X1 U618 ( .A(KEYINPUT111), .B(n554), .Z(n563) );
  NAND2_X1 U619 ( .A1(n581), .A2(n563), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT114), .Z(n558) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT113), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT52), .B(n559), .Z(n561) );
  NAND2_X1 U625 ( .A1(n563), .A2(n567), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n591), .A2(n563), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n572), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n581), .A2(n573), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  NAND2_X1 U634 ( .A1(n573), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT56), .Z(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1351GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n583) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT123), .B(n580), .Z(n594) );
  NAND2_X1 U647 ( .A1(n594), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(n584), .B(KEYINPUT59), .Z(n586) );
  XNOR2_X1 U650 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n589) );
  NAND2_X1 U653 ( .A1(n594), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G204GAT), .B(n590), .ZN(G1353GAT) );
  NAND2_X1 U656 ( .A1(n591), .A2(n594), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n596) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U661 ( .A(G218GAT), .B(n597), .ZN(G1355GAT) );
endmodule

