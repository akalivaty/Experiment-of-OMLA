//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n240), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  AND3_X1   g0052(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n249), .B2(new_n251), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G222), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n257), .B1(new_n258), .B2(new_n255), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT64), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n215), .B1(KEYINPUT65), .B2(new_n268), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n268), .A2(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n267), .A2(G274), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n265), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(G226), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n263), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G190), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(G200), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT67), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n209), .B2(new_n248), .ZN(new_n282));
  NAND4_X1  g0082(.A1(KEYINPUT67), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n215), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n264), .A2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G50), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n216), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G150), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n290), .A2(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n203), .A2(G50), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n216), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n284), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n289), .B(new_n298), .C1(G50), .C2(new_n285), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT9), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n278), .A2(new_n279), .A3(new_n280), .A4(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n255), .A2(G226), .A3(new_n256), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n250), .A2(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT66), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n307), .A2(G232), .A3(G1698), .A4(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n248), .B2(new_n205), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n262), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n272), .B1(G238), .B2(new_n274), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT70), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n311), .A2(new_n312), .B1(new_n313), .B2(KEYINPUT13), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(KEYINPUT13), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n312), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT13), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n320), .A2(G200), .A3(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n293), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n258), .B2(new_n291), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT11), .B1(new_n324), .B2(new_n284), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n285), .A2(G68), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT12), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n324), .A2(KEYINPUT11), .A3(new_n284), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n287), .A2(G68), .A3(new_n288), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n317), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n320), .A2(G169), .A3(new_n321), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n320), .A2(new_n335), .A3(G169), .A4(new_n321), .ZN(new_n336));
  INV_X1    g0136(.A(new_n316), .ZN(new_n337));
  OAI21_X1  g0137(.A(G179), .B1(new_n337), .B2(new_n314), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n332), .B1(new_n331), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n276), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n299), .C1(G179), .C2(new_n276), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n267), .A2(G274), .A3(new_n271), .ZN(new_n344));
  INV_X1    g0144(.A(G244), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n273), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n255), .A2(G232), .A3(new_n256), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n347), .B1(new_n206), .B2(new_n255), .C1(new_n259), .C2(new_n220), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n346), .B1(new_n348), .B2(new_n262), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n287), .A2(G77), .A3(new_n288), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT68), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n290), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n293), .B1(G20), .B2(G77), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT15), .B(G87), .Z(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n291), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n284), .B1(new_n258), .B2(new_n286), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n350), .A2(new_n341), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n349), .A2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n350), .A2(new_n303), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n349), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n353), .A2(new_n359), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n302), .A2(new_n340), .A3(new_n343), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G58), .A2(G68), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n203), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT3), .B(G33), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n375), .A2(new_n376), .A3(G20), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n249), .B2(new_n251), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT71), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n376), .C1(new_n375), .C2(G20), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT16), .B(new_n374), .C1(new_n382), .C2(new_n202), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n383), .A2(new_n284), .ZN(new_n384));
  INV_X1    g0184(.A(new_n374), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT73), .ZN(new_n386));
  AOI21_X1  g0186(.A(G20), .B1(new_n307), .B2(new_n308), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(KEYINPUT7), .ZN(new_n388));
  INV_X1    g0188(.A(new_n377), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n216), .B1(new_n253), .B2(new_n254), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(KEYINPUT73), .A3(new_n376), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n385), .B1(new_n392), .B2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n384), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n282), .A2(new_n215), .A3(new_n283), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n285), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n354), .A2(new_n288), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n396), .A2(new_n397), .B1(new_n285), .B2(new_n354), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G232), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n273), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n272), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n249), .A2(new_n251), .A3(G226), .A4(G1698), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT74), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n375), .A2(KEYINPUT74), .A3(G226), .A4(G1698), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT75), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n249), .A2(new_n251), .A3(G223), .A4(new_n256), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n407), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n262), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n405), .B2(new_n406), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n408), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n303), .B(new_n402), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n344), .B1(new_n400), .B2(new_n273), .ZN(new_n418));
  INV_X1    g0218(.A(new_n262), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n415), .B2(new_n408), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n407), .A2(new_n412), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT75), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n417), .B1(new_n423), .B2(G200), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n394), .A2(new_n399), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT76), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT76), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n394), .A2(new_n424), .A3(new_n427), .A4(new_n399), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n394), .A2(new_n424), .A3(new_n430), .A4(new_n399), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n394), .A2(new_n399), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n423), .A2(G179), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n341), .B2(new_n423), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n434), .B2(new_n436), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT77), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n426), .A2(new_n442), .A3(KEYINPUT17), .A4(new_n428), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n433), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(KEYINPUT78), .A2(G97), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT78), .A2(G97), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n248), .ZN(new_n448));
  AOI21_X1  g0248(.A(G20), .B1(G33), .B2(G283), .ZN(new_n449));
  INV_X1    g0249(.A(G116), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n448), .A2(new_n449), .B1(G20), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n284), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT20), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(new_n449), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(G20), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n284), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT86), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n451), .A2(KEYINPUT86), .A3(KEYINPUT20), .A4(new_n284), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n454), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n285), .A2(G116), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT85), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n287), .B1(G1), .B2(new_n248), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n465), .B2(G116), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n461), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n461), .B2(new_n466), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n307), .A2(new_n308), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G303), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT83), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n375), .A2(G257), .A3(new_n256), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n375), .A2(G264), .A3(G1698), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G303), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n307), .B2(new_n308), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n475), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT83), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n262), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT84), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n476), .A2(new_n480), .A3(new_n483), .A4(new_n262), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n271), .A2(G274), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n486), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n271), .A2(new_n489), .A3(G270), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT82), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n482), .A2(new_n484), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G169), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT88), .B1(new_n470), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT21), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  OAI211_X1 g0297(.A(KEYINPUT88), .B(new_n497), .C1(new_n470), .C2(new_n494), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n482), .A2(G179), .A3(new_n484), .A4(new_n492), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n468), .B2(new_n469), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n493), .A2(G200), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n470), .B(new_n502), .C1(new_n303), .C2(new_n493), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n496), .A2(new_n498), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n375), .A2(new_n216), .A3(G87), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n506), .A2(KEYINPUT89), .A3(KEYINPUT22), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT89), .B1(new_n506), .B2(KEYINPUT22), .ZN(new_n508));
  OR3_X1    g0308(.A1(new_n221), .A2(KEYINPUT22), .A3(G20), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n507), .A2(new_n508), .B1(new_n471), .B2(new_n509), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n216), .A2(KEYINPUT23), .A3(G107), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT23), .B1(new_n216), .B2(G107), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT90), .ZN(new_n514));
  OAI221_X1 g0314(.A(new_n511), .B1(G20), .B2(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n514), .B2(new_n513), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n505), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n510), .A2(new_n505), .A3(new_n516), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n395), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n375), .A2(G257), .A3(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G294), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n375), .A2(new_n256), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n222), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n271), .A2(new_n489), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n524), .A2(new_n262), .B1(new_n525), .B2(G264), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n488), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G200), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n303), .B2(new_n527), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n286), .A2(new_n206), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT25), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n465), .B2(G107), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n520), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n527), .A2(new_n341), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G179), .B2(new_n527), .ZN(new_n536));
  INV_X1    g0336(.A(new_n519), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n284), .B1(new_n537), .B2(new_n517), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n538), .B2(new_n532), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n525), .A2(G257), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n541), .A2(new_n488), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n375), .A2(G244), .A3(new_n256), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n543), .A2(new_n544), .B1(G33), .B2(G283), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n345), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n307), .A2(new_n256), .A3(new_n308), .A4(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n307), .A2(G250), .A3(G1698), .A4(new_n308), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n262), .ZN(new_n550));
  AOI21_X1  g0350(.A(G169), .B1(new_n542), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n542), .A2(new_n550), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n361), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n286), .A2(new_n205), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n465), .A2(G97), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n447), .A2(KEYINPUT6), .A3(new_n206), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT6), .B1(new_n207), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n559), .A2(new_n216), .B1(new_n258), .B2(new_n294), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n392), .B2(G107), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n554), .B(new_n555), .C1(new_n561), .C2(new_n395), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n553), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n562), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n552), .A2(G190), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n552), .A2(KEYINPUT79), .A3(new_n365), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n542), .A2(new_n550), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n567), .B1(new_n568), .B2(G200), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n375), .A2(new_n216), .A3(G68), .ZN(new_n571));
  INV_X1    g0371(.A(new_n447), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n291), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(KEYINPUT19), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n447), .A2(G87), .A3(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(new_n216), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n284), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n357), .A2(new_n286), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n221), .C2(new_n464), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n375), .A2(G244), .A3(G1698), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n512), .C1(new_n523), .C2(new_n220), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n486), .A2(new_n222), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n582), .A2(new_n262), .B1(new_n271), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n271), .A2(G274), .A3(new_n486), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT80), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n271), .A2(new_n587), .A3(G274), .A4(new_n486), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n303), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n365), .B1(new_n584), .B2(new_n589), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n580), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n465), .A2(new_n356), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n578), .A3(new_n579), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n590), .A2(G169), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n584), .A2(new_n589), .A3(G179), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT81), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(KEYINPUT81), .A3(new_n598), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n593), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n540), .A2(new_n563), .A3(new_n570), .A4(new_n603), .ZN(new_n604));
  NOR4_X1   g0404(.A1(new_n370), .A2(new_n444), .A3(new_n504), .A4(new_n604), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n339), .A2(new_n331), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n360), .A2(new_n362), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n332), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n433), .A3(new_n443), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n441), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n302), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n611), .A2(new_n343), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n370), .A2(new_n444), .ZN(new_n613));
  INV_X1    g0413(.A(new_n534), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n599), .A2(new_n595), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n593), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n563), .A2(new_n614), .A3(new_n570), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n539), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n496), .A2(new_n498), .A3(new_n501), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  INV_X1    g0422(.A(new_n563), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n603), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n580), .A2(new_n591), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n615), .B1(new_n626), .B2(new_n592), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT91), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n553), .B2(new_n562), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n625), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n630), .B2(new_n622), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n621), .A2(new_n615), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n612), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT92), .ZN(G369));
  AND3_X1   g0435(.A1(new_n496), .A2(new_n498), .A3(new_n501), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n264), .A2(new_n216), .A3(G13), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT93), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g0441(.A(KEYINPUT94), .B(G343), .Z(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n470), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n636), .A2(new_n503), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n636), .B2(new_n646), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n643), .B1(new_n520), .B2(new_n533), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n539), .B1(new_n614), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n539), .B2(new_n644), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n636), .A2(new_n643), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n652), .B1(new_n539), .B2(new_n644), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(G399));
  NAND2_X1  g0456(.A1(new_n575), .A2(new_n450), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n210), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(G1), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n213), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  INV_X1    g0464(.A(G330), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n504), .A2(new_n604), .A3(new_n643), .ZN(new_n666));
  NOR2_X1   g0466(.A1(KEYINPUT96), .A2(KEYINPUT30), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n526), .A2(new_n584), .A3(new_n589), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT95), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT95), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n526), .A2(new_n584), .A3(new_n589), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n552), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n667), .B1(new_n673), .B2(new_n499), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n527), .A2(new_n590), .A3(new_n361), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n493), .A2(new_n568), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n667), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n568), .B1(new_n669), .B2(new_n671), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n500), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n674), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT31), .B1(new_n680), .B2(new_n643), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT97), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n682), .A2(KEYINPUT97), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT98), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n666), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT98), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n665), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n603), .A2(new_n623), .ZN(new_n690));
  MUX2_X1   g0490(.A(new_n690), .B(new_n630), .S(KEYINPUT26), .Z(new_n691));
  AOI21_X1  g0491(.A(new_n616), .B1(new_n618), .B2(new_n620), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n643), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI211_X1 g0495(.A(KEYINPUT29), .B(new_n643), .C1(new_n692), .C2(new_n631), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n689), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n664), .B1(new_n697), .B2(G1), .ZN(G364));
  AND2_X1   g0498(.A1(new_n216), .A2(G13), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n264), .B1(new_n699), .B2(G45), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n660), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n649), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(G330), .B2(new_n648), .ZN(new_n704));
  INV_X1    g0504(.A(new_n702), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n216), .A2(G179), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(new_n303), .A3(G200), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT100), .Z(new_n708));
  NOR2_X1   g0508(.A1(new_n303), .A2(new_n365), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n706), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT101), .Z(new_n711));
  AOI22_X1  g0511(.A1(G283), .A2(new_n708), .B1(new_n711), .B2(G303), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G190), .A2(G200), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G329), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n216), .A2(new_n361), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n713), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(G326), .A2(new_n719), .B1(new_n721), .B2(G311), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n303), .A2(G179), .A3(G200), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n216), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n255), .B1(G294), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n712), .A2(new_n716), .A3(new_n722), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n717), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n728), .A2(new_n365), .A3(G190), .ZN(new_n729));
  XNOR2_X1  g0529(.A(KEYINPUT33), .B(G317), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n728), .A2(new_n303), .A3(G200), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(G322), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT102), .Z(new_n733));
  NAND2_X1  g0533(.A1(new_n708), .A2(G107), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n718), .A2(new_n241), .B1(new_n720), .B2(new_n258), .ZN(new_n735));
  INV_X1    g0535(.A(new_n710), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(G87), .B2(new_n736), .ZN(new_n737));
  AOI22_X1  g0537(.A1(G58), .A2(new_n731), .B1(new_n729), .B2(G68), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n734), .A2(new_n255), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G159), .ZN(new_n740));
  OR3_X1    g0540(.A1(new_n714), .A2(KEYINPUT32), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT32), .B1(new_n714), .B2(new_n740), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n741), .B(new_n742), .C1(new_n205), .C2(new_n724), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n727), .A2(new_n733), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n215), .B1(G20), .B2(new_n341), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n705), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n745), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n659), .A2(new_n375), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n246), .A2(new_n485), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n753), .B(new_n754), .C1(new_n485), .C2(new_n214), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n255), .A2(new_n210), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n210), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT99), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n755), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n746), .B1(new_n751), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT103), .ZN(new_n764));
  INV_X1    g0564(.A(new_n749), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n648), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n704), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(G396));
  NOR2_X1   g0568(.A1(new_n745), .A2(new_n747), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT104), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n705), .B1(new_n771), .B2(new_n258), .ZN(new_n772));
  INV_X1    g0572(.A(new_n745), .ZN(new_n773));
  INV_X1    g0573(.A(new_n708), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n221), .ZN(new_n775));
  INV_X1    g0575(.A(new_n711), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n206), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G303), .A2(new_n719), .B1(new_n721), .B2(G116), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n778), .B(new_n471), .C1(new_n205), .C2(new_n724), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n729), .A2(G283), .B1(G311), .B2(new_n715), .ZN(new_n780));
  INV_X1    g0580(.A(G294), .ZN(new_n781));
  INV_X1    g0581(.A(new_n731), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n775), .A2(new_n777), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n731), .A2(G143), .B1(new_n719), .B2(G137), .ZN(new_n785));
  INV_X1    g0585(.A(new_n729), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n785), .B1(new_n292), .B2(new_n786), .C1(new_n740), .C2(new_n720), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT105), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT34), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n708), .A2(G68), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n711), .A2(G50), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n725), .A2(G58), .ZN(new_n793));
  INV_X1    g0593(.A(new_n375), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n715), .B2(G132), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n791), .A2(new_n792), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n788), .B2(new_n789), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n784), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n367), .A2(new_n643), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT106), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n367), .A2(KEYINPUT106), .A3(new_n643), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n607), .B1(new_n368), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n363), .A2(new_n644), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n772), .B1(new_n773), .B2(new_n798), .C1(new_n807), .C2(new_n748), .ZN(new_n808));
  INV_X1    g0608(.A(new_n689), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n643), .B1(new_n692), .B2(new_n631), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(new_n807), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n702), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n809), .A2(new_n811), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(G384));
  INV_X1    g0615(.A(new_n559), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT35), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(KEYINPUT35), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n817), .A2(G116), .A3(new_n217), .A4(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT36), .Z(new_n820));
  NAND3_X1  g0620(.A1(new_n372), .A2(new_n214), .A3(G77), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n264), .B(G13), .C1(new_n821), .C2(new_n242), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT110), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n641), .B1(new_n438), .B2(new_n440), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n632), .A2(new_n644), .A3(new_n807), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n805), .ZN(new_n827));
  OR3_X1    g0627(.A1(new_n317), .A2(new_n322), .A3(new_n331), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n643), .A2(new_n331), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n606), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n331), .B(new_n643), .C1(new_n332), .C2(new_n339), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n374), .B1(new_n382), .B2(new_n202), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT16), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n383), .A2(new_n284), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n399), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n641), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n444), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n436), .B2(new_n839), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n426), .A2(new_n428), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT107), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT107), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n846), .A3(KEYINPUT37), .ZN(new_n847));
  XOR2_X1   g0647(.A(KEYINPUT109), .B(KEYINPUT37), .Z(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT7), .B1(new_n471), .B2(new_n216), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n377), .B1(new_n849), .B2(KEYINPUT73), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n202), .B1(new_n850), .B2(new_n388), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n835), .B1(new_n851), .B2(new_n385), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n398), .B1(new_n852), .B2(new_n384), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n848), .B1(new_n853), .B2(new_n641), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT108), .B1(new_n434), .B2(new_n436), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n426), .A2(new_n428), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n434), .A2(KEYINPUT108), .A3(new_n436), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n845), .A2(new_n847), .A3(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n841), .A2(new_n860), .A3(KEYINPUT38), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n841), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n824), .B(new_n825), .C1(new_n833), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n606), .A2(new_n643), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n841), .A2(new_n860), .A3(KEYINPUT38), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n853), .A2(new_n641), .ZN(new_n868));
  INV_X1    g0668(.A(new_n848), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n437), .A2(new_n425), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n869), .B1(new_n870), .B2(new_n868), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n444), .A2(new_n868), .B1(new_n859), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n867), .B1(KEYINPUT38), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n865), .A2(new_n866), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n864), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n825), .B1(new_n833), .B2(new_n863), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT110), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n613), .B1(new_n695), .B2(new_n696), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n612), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n880), .B(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n666), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n679), .A2(new_n676), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n677), .B1(new_n500), .B2(new_n678), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n643), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT31), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n613), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT111), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n806), .B1(new_n830), .B2(new_n831), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n666), .B2(new_n891), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n444), .A2(new_n868), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n859), .A2(new_n871), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n898), .B1(new_n861), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n841), .A2(new_n860), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n867), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n896), .B(new_n907), .C1(new_n666), .C2(new_n891), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n902), .A2(KEYINPUT40), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n895), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n895), .A2(new_n910), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(G330), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n883), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n264), .B2(new_n699), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n883), .A2(new_n913), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n823), .B1(new_n915), .B2(new_n916), .ZN(G367));
  OAI221_X1 g0717(.A(new_n750), .B1(new_n210), .B2(new_n357), .C1(new_n236), .C2(new_n753), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT116), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n705), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n729), .A2(G159), .B1(G137), .B2(new_n715), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n922), .B1(new_n201), .B2(new_n710), .C1(new_n292), .C2(new_n782), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n719), .A2(G143), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n924), .B1(new_n241), .B2(new_n720), .C1(new_n258), .C2(new_n707), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n724), .A2(new_n202), .ZN(new_n926));
  OR4_X1    g0726(.A1(new_n471), .A2(new_n923), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(G283), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n782), .A2(new_n477), .B1(new_n720), .B2(new_n928), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n375), .B(new_n929), .C1(G311), .C2(new_n719), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n710), .A2(new_n450), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n930), .B1(KEYINPUT46), .B2(new_n931), .C1(new_n206), .C2(new_n724), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n711), .A2(KEYINPUT46), .A3(G116), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n729), .A2(G294), .ZN(new_n934));
  INV_X1    g0734(.A(new_n707), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n447), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n715), .A2(G317), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n933), .A2(new_n934), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n927), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT47), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n921), .B1(new_n940), .B2(new_n745), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n580), .A2(new_n643), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n617), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n615), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n749), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n570), .B(new_n563), .C1(new_n564), .C2(new_n644), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n563), .B2(new_n644), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n654), .A2(new_n652), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n563), .B1(new_n949), .B2(new_n619), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n644), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT113), .Z(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n959));
  NAND2_X1  g0759(.A1(new_n946), .A2(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n956), .A2(new_n958), .B1(KEYINPUT114), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(KEYINPUT114), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n653), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n950), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT115), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT115), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n964), .A2(new_n971), .A3(new_n968), .A4(new_n965), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n966), .A2(new_n969), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n655), .A2(new_n950), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT45), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n655), .A2(new_n950), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n967), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n977), .A2(new_n653), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n654), .B(new_n652), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n649), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n697), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n697), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n660), .B(KEYINPUT41), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n701), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n948), .B1(new_n975), .B2(new_n990), .ZN(G387));
  OAI22_X1  g0791(.A1(new_n786), .A2(new_n290), .B1(new_n258), .B2(new_n710), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n794), .B(new_n992), .C1(G150), .C2(new_n715), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n725), .A2(new_n356), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n708), .A2(G97), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n782), .A2(new_n241), .B1(new_n718), .B2(new_n740), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G68), .B2(new_n721), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n375), .B1(new_n715), .B2(G326), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n724), .A2(new_n928), .B1(new_n710), .B2(new_n781), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n731), .A2(G317), .B1(new_n719), .B2(G322), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n729), .A2(G311), .B1(G303), .B2(new_n721), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT49), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n999), .B1(new_n450), .B2(new_n707), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n998), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n773), .B1(new_n1010), .B2(KEYINPUT117), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(KEYINPUT117), .B2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n752), .B1(new_n233), .B2(new_n485), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n658), .B2(new_n756), .ZN(new_n1014));
  AOI21_X1  g0814(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT50), .B1(new_n290), .B2(G50), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n290), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n658), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1014), .A2(new_n1018), .B1(new_n206), .B2(new_n659), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1012), .B(new_n702), .C1(new_n751), .C2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n652), .A2(new_n765), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT118), .Z(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n985), .B2(new_n701), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n986), .A2(new_n660), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n697), .A2(new_n985), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(G393));
  AND2_X1   g0827(.A1(new_n981), .A2(new_n982), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n986), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n661), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1029), .B1(new_n981), .B2(new_n982), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(KEYINPUT121), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT121), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n660), .B1(new_n983), .B2(new_n986), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n1031), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1028), .A2(new_n701), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n750), .B1(new_n210), .B2(new_n572), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n240), .B2(new_n752), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n731), .A2(G159), .B1(new_n719), .B2(G150), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n775), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G68), .A2(new_n736), .B1(new_n715), .B2(G143), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n729), .A2(G50), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n725), .A2(G77), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n794), .B1(new_n721), .B2(new_n354), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n731), .A2(G311), .B1(new_n719), .B2(G317), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G283), .A2(new_n736), .B1(new_n715), .B2(G322), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n729), .A2(G303), .B1(G294), .B2(new_n721), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n255), .B1(G116), .B2(new_n725), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n734), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1044), .A2(new_n1049), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n705), .B(new_n1040), .C1(new_n1056), .C2(new_n745), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT120), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n950), .B2(new_n765), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1038), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1037), .A2(new_n1061), .ZN(G390));
  NAND3_X1  g0862(.A1(new_n893), .A2(G330), .A3(new_n896), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n866), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n865), .A2(new_n875), .B1(new_n833), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n805), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n693), .B2(new_n804), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n832), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n873), .B(new_n1065), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1064), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1067), .B1(new_n810), .B2(new_n807), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1065), .B1(new_n1073), .B2(new_n1069), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n906), .A2(new_n874), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n899), .A2(new_n900), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n904), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT39), .B1(new_n1077), .B2(new_n867), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n689), .A2(new_n807), .A3(new_n832), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1070), .A3(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1072), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n893), .A2(G330), .A3(new_n613), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n881), .A2(new_n612), .A3(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT122), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n832), .B1(new_n689), .B2(new_n807), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n827), .B1(new_n1086), .B2(new_n1064), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n893), .A2(G330), .A3(new_n807), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n1069), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1080), .A2(new_n1068), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1082), .A2(new_n1085), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1085), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1072), .A2(new_n1081), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1095), .A3(new_n660), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1082), .A2(new_n701), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n747), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n702), .B1(new_n770), .B2(new_n354), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n711), .A2(G87), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n721), .A2(new_n447), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n731), .A2(G116), .B1(new_n719), .B2(G283), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n791), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n729), .A2(G107), .B1(G294), .B2(new_n715), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n471), .A3(new_n1047), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n710), .A2(new_n292), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT54), .B(G143), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G128), .A2(new_n719), .B1(new_n721), .B2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n729), .A2(G137), .B1(G125), .B2(new_n715), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1107), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n731), .A2(G132), .B1(G50), .B2(new_n935), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n255), .C1(new_n740), .C2(new_n724), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1103), .A2(new_n1105), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1099), .B1(new_n1115), .B2(new_n745), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1098), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n1097), .A3(new_n1117), .ZN(G378));
  INV_X1    g0918(.A(KEYINPUT125), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n839), .A2(new_n299), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n302), .A2(new_n343), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n302), .B2(new_n343), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n910), .B2(new_n665), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n907), .B1(new_n873), .B2(new_n898), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n908), .B1(new_n905), .B2(new_n867), .ZN(new_n1131));
  OAI211_X1 g0931(.A(G330), .B(new_n1127), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT124), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1119), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(KEYINPUT124), .B(KEYINPUT125), .C1(new_n1129), .C2(new_n1132), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n880), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1132), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n909), .B1(new_n861), .B2(new_n862), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n897), .B1(new_n1077), .B2(new_n867), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n907), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1127), .B1(new_n1141), .B2(G330), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1134), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT125), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n880), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1133), .A2(new_n1134), .A3(new_n1119), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1137), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT122), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1084), .B(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1082), .B2(new_n1091), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT57), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n880), .A2(new_n1133), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n877), .A2(new_n879), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT57), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n660), .B1(new_n1157), .B2(new_n1151), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1128), .A2(new_n747), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n702), .B1(new_n770), .B2(G50), .ZN(new_n1161));
  INV_X1    g0961(.A(G41), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n794), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n729), .B2(G97), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n450), .B2(new_n718), .C1(new_n206), .C2(new_n782), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n357), .A2(new_n720), .B1(new_n258), .B2(new_n710), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n707), .A2(new_n201), .B1(new_n714), .B2(new_n928), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1165), .A2(new_n926), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT58), .Z(new_n1169));
  OAI211_X1 g0969(.A(new_n1163), .B(new_n241), .C1(G33), .C2(G41), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n721), .A2(G137), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n731), .A2(G128), .B1(new_n719), .B2(G125), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n729), .A2(G132), .B1(new_n736), .B2(new_n1109), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n725), .A2(G150), .ZN(new_n1174));
  AND4_X1   g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n248), .B(new_n1162), .C1(new_n707), .C2(new_n740), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G124), .B2(new_n715), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1169), .B(new_n1170), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT123), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n773), .B1(new_n1182), .B2(KEYINPUT123), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1161), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1160), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1148), .B2(new_n701), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1159), .A2(new_n1188), .ZN(G375));
  NAND2_X1  g0989(.A1(new_n1069), .A2(new_n747), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n702), .B1(new_n770), .B2(G68), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1109), .A2(new_n729), .B1(new_n731), .B2(G137), .ZN(new_n1192));
  INV_X1    g0992(.A(G132), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n718), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G159), .B2(new_n711), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n725), .A2(G50), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n794), .B1(new_n935), .B2(G58), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G150), .A2(new_n721), .B1(new_n715), .B2(G128), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n471), .B1(new_n477), .B2(new_n714), .C1(new_n782), .C2(new_n928), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n356), .B2(new_n725), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n258), .B2(new_n774), .C1(new_n205), .C2(new_n776), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G294), .A2(new_n719), .B1(new_n721), .B2(G107), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n450), .B2(new_n786), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT126), .Z(new_n1205));
  OAI21_X1  g1005(.A(new_n1199), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1191), .B1(new_n1206), .B2(new_n745), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1091), .A2(new_n701), .B1(new_n1190), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1093), .A2(new_n989), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1091), .A2(new_n1085), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(G381));
  NAND2_X1  g1011(.A1(new_n987), .A2(new_n989), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n700), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n970), .A2(new_n972), .B1(new_n966), .B2(new_n969), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1213), .A2(new_n1214), .B1(new_n947), .B2(new_n941), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1060), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  OR4_X1    g1018(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1218), .ZN(G407));
  AND3_X1   g1019(.A1(new_n1096), .A2(new_n1097), .A3(new_n1117), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n642), .A2(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G375), .C2(new_n1223), .ZN(G409));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1091), .B2(new_n1085), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(new_n1210), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n1087), .A4(new_n1090), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n660), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1208), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(G384), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G384), .B(new_n1208), .C1(new_n1227), .C2(new_n1229), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1222), .A2(G2897), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G378), .B(new_n1188), .C1(new_n1153), .C2(new_n1158), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n988), .B(new_n1151), .C1(new_n1137), .C2(new_n1147), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1156), .A2(new_n701), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1186), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1220), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1221), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT61), .B1(new_n1240), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1247), .B2(new_n1234), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G387), .A2(new_n1216), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT127), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(G393), .B(G396), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G390), .A2(new_n1215), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1251), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1255), .A2(new_n1251), .A3(new_n1258), .A4(new_n1253), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1222), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1234), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(KEYINPUT63), .A3(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1248), .A2(new_n1250), .A3(new_n1260), .A4(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1261), .A2(new_n1265), .A3(new_n1262), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1261), .B2(new_n1239), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1265), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1264), .B1(new_n1270), .B2(new_n1260), .ZN(G405));
  AOI22_X1  g1071(.A1(new_n1252), .A2(new_n1253), .B1(new_n1255), .B2(new_n1251), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1259), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G378), .B1(new_n1159), .B2(new_n1188), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1241), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1262), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G375), .A2(new_n1220), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1234), .A3(new_n1241), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1274), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1274), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(G402));
endmodule


