

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U559 ( .A1(n1001), .A2(n731), .ZN(n735) );
  NOR2_X2 U560 ( .A1(n791), .A2(n790), .ZN(n800) );
  XNOR2_X1 U561 ( .A(n752), .B(n751), .ZN(n759) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n751) );
  NOR2_X1 U563 ( .A1(n722), .A2(n721), .ZN(n753) );
  INV_X1 U564 ( .A(n753), .ZN(n771) );
  INV_X1 U565 ( .A(G2104), .ZN(n528) );
  NOR2_X1 U566 ( .A1(G651), .A2(n635), .ZN(n643) );
  NAND2_X1 U567 ( .A1(n528), .A2(G2105), .ZN(n526) );
  XNOR2_X2 U568 ( .A(n526), .B(KEYINPUT65), .ZN(n889) );
  NAND2_X1 U569 ( .A1(n889), .A2(G125), .ZN(n527) );
  XNOR2_X1 U570 ( .A(KEYINPUT66), .B(n527), .ZN(n531) );
  NOR2_X1 U571 ( .A1(G2105), .A2(n528), .ZN(n884) );
  NAND2_X1 U572 ( .A1(n884), .A2(G101), .ZN(n529) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  NAND2_X1 U574 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U575 ( .A(n532), .B(KEYINPUT67), .ZN(n686) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XOR2_X1 U577 ( .A(KEYINPUT17), .B(n533), .Z(n885) );
  NAND2_X1 U578 ( .A1(G137), .A2(n885), .ZN(n683) );
  AND2_X1 U579 ( .A1(n686), .A2(n683), .ZN(n535) );
  AND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U581 ( .A1(n888), .A2(G113), .ZN(n534) );
  XNOR2_X1 U582 ( .A(KEYINPUT68), .B(n534), .ZN(n682) );
  AND2_X1 U583 ( .A1(n535), .A2(n682), .ZN(G160) );
  INV_X1 U584 ( .A(G651), .ZN(n541) );
  NOR2_X1 U585 ( .A1(G543), .A2(n541), .ZN(n537) );
  XNOR2_X1 U586 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n537), .B(n536), .ZN(n639) );
  NAND2_X1 U588 ( .A1(G65), .A2(n639), .ZN(n540) );
  NOR2_X1 U589 ( .A1(G543), .A2(G651), .ZN(n538) );
  XNOR2_X1 U590 ( .A(n538), .B(KEYINPUT64), .ZN(n638) );
  NAND2_X1 U591 ( .A1(G91), .A2(n638), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n545) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  NOR2_X1 U594 ( .A1(n635), .A2(n541), .ZN(n642) );
  NAND2_X1 U595 ( .A1(G78), .A2(n642), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G53), .A2(n643), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U598 ( .A1(n545), .A2(n544), .ZN(G299) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U600 ( .A1(G99), .A2(n884), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G111), .A2(n888), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G123), .A2(n889), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n548), .B(KEYINPUT18), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n885), .A2(G135), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n552), .A2(n551), .ZN(n931) );
  XNOR2_X1 U608 ( .A(n931), .B(G2096), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n553), .B(KEYINPUT77), .ZN(n554) );
  OR2_X1 U610 ( .A1(G2100), .A2(n554), .ZN(G156) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  INV_X1 U612 ( .A(G132), .ZN(G219) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  NAND2_X1 U614 ( .A1(n642), .A2(G75), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G88), .A2(n638), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT82), .B(n557), .Z(n561) );
  NAND2_X1 U618 ( .A1(G62), .A2(n639), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G50), .A2(n643), .ZN(n558) );
  AND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(G303) );
  INV_X1 U622 ( .A(G303), .ZN(G166) );
  NAND2_X1 U623 ( .A1(n638), .A2(G89), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n562), .B(KEYINPUT74), .ZN(n563) );
  XNOR2_X1 U625 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G76), .A2(n642), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U628 ( .A(n566), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n643), .A2(G51), .ZN(n567) );
  XOR2_X1 U630 ( .A(KEYINPUT75), .B(n567), .Z(n569) );
  NAND2_X1 U631 ( .A1(n639), .A2(G63), .ZN(n568) );
  NAND2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U635 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U637 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n575) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G223) );
  XOR2_X1 U640 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n577) );
  INV_X1 U641 ( .A(G223), .ZN(n837) );
  NAND2_X1 U642 ( .A1(G567), .A2(n837), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G234) );
  NAND2_X1 U644 ( .A1(G56), .A2(n639), .ZN(n578) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n578), .Z(n584) );
  NAND2_X1 U646 ( .A1(G81), .A2(n638), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G68), .A2(n642), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  NOR2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U652 ( .A1(n643), .A2(G43), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n1001) );
  INV_X1 U654 ( .A(G860), .ZN(n606) );
  OR2_X1 U655 ( .A1(n1001), .A2(n606), .ZN(G153) );
  NAND2_X1 U656 ( .A1(n642), .A2(G77), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G90), .A2(n638), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U659 ( .A(KEYINPUT9), .B(n589), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G64), .A2(n639), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G52), .A2(n643), .ZN(n590) );
  AND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(G301) );
  INV_X1 U664 ( .A(G301), .ZN(G171) );
  INV_X1 U665 ( .A(G868), .ZN(n658) );
  NOR2_X1 U666 ( .A1(n658), .A2(G171), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT73), .ZN(n603) );
  NAND2_X1 U668 ( .A1(G66), .A2(n639), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G92), .A2(n638), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G79), .A2(n642), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G54), .A2(n643), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U675 ( .A(KEYINPUT15), .B(n601), .Z(n995) );
  OR2_X1 U676 ( .A1(G868), .A2(n995), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(G284) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U679 ( .A1(G286), .A2(n658), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U681 ( .A1(G559), .A2(n606), .ZN(n607) );
  XNOR2_X1 U682 ( .A(KEYINPUT76), .B(n607), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n608), .A2(n995), .ZN(n609) );
  XNOR2_X1 U684 ( .A(KEYINPUT16), .B(n609), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n1001), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G868), .A2(n995), .ZN(n610) );
  NOR2_X1 U687 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U688 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U689 ( .A1(G67), .A2(n639), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n613), .B(KEYINPUT78), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n642), .A2(G80), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G93), .A2(n638), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G55), .A2(n643), .ZN(n616) );
  XNOR2_X1 U695 ( .A(KEYINPUT79), .B(n616), .ZN(n617) );
  NOR2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n659) );
  NAND2_X1 U698 ( .A1(n995), .A2(G559), .ZN(n656) );
  XNOR2_X1 U699 ( .A(n1001), .B(n656), .ZN(n621) );
  NOR2_X1 U700 ( .A1(G860), .A2(n621), .ZN(n622) );
  XOR2_X1 U701 ( .A(n659), .B(n622), .Z(G145) );
  NAND2_X1 U702 ( .A1(G61), .A2(n639), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n623), .B(KEYINPUT80), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n642), .A2(G73), .ZN(n624) );
  XNOR2_X1 U705 ( .A(n624), .B(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G48), .A2(n643), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G86), .A2(n638), .ZN(n627) );
  XNOR2_X1 U709 ( .A(KEYINPUT81), .B(n627), .ZN(n628) );
  NOR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U712 ( .A1(G49), .A2(n643), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U715 ( .A1(n639), .A2(n634), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n635), .A2(G87), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G85), .A2(n638), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n639), .A2(G60), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G72), .A2(n642), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G47), .A2(n643), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U725 ( .A(KEYINPUT70), .B(n648), .Z(G290) );
  XOR2_X1 U726 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n649) );
  XNOR2_X1 U727 ( .A(G288), .B(n649), .ZN(n650) );
  XNOR2_X1 U728 ( .A(G305), .B(n650), .ZN(n652) );
  XNOR2_X1 U729 ( .A(G290), .B(G166), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n653), .B(G299), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(n659), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(n1001), .ZN(n908) );
  XNOR2_X1 U734 ( .A(n908), .B(n656), .ZN(n657) );
  NOR2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n661) );
  NOR2_X1 U736 ( .A1(G868), .A2(n659), .ZN(n660) );
  NOR2_X1 U737 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U744 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U745 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U746 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U747 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U748 ( .A1(G96), .A2(n668), .ZN(n841) );
  NAND2_X1 U749 ( .A1(n841), .A2(G2106), .ZN(n672) );
  NAND2_X1 U750 ( .A1(G69), .A2(G120), .ZN(n669) );
  NOR2_X1 U751 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U752 ( .A1(G108), .A2(n670), .ZN(n842) );
  NAND2_X1 U753 ( .A1(n842), .A2(G567), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(n843) );
  NOR2_X1 U755 ( .A1(n673), .A2(n843), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n674), .B(KEYINPUT84), .ZN(n840) );
  NAND2_X1 U757 ( .A1(n840), .A2(G36), .ZN(n675) );
  XOR2_X1 U758 ( .A(KEYINPUT85), .B(n675), .Z(G176) );
  NAND2_X1 U759 ( .A1(G102), .A2(n884), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G138), .A2(n885), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U762 ( .A1(G114), .A2(n888), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G126), .A2(n889), .ZN(n678) );
  NAND2_X1 U764 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n681), .A2(n680), .ZN(G164) );
  XNOR2_X1 U766 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n836) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n720) );
  AND2_X1 U768 ( .A1(G40), .A2(n682), .ZN(n684) );
  AND2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U770 ( .A1(n686), .A2(n685), .ZN(n721) );
  NOR2_X1 U771 ( .A1(n720), .A2(n721), .ZN(n831) );
  NAND2_X1 U772 ( .A1(G104), .A2(n884), .ZN(n688) );
  NAND2_X1 U773 ( .A1(G140), .A2(n885), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT34), .B(n689), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G116), .A2(n888), .ZN(n691) );
  NAND2_X1 U777 ( .A1(G128), .A2(n889), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U779 ( .A(KEYINPUT87), .B(n692), .ZN(n693) );
  XNOR2_X1 U780 ( .A(KEYINPUT35), .B(n693), .ZN(n694) );
  NOR2_X1 U781 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U782 ( .A(n696), .B(KEYINPUT36), .ZN(n697) );
  XNOR2_X1 U783 ( .A(n697), .B(KEYINPUT88), .ZN(n898) );
  XNOR2_X1 U784 ( .A(G2067), .B(KEYINPUT37), .ZN(n698) );
  XNOR2_X1 U785 ( .A(n698), .B(KEYINPUT86), .ZN(n829) );
  NOR2_X1 U786 ( .A1(n898), .A2(n829), .ZN(n940) );
  NAND2_X1 U787 ( .A1(n831), .A2(n940), .ZN(n827) );
  NAND2_X1 U788 ( .A1(G95), .A2(n884), .ZN(n700) );
  NAND2_X1 U789 ( .A1(G107), .A2(n888), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n705) );
  NAND2_X1 U791 ( .A1(G119), .A2(n889), .ZN(n701) );
  XOR2_X1 U792 ( .A(KEYINPUT89), .B(n701), .Z(n703) );
  NAND2_X1 U793 ( .A1(n885), .A2(G131), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  OR2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n902) );
  AND2_X1 U796 ( .A1(n902), .A2(G1991), .ZN(n715) );
  NAND2_X1 U797 ( .A1(G141), .A2(n885), .ZN(n706) );
  XNOR2_X1 U798 ( .A(n706), .B(KEYINPUT90), .ZN(n713) );
  NAND2_X1 U799 ( .A1(G117), .A2(n888), .ZN(n708) );
  NAND2_X1 U800 ( .A1(G129), .A2(n889), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n884), .A2(G105), .ZN(n709) );
  XOR2_X1 U803 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U804 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n897) );
  AND2_X1 U806 ( .A1(n897), .A2(G1996), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n934) );
  INV_X1 U808 ( .A(n831), .ZN(n716) );
  NOR2_X1 U809 ( .A1(n934), .A2(n716), .ZN(n824) );
  INV_X1 U810 ( .A(n824), .ZN(n717) );
  NAND2_X1 U811 ( .A1(n827), .A2(n717), .ZN(n819) );
  NOR2_X1 U812 ( .A1(G1981), .A2(G305), .ZN(n718) );
  XOR2_X1 U813 ( .A(n718), .B(KEYINPUT24), .Z(n719) );
  XNOR2_X1 U814 ( .A(n719), .B(KEYINPUT91), .ZN(n723) );
  INV_X1 U815 ( .A(n720), .ZN(n722) );
  NAND2_X1 U816 ( .A1(n771), .A2(G8), .ZN(n801) );
  INV_X1 U817 ( .A(n801), .ZN(n803) );
  NAND2_X1 U818 ( .A1(n723), .A2(n803), .ZN(n796) );
  NAND2_X1 U819 ( .A1(G8), .A2(G166), .ZN(n724) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n724), .ZN(n725) );
  XNOR2_X1 U821 ( .A(n725), .B(KEYINPUT105), .ZN(n793) );
  XOR2_X1 U822 ( .A(KEYINPUT92), .B(n771), .Z(n739) );
  NAND2_X1 U823 ( .A1(n739), .A2(G2067), .ZN(n727) );
  NAND2_X1 U824 ( .A1(G1348), .A2(n771), .ZN(n726) );
  NAND2_X1 U825 ( .A1(n727), .A2(n726), .ZN(n734) );
  INV_X1 U826 ( .A(G1996), .ZN(n954) );
  NOR2_X1 U827 ( .A1(n771), .A2(n954), .ZN(n728) );
  XOR2_X1 U828 ( .A(n728), .B(KEYINPUT26), .Z(n730) );
  NAND2_X1 U829 ( .A1(n771), .A2(G1341), .ZN(n729) );
  NAND2_X1 U830 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U831 ( .A1(n995), .A2(n735), .ZN(n732) );
  XOR2_X1 U832 ( .A(KEYINPUT95), .B(n732), .Z(n733) );
  NAND2_X1 U833 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U834 ( .A1(n995), .A2(n735), .ZN(n736) );
  XOR2_X1 U835 ( .A(KEYINPUT96), .B(n736), .Z(n737) );
  NAND2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n746) );
  INV_X1 U837 ( .A(n739), .ZN(n754) );
  INV_X1 U838 ( .A(G2072), .ZN(n945) );
  NOR2_X1 U839 ( .A1(n754), .A2(n945), .ZN(n741) );
  XNOR2_X1 U840 ( .A(KEYINPUT94), .B(KEYINPUT27), .ZN(n740) );
  XNOR2_X1 U841 ( .A(n741), .B(n740), .ZN(n743) );
  NAND2_X1 U842 ( .A1(n754), .A2(G1956), .ZN(n742) );
  NAND2_X1 U843 ( .A1(n743), .A2(n742), .ZN(n747) );
  NOR2_X1 U844 ( .A1(G299), .A2(n747), .ZN(n744) );
  XNOR2_X1 U845 ( .A(n744), .B(KEYINPUT97), .ZN(n745) );
  NAND2_X1 U846 ( .A1(n746), .A2(n745), .ZN(n750) );
  NAND2_X1 U847 ( .A1(G299), .A2(n747), .ZN(n748) );
  XNOR2_X1 U848 ( .A(n748), .B(KEYINPUT28), .ZN(n749) );
  NAND2_X1 U849 ( .A1(n750), .A2(n749), .ZN(n752) );
  NOR2_X1 U850 ( .A1(n753), .A2(G1961), .ZN(n756) );
  XOR2_X1 U851 ( .A(KEYINPUT25), .B(G2078), .Z(n957) );
  NOR2_X1 U852 ( .A1(n957), .A2(n754), .ZN(n755) );
  NOR2_X1 U853 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U854 ( .A(n757), .B(KEYINPUT93), .Z(n765) );
  OR2_X1 U855 ( .A1(n765), .A2(G301), .ZN(n758) );
  NAND2_X1 U856 ( .A1(n759), .A2(n758), .ZN(n784) );
  XNOR2_X1 U857 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n769) );
  NOR2_X1 U858 ( .A1(G1966), .A2(n801), .ZN(n789) );
  NOR2_X1 U859 ( .A1(G2084), .A2(n771), .ZN(n785) );
  NOR2_X1 U860 ( .A1(n789), .A2(n785), .ZN(n760) );
  NAND2_X1 U861 ( .A1(G8), .A2(n760), .ZN(n762) );
  XNOR2_X1 U862 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n761) );
  XNOR2_X1 U863 ( .A(n762), .B(n761), .ZN(n763) );
  NOR2_X1 U864 ( .A1(G168), .A2(n763), .ZN(n764) );
  XNOR2_X1 U865 ( .A(n764), .B(KEYINPUT99), .ZN(n767) );
  NAND2_X1 U866 ( .A1(n765), .A2(G301), .ZN(n766) );
  NAND2_X1 U867 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U868 ( .A(n769), .B(n768), .ZN(n783) );
  NOR2_X1 U869 ( .A1(G1971), .A2(n801), .ZN(n770) );
  XNOR2_X1 U870 ( .A(KEYINPUT101), .B(n770), .ZN(n774) );
  NOR2_X1 U871 ( .A1(G2090), .A2(n771), .ZN(n772) );
  NOR2_X1 U872 ( .A1(G166), .A2(n772), .ZN(n773) );
  NAND2_X1 U873 ( .A1(n774), .A2(n773), .ZN(n776) );
  AND2_X1 U874 ( .A1(n783), .A2(n776), .ZN(n775) );
  NAND2_X1 U875 ( .A1(n784), .A2(n775), .ZN(n780) );
  INV_X1 U876 ( .A(n776), .ZN(n777) );
  OR2_X1 U877 ( .A1(n777), .A2(G286), .ZN(n778) );
  AND2_X1 U878 ( .A1(n778), .A2(G8), .ZN(n779) );
  NAND2_X1 U879 ( .A1(n780), .A2(n779), .ZN(n782) );
  XOR2_X1 U880 ( .A(KEYINPUT32), .B(KEYINPUT102), .Z(n781) );
  XNOR2_X1 U881 ( .A(n782), .B(n781), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U883 ( .A1(G8), .A2(n785), .ZN(n786) );
  NAND2_X1 U884 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U885 ( .A1(n789), .A2(n788), .ZN(n790) );
  INV_X1 U886 ( .A(n800), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n801), .A2(n794), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n817) );
  NOR2_X1 U890 ( .A1(G1971), .A2(G303), .ZN(n797) );
  NOR2_X1 U891 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NOR2_X1 U892 ( .A1(n797), .A2(n983), .ZN(n798) );
  XNOR2_X1 U893 ( .A(n798), .B(KEYINPUT103), .ZN(n799) );
  NOR2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n802) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n809) );
  NAND2_X1 U896 ( .A1(G1976), .A2(G288), .ZN(n982) );
  INV_X1 U897 ( .A(KEYINPUT33), .ZN(n811) );
  NAND2_X1 U898 ( .A1(n803), .A2(n983), .ZN(n804) );
  NOR2_X1 U899 ( .A1(n811), .A2(n804), .ZN(n805) );
  XOR2_X1 U900 ( .A(n805), .B(KEYINPUT104), .Z(n810) );
  AND2_X1 U901 ( .A1(n982), .A2(n810), .ZN(n807) );
  XNOR2_X1 U902 ( .A(G1981), .B(G305), .ZN(n993) );
  INV_X1 U903 ( .A(n993), .ZN(n806) );
  AND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n815) );
  INV_X1 U906 ( .A(n810), .ZN(n812) );
  OR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U908 ( .A1(n993), .A2(n813), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n821) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U913 ( .A1(n990), .A2(n831), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n834) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n897), .ZN(n929) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n902), .ZN(n932) );
  NOR2_X1 U918 ( .A1(n822), .A2(n932), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U920 ( .A1(n929), .A2(n825), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n826), .B(KEYINPUT39), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n898), .A2(n829), .ZN(n942) );
  NAND2_X1 U924 ( .A1(n830), .A2(n942), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U927 ( .A(n836), .B(n835), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U930 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U932 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  INV_X1 U939 ( .A(n843), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2474), .B(G1981), .Z(n845) );
  XNOR2_X1 U941 ( .A(G1961), .B(G1966), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U943 ( .A(n846), .B(KEYINPUT109), .Z(n848) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U946 ( .A(G1976), .B(G1956), .Z(n850) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1971), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U950 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(G229) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2090), .B(G2678), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(n857), .B(KEYINPUT108), .Z(n859) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2100), .Z(n861) );
  XNOR2_X1 U959 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(G227) );
  NAND2_X1 U962 ( .A1(n888), .A2(G112), .ZN(n864) );
  XOR2_X1 U963 ( .A(KEYINPUT111), .B(n864), .Z(n866) );
  NAND2_X1 U964 ( .A1(n884), .A2(G100), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U966 ( .A(KEYINPUT112), .B(n867), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G124), .A2(n889), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n885), .A2(G136), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n883) );
  NAND2_X1 U973 ( .A1(G106), .A2(n884), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G142), .A2(n885), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n875), .B(KEYINPUT45), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G118), .A2(n888), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G130), .A2(n889), .ZN(n878) );
  XNOR2_X1 U980 ( .A(KEYINPUT113), .B(n878), .ZN(n879) );
  NOR2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U982 ( .A(G164), .B(n881), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n896) );
  NAND2_X1 U984 ( .A1(G103), .A2(n884), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G139), .A2(n885), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n895) );
  NAND2_X1 U987 ( .A1(G115), .A2(n888), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G127), .A2(n889), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  XNOR2_X1 U991 ( .A(KEYINPUT114), .B(n893), .ZN(n894) );
  NOR2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n944) );
  XOR2_X1 U993 ( .A(n896), .B(n944), .Z(n900) );
  XOR2_X1 U994 ( .A(n898), .B(n897), .Z(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U996 ( .A(n901), .B(n931), .Z(n904) );
  XOR2_X1 U997 ( .A(n902), .B(G162), .Z(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U999 ( .A(G160), .B(n905), .Z(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(n907) );
  XOR2_X1 U1001 ( .A(KEYINPUT115), .B(n907), .Z(G395) );
  XOR2_X1 U1002 ( .A(n908), .B(n995), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G286), .B(G171), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n911), .ZN(G397) );
  XOR2_X1 U1006 ( .A(KEYINPUT107), .B(G2451), .Z(n913) );
  XNOR2_X1 U1007 ( .A(G2446), .B(G2427), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n920) );
  XOR2_X1 U1009 ( .A(G2438), .B(G2435), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2430), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1012 ( .A(n916), .B(G2454), .Z(n918) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n920), .B(n919), .ZN(n921) );
  NAND2_X1 U1016 ( .A1(n921), .A2(G14), .ZN(n927) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G108), .ZN(G238) );
  INV_X1 U1025 ( .A(n927), .ZN(G401) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1028 ( .A(KEYINPUT51), .B(n930), .Z(n938) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n936) );
  XOR2_X1 U1031 ( .A(G160), .B(G2084), .Z(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(n941), .B(KEYINPUT116), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n950) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n947) );
  XNOR2_X1 U1038 ( .A(n945), .B(n944), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1040 ( .A(KEYINPUT50), .B(n948), .Z(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n976), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n953), .A2(G29), .ZN(n1037) );
  XNOR2_X1 U1046 ( .A(G32), .B(n954), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n955), .A2(G28), .ZN(n967) );
  XNOR2_X1 U1048 ( .A(G25), .B(G1991), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(n956), .B(KEYINPUT117), .ZN(n965) );
  XNOR2_X1 U1050 ( .A(n957), .B(G27), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(n958), .B(KEYINPUT118), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(G33), .B(G2072), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT119), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n969), .B(n968), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(G35), .B(G2090), .ZN(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1063 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n976), .B(n975), .ZN(n978) );
  INV_X1 U1067 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n979), .ZN(n1035) );
  INV_X1 U1070 ( .A(G16), .ZN(n1031) );
  XNOR2_X1 U1071 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n1031), .B(n980), .ZN(n1007) );
  XOR2_X1 U1073 ( .A(G1956), .B(G299), .Z(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(n983), .B(KEYINPUT123), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G166), .B(G1971), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(KEYINPUT124), .B(n988), .Z(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1081 ( .A(KEYINPUT125), .B(n991), .Z(n1005) );
  XOR2_X1 U1082 ( .A(G1966), .B(G168), .Z(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1084 ( .A(KEYINPUT57), .B(n994), .Z(n1000) );
  XOR2_X1 U1085 ( .A(G1348), .B(n995), .Z(n996) );
  XNOR2_X1 U1086 ( .A(KEYINPUT122), .B(n996), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G1961), .B(G301), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G1341), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1033) );
  XOR2_X1 U1094 ( .A(G1348), .B(KEYINPUT59), .Z(n1008) );
  XNOR2_X1 U1095 ( .A(G4), .B(n1008), .ZN(n1016) );
  XOR2_X1 U1096 ( .A(G1956), .B(G20), .Z(n1011) );
  XOR2_X1 U1097 ( .A(G19), .B(KEYINPUT126), .Z(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(G1341), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G6), .B(G1981), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1014), .B(KEYINPUT127), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1017), .ZN(n1026) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G21), .ZN(n1024) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XOR2_X1 U1109 ( .A(G1986), .B(G24), .Z(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(G5), .B(G1961), .ZN(n1027) );
  NOR2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1038), .Z(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

