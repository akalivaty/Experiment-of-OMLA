//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT67), .A3(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(KEYINPUT68), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n199), .B2(KEYINPUT69), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(G116), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G119), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n189), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(KEYINPUT69), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n201), .A3(G119), .ZN(new_n206));
  INV_X1    g020(.A(new_n189), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n195), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT70), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(KEYINPUT70), .A3(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT64), .A2(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT64), .A2(G146), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT65), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT0), .B(G128), .Z(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT64), .A2(G146), .ZN(new_n222));
  AOI21_X1  g036(.A(G143), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT65), .B1(new_n220), .B2(G143), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n217), .B(new_n218), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(G143), .A3(new_n222), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n214), .A2(G146), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(KEYINPUT0), .A3(G128), .A4(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  INV_X1    g045(.A(G134), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G137), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT11), .A3(G134), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(G137), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n233), .A2(new_n235), .A3(new_n239), .A4(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n230), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n227), .A2(new_n243), .A3(G128), .A4(new_n228), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n217), .B1(new_n223), .B2(new_n225), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n227), .B2(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT66), .B1(new_n232), .B2(G137), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n234), .A3(G134), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n251), .A3(new_n236), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G131), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n253), .A2(new_n240), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n242), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n188), .B1(new_n213), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(G237), .A2(G953), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT27), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n262), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n248), .A2(new_n270), .A3(new_n254), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n271), .A3(new_n242), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n272), .B2(new_n213), .ZN(new_n273));
  INV_X1    g087(.A(new_n212), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT70), .B1(new_n204), .B2(new_n208), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n241), .A2(new_n229), .A3(new_n226), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n253), .A2(new_n240), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n215), .A2(new_n216), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n224), .B1(new_n279), .B2(G143), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n243), .B1(new_n279), .B2(G143), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n280), .B(new_n217), .C1(new_n281), .C2(new_n246), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n282), .B2(new_n244), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n277), .B1(new_n283), .B2(new_n270), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n276), .A2(new_n284), .A3(new_n285), .A4(new_n269), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n273), .A2(new_n286), .B1(new_n213), .B2(new_n272), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n257), .B(new_n268), .C1(new_n287), .C2(new_n188), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n242), .A2(new_n271), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n270), .B1(new_n248), .B2(new_n254), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT30), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n242), .A2(new_n292), .A3(new_n255), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n213), .A2(new_n294), .B1(new_n273), .B2(new_n286), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n267), .B1(new_n295), .B2(new_n265), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n273), .A2(KEYINPUT28), .A3(new_n286), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n265), .B(KEYINPUT73), .Z(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n213), .A2(new_n256), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n257), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n297), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n187), .B(new_n288), .C1(new_n296), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G472), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n299), .B1(new_n297), .B2(new_n301), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT31), .B1(new_n295), .B2(new_n265), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n273), .A2(new_n286), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n292), .B1(new_n284), .B2(new_n269), .ZN(new_n309));
  INV_X1    g123(.A(new_n293), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n213), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AND4_X1   g125(.A1(KEYINPUT31), .A2(new_n308), .A3(new_n311), .A4(new_n265), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n306), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT32), .B1(new_n315), .B2(KEYINPUT74), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n311), .A3(new_n265), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT31), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n308), .A2(new_n311), .A3(KEYINPUT31), .A4(new_n265), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n305), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n314), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT74), .B(KEYINPUT32), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n304), .B1(new_n316), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT78), .A4(G125), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(G125), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n220), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n327), .A2(G146), .A3(new_n330), .A4(new_n333), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n193), .A2(G128), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n337), .A2(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n193), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(KEYINPUT75), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT24), .B(G110), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n335), .A2(new_n336), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n337), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n339), .C1(new_n337), .C2(new_n347), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G110), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n344), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI22_X1  g169(.A1(new_n341), .A2(new_n343), .B1(new_n350), .B2(G110), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n279), .A2(new_n326), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n336), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  INV_X1    g174(.A(G953), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n361), .A2(G221), .A3(G234), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n360), .B(new_n362), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n355), .A2(new_n358), .A3(new_n363), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n187), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(G234), .B2(new_n187), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n366), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n371), .A2(G902), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n369), .A2(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(G221), .B1(new_n376), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT82), .B1(new_n378), .B2(G104), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G107), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n379), .B(new_n382), .C1(new_n381), .C2(G107), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G101), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT81), .B(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(G107), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n378), .A3(G104), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n384), .B1(new_n383), .B2(G101), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n282), .B(new_n244), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n227), .A2(new_n228), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n220), .A2(G143), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n246), .B1(new_n396), .B2(KEYINPUT1), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n244), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n383), .A2(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT83), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n398), .A2(new_n400), .A3(new_n385), .A4(new_n391), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n241), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT12), .B1(new_n241), .B2(KEYINPUT84), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n404), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n241), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(KEYINPUT86), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n406), .B1(new_n402), .B2(new_n241), .ZN(new_n410));
  INV_X1    g224(.A(new_n241), .ZN(new_n411));
  AOI211_X1 g225(.A(new_n411), .B(new_n404), .C1(new_n394), .C2(new_n401), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT10), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n401), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n392), .A2(new_n393), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT10), .A3(new_n248), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n391), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n388), .A2(new_n390), .A3(new_n387), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G101), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(KEYINPUT80), .B2(new_n418), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n418), .A2(KEYINPUT80), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(G101), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n230), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n415), .A2(new_n417), .A3(new_n426), .A4(new_n411), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G140), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT79), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n361), .A2(G227), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n408), .A2(new_n413), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n431), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n415), .A2(new_n417), .A3(new_n426), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n435), .A2(new_n241), .ZN(new_n436));
  INV_X1    g250(.A(new_n427), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n187), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n187), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n410), .A2(new_n412), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT85), .B1(new_n445), .B2(new_n437), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT85), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(new_n427), .C1(new_n410), .C2(new_n412), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n431), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n427), .A2(new_n431), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n436), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n449), .A2(new_n440), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n377), .B1(new_n444), .B2(new_n452), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n376), .A2(new_n370), .A3(G953), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n214), .B2(G128), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n246), .A2(KEYINPUT89), .A3(G143), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n214), .A2(G128), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G134), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT88), .B(G122), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G116), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n202), .A2(G122), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n378), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n461), .A2(new_n232), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n466), .A2(KEYINPUT14), .B1(G116), .B2(new_n464), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n202), .A2(new_n471), .A3(G122), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n378), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n232), .B1(new_n459), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n462), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n476), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n465), .A2(new_n466), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G107), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n477), .A2(new_n478), .B1(new_n480), .B2(new_n467), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n455), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n468), .A2(new_n467), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n470), .A2(new_n472), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n463), .B(new_n483), .C1(new_n484), .C2(new_n378), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n467), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n462), .A2(new_n476), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n462), .A2(new_n476), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n489), .A3(new_n454), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n482), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n491), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G237), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n361), .A3(G214), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n214), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n258), .A2(G143), .A3(G214), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G131), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n239), .A3(new_n499), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n326), .A2(KEYINPUT19), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n326), .A2(KEYINPUT19), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n279), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n336), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(KEYINPUT18), .A3(G131), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n357), .B1(new_n220), .B2(new_n326), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT18), .A2(G131), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n498), .A2(new_n499), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(G113), .B(G122), .Z(new_n514));
  XOR2_X1   g328(.A(KEYINPUT87), .B(G104), .Z(new_n515));
  XOR2_X1   g329(.A(new_n514), .B(new_n515), .Z(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n501), .A2(new_n518), .A3(new_n502), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n500), .A2(KEYINPUT17), .A3(G131), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n335), .A4(new_n336), .ZN(new_n521));
  INV_X1    g335(.A(new_n516), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n512), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  NOR2_X1   g339(.A1(G475), .A2(G902), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n525), .B1(new_n524), .B2(new_n526), .ZN(new_n528));
  INV_X1    g342(.A(G475), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n521), .A2(new_n512), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n516), .ZN(new_n531));
  AOI21_X1  g345(.A(G902), .B1(new_n531), .B2(new_n523), .ZN(new_n532));
  OAI22_X1  g346(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n495), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n361), .A2(G952), .ZN(new_n535));
  INV_X1    g349(.A(G234), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n496), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT21), .B(G898), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT90), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n187), .B(new_n361), .C1(G234), .C2(G237), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G214), .B1(G237), .B2(G902), .ZN(new_n545));
  XNOR2_X1  g359(.A(G110), .B(G122), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n211), .B2(new_n212), .ZN(new_n549));
  INV_X1    g363(.A(G113), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n191), .A2(G119), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT5), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n205), .A2(new_n206), .A3(new_n195), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(new_n552), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n416), .A2(new_n208), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n547), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n425), .B1(new_n274), .B2(new_n275), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n556), .A3(new_n546), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(KEYINPUT6), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT6), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n547), .C1(new_n549), .C2(new_n557), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n230), .A2(G125), .ZN(new_n564));
  INV_X1    g378(.A(G125), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n248), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G224), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G953), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n567), .B(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n561), .A2(new_n563), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n567), .B1(new_n573), .B2(new_n569), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n564), .A2(KEYINPUT7), .A3(new_n566), .A4(new_n570), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n555), .A2(new_n208), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n400), .A2(new_n385), .A3(new_n391), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n556), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n546), .B(KEYINPUT8), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n574), .A2(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n581), .B2(new_n560), .ZN(new_n582));
  OAI21_X1  g396(.A(G210), .B1(G237), .B2(G902), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n572), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n572), .B2(new_n582), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n545), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n453), .A2(new_n544), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n325), .A2(new_n375), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(new_n386), .Z(G3));
  OAI21_X1  g403(.A(G472), .B1(new_n321), .B2(G902), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n315), .A3(new_n375), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n545), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n572), .A2(new_n582), .ZN(new_n594));
  INV_X1    g408(.A(new_n583), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n572), .A2(new_n582), .A3(new_n583), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n542), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n474), .A2(new_n481), .A3(new_n455), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n454), .B1(new_n485), .B2(new_n489), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT33), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n482), .A2(new_n490), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(G478), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n492), .A2(new_n187), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n491), .B2(new_n492), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n524), .A2(new_n526), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT20), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n611));
  INV_X1    g425(.A(new_n532), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(G475), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n599), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n377), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n433), .B2(new_n438), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n442), .B1(new_n618), .B2(new_n440), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n405), .A2(new_n407), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n447), .B1(new_n620), .B2(new_n427), .ZN(new_n621));
  INV_X1    g435(.A(new_n448), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n434), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n451), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(G469), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n617), .B1(new_n619), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n592), .A2(new_n616), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  NAND2_X1  g443(.A1(new_n495), .A2(new_n613), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n543), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT91), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n626), .A2(new_n598), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n632), .A2(new_n633), .A3(new_n591), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NAND2_X1  g450(.A1(new_n590), .A2(new_n315), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n359), .B(new_n638), .Z(new_n639));
  INV_X1    g453(.A(new_n374), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n369), .B2(new_n371), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n587), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  INV_X1    g460(.A(KEYINPUT93), .ZN(new_n647));
  INV_X1    g461(.A(new_n633), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n537), .B(KEYINPUT92), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(new_n540), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n642), .A2(new_n630), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n325), .A2(new_n647), .A3(new_n648), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n304), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT32), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n321), .A2(new_n322), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT74), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n655), .B1(new_n659), .B2(new_n323), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n653), .A2(new_n626), .A3(new_n598), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT93), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XOR2_X1   g478(.A(new_n652), .B(KEYINPUT39), .Z(new_n665));
  AND2_X1   g479(.A1(new_n626), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT40), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n659), .A2(new_n323), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n317), .B1(new_n299), .B2(new_n287), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n187), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G472), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n596), .A2(new_n597), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n369), .A2(new_n371), .ZN(new_n676));
  INV_X1    g490(.A(new_n641), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n495), .A2(new_n533), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n678), .A2(new_n593), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n667), .A2(new_n672), .A3(new_n675), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT95), .B(G143), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G45));
  INV_X1    g497(.A(new_n652), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n614), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT96), .B1(new_n586), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT96), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n608), .A2(new_n613), .A3(new_n652), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n598), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n453), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n325), .A2(new_n690), .A3(new_n678), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT97), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT97), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n325), .A2(new_n690), .A3(new_n693), .A4(new_n678), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  INV_X1    g510(.A(KEYINPUT99), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n618), .B2(new_n440), .ZN(new_n698));
  OAI21_X1  g512(.A(G469), .B1(new_n618), .B2(KEYINPUT98), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n435), .A2(new_n241), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n431), .B1(new_n700), .B2(new_n427), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n450), .B1(new_n445), .B2(KEYINPUT86), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n701), .B1(new_n702), .B2(new_n413), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT98), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n703), .A2(new_n704), .A3(G902), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n698), .B1(new_n699), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n704), .B1(new_n703), .B2(G902), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n618), .A2(KEYINPUT98), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n697), .A4(G469), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n617), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n325), .A2(new_n375), .A3(new_n616), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND2_X1  g527(.A1(new_n706), .A2(new_n709), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n598), .A3(new_n377), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n660), .ZN(new_n716));
  INV_X1    g530(.A(new_n375), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n632), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NOR2_X1   g534(.A1(new_n544), .A2(new_n642), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  NOR2_X1   g537(.A1(new_n599), .A2(new_n679), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n257), .B1(new_n287), .B2(new_n188), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT100), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT100), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n727), .B(new_n257), .C1(new_n287), .C2(new_n188), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n298), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n319), .A2(new_n320), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n322), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(G472), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n313), .B2(new_n187), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n710), .A2(new_n724), .A3(new_n375), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NAND2_X1  g550(.A1(new_n729), .A2(new_n730), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n314), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n590), .A3(new_n678), .A4(new_n688), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n715), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n565), .ZN(G27));
  NAND3_X1  g555(.A1(new_n596), .A2(new_n545), .A3(new_n597), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n453), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n325), .A2(new_n375), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n742), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n626), .A2(new_n746), .A3(new_n614), .A4(new_n684), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n656), .B1(new_n321), .B2(new_n322), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n314), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n304), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n375), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT101), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT101), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n753), .A3(new_n375), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n747), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n745), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n239), .ZN(G33));
  NOR2_X1   g572(.A1(new_n630), .A2(new_n652), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n325), .A2(new_n375), .A3(new_n759), .A4(new_n743), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n449), .B2(new_n451), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n623), .A2(KEYINPUT45), .A3(new_n624), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(G469), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n443), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n443), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n441), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n377), .A3(new_n665), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT102), .ZN(new_n772));
  INV_X1    g586(.A(new_n441), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n766), .B2(new_n767), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n617), .B1(new_n774), .B2(new_n769), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT102), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n665), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT43), .B1(new_n608), .B2(new_n533), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n613), .A2(new_n780), .A3(new_n605), .A4(new_n607), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT103), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n678), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n782), .B1(new_n779), .B2(new_n781), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n637), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT104), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n746), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n637), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n788), .B1(new_n787), .B2(new_n746), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n778), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  INV_X1    g611(.A(KEYINPUT105), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n770), .A2(new_n377), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n798), .B1(new_n799), .B2(KEYINPUT47), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n775), .A2(KEYINPUT105), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT106), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n804), .A3(KEYINPUT47), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT106), .B1(new_n775), .B2(new_n801), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n325), .A2(new_n375), .A3(new_n685), .A4(new_n742), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n803), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  XOR2_X1   g624(.A(new_n714), .B(KEYINPUT49), .Z(new_n811));
  NOR2_X1   g625(.A1(new_n608), .A2(new_n533), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n375), .A2(new_n545), .A3(new_n377), .A4(new_n812), .ZN(new_n813));
  OR4_X1    g627(.A1(new_n672), .A2(new_n811), .A3(new_n675), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n710), .A2(new_n593), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(KEYINPUT112), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n779), .A2(new_n781), .A3(new_n650), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n734), .A2(new_n375), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n816), .A2(new_n675), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(KEYINPUT112), .B2(new_n815), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT50), .Z(new_n822));
  AOI22_X1  g636(.A1(new_n803), .A2(new_n807), .B1(new_n617), .B2(new_n714), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n823), .A2(new_n742), .A3(new_n819), .ZN(new_n824));
  INV_X1    g638(.A(new_n672), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n710), .A2(new_n746), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n717), .A2(new_n537), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n533), .B1(new_n605), .B2(new_n607), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n826), .A2(new_n818), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n299), .B1(new_n725), .B2(KEYINPUT100), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n832), .A2(new_n728), .B1(new_n319), .B2(new_n320), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n590), .B(new_n678), .C1(new_n833), .C2(new_n322), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n829), .A2(new_n830), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n822), .A2(new_n824), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n822), .A2(new_n824), .A3(KEYINPUT113), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(KEYINPUT51), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(KEYINPUT51), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n837), .ZN(new_n842));
  OAI221_X1 g656(.A(new_n535), .B1(new_n819), .B2(new_n715), .C1(new_n828), .C2(new_n615), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT114), .Z(new_n844));
  NAND2_X1  g658(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n750), .A2(new_n753), .A3(new_n375), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n753), .B1(new_n750), .B2(new_n375), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n831), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n848), .B(new_n849), .Z(new_n850));
  NAND4_X1  g664(.A1(new_n840), .A2(new_n842), .A3(new_n844), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n586), .B(new_n617), .C1(new_n706), .C2(new_n709), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n853), .B(new_n325), .C1(new_n718), .C2(new_n721), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n633), .A2(new_n591), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n855), .A2(new_n631), .B1(new_n587), .B2(new_n643), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n856), .A3(new_n711), .A4(new_n735), .ZN(new_n857));
  INV_X1    g671(.A(new_n599), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n614), .B(KEYINPUT107), .Z(new_n859));
  NAND4_X1  g673(.A1(new_n592), .A2(new_n626), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n588), .A2(KEYINPUT108), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT108), .B1(new_n588), .B2(new_n860), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n857), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n740), .B1(new_n654), .B2(new_n662), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  INV_X1    g679(.A(new_n679), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n598), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n642), .A2(new_n684), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT110), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n672), .A2(new_n626), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n695), .A2(new_n864), .A3(new_n865), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n747), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(KEYINPUT109), .A3(new_n835), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT109), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n747), .B2(new_n834), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n453), .A2(new_n534), .A3(new_n652), .A4(new_n742), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n325), .A3(new_n678), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n760), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n757), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n863), .A2(new_n872), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n695), .A2(new_n864), .A3(new_n871), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n883), .A2(KEYINPUT52), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n852), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n856), .A2(new_n711), .A3(new_n735), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n588), .A2(new_n860), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT108), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n588), .A2(KEYINPUT108), .A3(new_n860), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n886), .A2(new_n889), .A3(new_n890), .A4(new_n854), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n760), .A2(new_n879), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n873), .B1(new_n846), .B2(new_n847), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT42), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n892), .A2(new_n894), .A3(new_n745), .A4(new_n877), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n883), .A2(KEYINPUT52), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(KEYINPUT53), .A3(new_n897), .A4(new_n872), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n885), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(KEYINPUT111), .A3(KEYINPUT54), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT111), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n885), .A2(new_n898), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n851), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(G952), .A2(G953), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n814), .B1(new_n906), .B2(new_n907), .ZN(G75));
  NOR2_X1   g722(.A1(new_n361), .A2(G952), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n187), .B1(new_n885), .B2(new_n898), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT56), .B1(new_n911), .B2(G210), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n561), .A2(new_n563), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n571), .ZN(new_n914));
  XNOR2_X1  g728(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT117), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n914), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n910), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n911), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n911), .A2(new_n919), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n595), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n917), .B(KEYINPUT119), .Z(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(KEYINPUT56), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n918), .B1(new_n923), .B2(new_n925), .ZN(G51));
  INV_X1    g740(.A(new_n765), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n920), .A2(new_n927), .A3(new_n921), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(KEYINPUT120), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n901), .A2(new_n904), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n442), .B(KEYINPUT57), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n703), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(KEYINPUT120), .B2(new_n928), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n909), .B1(new_n929), .B2(new_n933), .ZN(G54));
  NAND2_X1  g748(.A1(KEYINPUT58), .A2(G475), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n922), .A2(new_n524), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n524), .B1(new_n922), .B2(new_n936), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n909), .ZN(G60));
  XNOR2_X1  g753(.A(new_n606), .B(KEYINPUT59), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n905), .A2(new_n900), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n602), .A2(new_n604), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n940), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n909), .B1(new_n930), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n944), .A2(KEYINPUT121), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT60), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n885), .B2(new_n898), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n910), .B1(new_n954), .B2(new_n373), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n957));
  INV_X1    g771(.A(new_n954), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n956), .B(new_n957), .C1(new_n639), .C2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT61), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n639), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT123), .B1(new_n962), .B2(new_n955), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n959), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(G66));
  INV_X1    g780(.A(new_n539), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n967), .B2(new_n568), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n863), .B2(G953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n913), .B1(G898), .B2(new_n361), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  XNOR2_X1  g785(.A(new_n294), .B(KEYINPUT124), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n504), .A2(new_n505), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n630), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n666), .B(new_n746), .C1(new_n975), .C2(new_n859), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n976), .A2(new_n660), .A3(new_n717), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n778), .B2(new_n795), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n809), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n681), .A2(new_n695), .A3(new_n864), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n974), .B1(new_n984), .B2(G953), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n361), .B1(G227), .B2(G900), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n695), .A2(new_n864), .ZN(new_n988));
  INV_X1    g802(.A(new_n760), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n988), .A2(new_n757), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n867), .B1(new_n752), .B2(new_n754), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n778), .B1(new_n795), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n990), .A2(new_n809), .A3(new_n992), .A4(new_n361), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n974), .B1(G900), .B2(G953), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n985), .A2(new_n987), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n993), .A2(KEYINPUT125), .A3(new_n994), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n985), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n1000), .A2(new_n1001), .A3(new_n986), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n1000), .B2(new_n986), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n996), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g820(.A(KEYINPUT127), .B(new_n996), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(G72));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  XNOR2_X1  g824(.A(new_n295), .B(new_n265), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n899), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n984), .A2(new_n863), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(new_n265), .A3(new_n1010), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n990), .A2(new_n809), .A3(new_n863), .A4(new_n992), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n266), .A2(new_n1010), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g831(.A(new_n909), .B(new_n1012), .C1(new_n1014), .C2(new_n1017), .ZN(G57));
endmodule


