//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OR3_X1    g0008(.A1(new_n208), .A2(KEYINPUT64), .A3(G13), .ZN(new_n209));
  OAI21_X1  g0009(.A(KEYINPUT64), .B1(new_n208), .B2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G250), .B1(G257), .B2(G264), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n206), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n214), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n222), .B1(KEYINPUT0), .B2(new_n214), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G238), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n229), .B1(new_n217), .B2(new_n230), .C1(new_n218), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n208), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n223), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n230), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n215), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT66), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n206), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT66), .B1(G20), .B2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n206), .A2(G33), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n261), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n252), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(KEYINPUT68), .B(new_n252), .C1(new_n260), .C2(new_n262), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(KEYINPUT11), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(KEYINPUT11), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G68), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT12), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n272), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  INV_X1    g0077(.A(new_n270), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n252), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n205), .A2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G68), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n268), .A2(new_n269), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT65), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n286), .B(new_n205), .C1(G41), .C2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G1), .A3(G13), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n231), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n290), .A2(G274), .ZN(new_n293));
  INV_X1    g0093(.A(new_n284), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G226), .A2(G1698), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n230), .B2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n254), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n297), .A2(new_n301), .B1(G33), .B2(G97), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n302), .B2(new_n290), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT13), .B1(new_n292), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n290), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n308), .B1(new_n285), .B2(new_n287), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G238), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n309), .A2(new_n310), .A3(new_n295), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(G169), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n314), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n315), .B1(new_n314), .B2(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n283), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n269), .A2(new_n282), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n314), .A2(G200), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n304), .A2(G190), .A3(new_n313), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n268), .A4(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n279), .A2(G50), .A3(new_n280), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n329), .A2(new_n261), .B1(new_n206), .B2(new_n201), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G150), .B2(new_n257), .ZN(new_n331));
  INV_X1    g0131(.A(new_n252), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n328), .B1(G50), .B2(new_n270), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G222), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G223), .A2(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n301), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n308), .C1(G77), .C2(new_n301), .ZN(new_n338));
  INV_X1    g0138(.A(G226), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n338), .B(new_n295), .C1(new_n339), .C2(new_n291), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n333), .B(new_n342), .C1(G179), .C2(new_n340), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT67), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(KEYINPUT67), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G238), .A2(G1698), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n301), .B(new_n348), .C1(new_n230), .C2(G1698), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n308), .C1(G107), .C2(new_n301), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n295), .C1(new_n225), .C2(new_n291), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n341), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G20), .A2(G77), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n353), .B1(new_n261), .B2(new_n354), .C1(new_n258), .C2(new_n329), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n355), .A2(new_n252), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n279), .A2(G77), .A3(new_n280), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G77), .B2(new_n270), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n352), .B1(G179), .B2(new_n351), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n356), .A2(new_n358), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n351), .A2(G200), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n361), .C1(new_n362), .C2(new_n351), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n347), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G200), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n339), .B2(G1698), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n301), .B1(G33), .B2(G87), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n295), .B1(new_n369), .B2(new_n290), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n288), .A2(G232), .A3(new_n290), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n301), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n308), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n311), .A2(G232), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n362), .A4(new_n295), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n299), .A2(new_n206), .A3(new_n300), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n299), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n300), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n218), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT71), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT71), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(G58), .A3(G68), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n389), .A3(new_n219), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n257), .A2(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n380), .B1(new_n385), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(KEYINPUT3), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT3), .A2(G33), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n382), .A3(new_n206), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n381), .A2(KEYINPUT7), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(G68), .ZN(new_n400));
  AOI22_X1  g0200(.A1(G20), .A2(new_n390), .B1(new_n257), .B2(G159), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n394), .A2(new_n252), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n329), .B1(new_n205), .B2(G20), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(new_n279), .B1(new_n278), .B2(new_n329), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n379), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT17), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n402), .A2(new_n252), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n395), .A2(new_n396), .A3(G20), .ZN(new_n410));
  XOR2_X1   g0210(.A(KEYINPUT70), .B(KEYINPUT7), .Z(new_n411));
  OAI21_X1  g0211(.A(new_n384), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G68), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT16), .B1(new_n413), .B2(new_n401), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n405), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(G169), .B1(new_n370), .B2(new_n371), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n376), .A2(new_n377), .A3(G179), .A4(new_n295), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n403), .A2(new_n405), .B1(new_n416), .B2(new_n417), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT72), .B1(new_n422), .B2(KEYINPUT18), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT72), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n419), .A2(new_n424), .A3(new_n420), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n408), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT9), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n333), .B(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n340), .A2(G200), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n362), .B2(new_n340), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT10), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n333), .B(KEYINPUT9), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT10), .ZN(new_n434));
  INV_X1    g0234(.A(new_n431), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n327), .A2(new_n365), .A3(new_n427), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT75), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n231), .A2(G1698), .ZN(new_n440));
  AND2_X1   g0240(.A1(G244), .A2(G1698), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n440), .A2(new_n441), .B1(new_n395), .B2(new_n396), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G116), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n308), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n227), .B1(new_n446), .B2(G1), .ZN(new_n447));
  INV_X1    g0247(.A(G274), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n205), .A2(new_n448), .A3(G45), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n290), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(G169), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n290), .B1(new_n442), .B2(new_n443), .ZN(new_n452));
  INV_X1    g0252(.A(new_n450), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n452), .A2(G179), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n439), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT19), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n206), .B1(new_n306), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n226), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT76), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n218), .A2(G20), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n206), .A2(G33), .A3(G97), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n301), .A2(new_n463), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT76), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n457), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n252), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n354), .A2(new_n278), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n205), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n270), .A2(new_n471), .A3(new_n215), .A4(new_n251), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n354), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n469), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G244), .A2(G1698), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n231), .B2(G1698), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n301), .A2(new_n478), .B1(G33), .B2(G116), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n317), .B(new_n450), .C1(new_n479), .C2(new_n290), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n452), .A2(new_n453), .ZN(new_n481));
  OAI211_X1 g0281(.A(KEYINPUT75), .B(new_n480), .C1(new_n481), .C2(G169), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n455), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n445), .A2(new_n450), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G200), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n468), .A2(new_n252), .B1(new_n278), .B2(new_n354), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n473), .A2(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(G190), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G1698), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(G244), .C1(new_n396), .C2(new_n395), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n225), .B1(new_n299), .B2(new_n300), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n493), .B(new_n494), .C1(new_n495), .C2(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g0296(.A(G250), .B1(new_n395), .B2(new_n396), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n334), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n308), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G41), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n205), .B(G45), .C1(new_n500), .C2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(G41), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n293), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(G41), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n506), .A2(new_n507), .A3(new_n205), .A4(G45), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G257), .A3(new_n290), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n499), .A2(new_n511), .A3(G179), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n495), .A2(new_n492), .B1(G33), .B2(G283), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n491), .B1(new_n397), .B2(new_n225), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n491), .B1(new_n301), .B2(G250), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n334), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n516), .B2(new_n308), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n512), .B1(new_n517), .B2(new_n341), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n412), .A2(G107), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n202), .B1(new_n255), .B2(new_n256), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  AND2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT73), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n525), .A2(new_n459), .A3(KEYINPUT6), .A4(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(KEYINPUT6), .A2(G97), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT73), .B1(new_n527), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n520), .B1(new_n529), .B2(G20), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n332), .B1(new_n519), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n270), .A2(G97), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n473), .B2(G97), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n518), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT74), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n531), .B2(new_n534), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n529), .A2(G20), .ZN(new_n540));
  INV_X1    g0340(.A(new_n520), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n459), .B1(new_n383), .B2(new_n384), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n252), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(KEYINPUT74), .A3(new_n533), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n517), .A2(G200), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n499), .A2(new_n511), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G190), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n539), .B(new_n545), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n490), .A2(new_n537), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G257), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(new_n334), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n301), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G250), .B(new_n334), .C1(new_n395), .C2(new_n396), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G294), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n308), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT82), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n508), .A2(G264), .A3(new_n290), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n505), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(KEYINPUT82), .A3(new_n308), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G169), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(G179), .A3(new_n557), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n226), .A2(G20), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n301), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g0369(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n570), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n572), .A2(KEYINPUT79), .A3(new_n301), .A4(new_n568), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(KEYINPUT22), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(new_n459), .A3(G20), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n576), .B(new_n578), .C1(G20), .C2(new_n443), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT80), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT24), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n332), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT25), .ZN(new_n587));
  AOI211_X1 g0387(.A(G107), .B(new_n270), .C1(KEYINPUT81), .C2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(KEYINPUT81), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(G107), .B2(new_n473), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n566), .B1(new_n586), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n494), .B(new_n206), .C1(G33), .C2(new_n458), .ZN(new_n595));
  INV_X1    g0395(.A(G116), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G20), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n252), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n595), .A2(KEYINPUT20), .A3(new_n252), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n278), .A2(new_n596), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n472), .B2(new_n596), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G179), .ZN(new_n607));
  INV_X1    g0407(.A(G303), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n397), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G264), .A2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n551), .B2(G1698), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(new_n308), .C1(new_n397), .C2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G270), .B(new_n290), .C1(new_n501), .C2(new_n503), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT77), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT77), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n508), .A2(new_n615), .A3(G270), .A4(new_n290), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n612), .A2(new_n614), .A3(new_n505), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n607), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n606), .A2(new_n617), .A3(G169), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT21), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n604), .B1(new_n601), .B2(new_n600), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n341), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(new_n617), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n618), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n606), .B1(G200), .B2(new_n617), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n362), .B2(new_n617), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n575), .A2(new_n581), .A3(new_n584), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n584), .B1(new_n575), .B2(new_n581), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n252), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n559), .A2(new_n362), .A3(new_n561), .A4(new_n562), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n561), .A2(new_n557), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n366), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n630), .A2(new_n592), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n594), .A2(new_n625), .A3(new_n627), .A4(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n438), .A2(new_n550), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT83), .ZN(G372));
  XNOR2_X1  g0438(.A(new_n422), .B(KEYINPUT18), .ZN(new_n639));
  INV_X1    g0439(.A(new_n359), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n321), .B1(new_n325), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n639), .B1(new_n641), .B2(new_n408), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT87), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n437), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n432), .A2(KEYINPUT87), .A3(new_n436), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n347), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n547), .A2(G169), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n545), .A2(new_n539), .B1(new_n648), .B2(new_n512), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT84), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n450), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n290), .A2(new_n447), .A3(new_n449), .A4(KEYINPUT84), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n651), .B(new_n652), .C1(new_n479), .C2(new_n290), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n341), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n654), .A2(KEYINPUT85), .A3(new_n480), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT85), .B1(new_n654), .B2(new_n480), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n476), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n653), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n488), .B1(new_n658), .B2(new_n366), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n469), .A2(new_n470), .A3(new_n487), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n649), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT86), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n535), .B1(new_n648), .B2(new_n512), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n490), .A2(new_n666), .A3(KEYINPUT26), .A4(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n483), .A2(new_n518), .A3(new_n536), .A4(new_n489), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT86), .B1(new_n669), .B2(new_n664), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n665), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT85), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n444), .A2(new_n308), .B1(new_n650), .B2(new_n450), .ZN(new_n673));
  AOI21_X1  g0473(.A(G169), .B1(new_n673), .B2(new_n652), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n674), .B2(new_n454), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n654), .A2(KEYINPUT85), .A3(new_n480), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n661), .B1(new_n677), .B2(new_n476), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(new_n537), .A3(new_n549), .A4(new_n635), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n630), .A2(new_n592), .B1(new_n564), .B2(new_n565), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n620), .A2(new_n624), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n607), .A2(new_n617), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n657), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n671), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n647), .B1(new_n438), .B2(new_n686), .ZN(G369));
  NAND3_X1  g0487(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n621), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n683), .A2(KEYINPUT88), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT88), .ZN(new_n697));
  INV_X1    g0497(.A(new_n695), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n625), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n625), .A2(new_n627), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n696), .B(new_n699), .C1(new_n700), .C2(new_n695), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n630), .A2(new_n592), .A3(new_n634), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n680), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n693), .B1(new_n586), .B2(new_n593), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n594), .B2(new_n694), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n625), .A2(new_n693), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT90), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n709), .A2(new_n712), .B1(new_n680), .B2(new_n694), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(G399));
  NOR2_X1   g0514(.A1(new_n212), .A2(G41), .ZN(new_n715));
  NOR4_X1   g0515(.A1(new_n715), .A2(new_n205), .A3(G116), .A4(new_n460), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n221), .B2(new_n715), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT28), .Z(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n686), .B2(new_n693), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n549), .A2(new_n537), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n594), .A2(new_n625), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n635), .A4(new_n678), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n665), .A2(new_n668), .A3(new_n670), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(new_n657), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(KEYINPUT94), .A3(new_n694), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n720), .A2(new_n721), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(KEYINPUT26), .B2(new_n669), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n694), .B1(new_n685), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n550), .ZN(new_n735));
  INV_X1    g0535(.A(new_n700), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n706), .A4(new_n694), .ZN(new_n737));
  XNOR2_X1  g0537(.A(KEYINPUT92), .B(KEYINPUT30), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n612), .A2(G179), .A3(new_n560), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n614), .A2(new_n505), .A3(new_n616), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(new_n481), .A4(new_n557), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT91), .B1(new_n741), .B2(new_n547), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n481), .A2(new_n557), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n612), .A2(G179), .A3(new_n560), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT91), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n517), .A3(new_n746), .A4(new_n740), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n738), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n517), .A3(new_n740), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n658), .A2(KEYINPUT93), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT93), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n653), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n751), .A2(new_n632), .A3(new_n753), .A4(new_n317), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n547), .A2(new_n617), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n749), .A2(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n693), .B1(new_n748), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(KEYINPUT31), .B(new_n693), .C1(new_n748), .C2(new_n756), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n737), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G330), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n734), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n718), .B1(new_n764), .B2(G1), .ZN(G364));
  AND2_X1   g0565(.A1(new_n206), .A2(G13), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n205), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n715), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n704), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G330), .B2(new_n702), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n215), .B1(G20), .B2(new_n341), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n206), .A2(new_n317), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n775), .A2(new_n366), .A3(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G179), .A2(G200), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n206), .B1(new_n777), .B2(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n776), .A2(G68), .B1(G97), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT97), .Z(new_n781));
  NAND3_X1  g0581(.A1(new_n777), .A2(G20), .A3(new_n362), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G159), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT32), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n774), .A2(G190), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n366), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n301), .B1(new_n791), .B2(new_n259), .C1(new_n202), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n789), .A2(G200), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n206), .A2(new_n366), .A3(G179), .A4(G190), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n795), .A2(G58), .B1(G107), .B2(new_n796), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n206), .A2(new_n362), .A3(new_n366), .A4(G179), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n797), .B1(new_n226), .B2(new_n799), .ZN(new_n800));
  OR4_X1    g0600(.A1(new_n781), .A2(new_n788), .A3(new_n794), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n776), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  INV_X1    g0603(.A(new_n795), .ZN(new_n804));
  INV_X1    g0604(.A(G322), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  INV_X1    g0607(.A(G326), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n791), .A2(new_n808), .B1(new_n778), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G283), .B2(new_n796), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n397), .B1(new_n608), .B2(new_n799), .C1(new_n793), .C2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G329), .B2(new_n786), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n807), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n773), .B1(new_n801), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n211), .A2(G355), .A3(new_n301), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(G116), .B2(new_n211), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n212), .A2(new_n301), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n446), .B2(new_n221), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n246), .A2(G45), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G13), .A2(G33), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(G20), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n772), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n769), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n830), .A2(KEYINPUT95), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(KEYINPUT95), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n816), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n826), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n702), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n771), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NOR2_X1   g0638(.A1(new_n364), .A2(new_n693), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n671), .B2(new_n685), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n720), .A2(new_n728), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n363), .B1(new_n360), .B2(new_n694), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n359), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n359), .A2(new_n693), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n840), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n769), .B1(new_n848), .B2(new_n762), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n762), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n772), .A2(new_n824), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n833), .B1(new_n202), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G150), .A2(new_n776), .B1(new_n792), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  INV_X1    g0654(.A(G143), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n854), .B2(new_n791), .C1(new_n855), .C2(new_n804), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT34), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n301), .B1(new_n778), .B2(new_n217), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n798), .A2(G50), .B1(new_n796), .B2(G68), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT100), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n858), .B(new_n860), .C1(G132), .C2(new_n786), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n397), .B1(new_n793), .B2(new_n596), .C1(new_n862), .C2(new_n802), .ZN(new_n863));
  INV_X1    g0663(.A(new_n796), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n226), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n791), .A2(new_n608), .B1(new_n459), .B2(new_n799), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n785), .A2(new_n812), .ZN(new_n867));
  NOR4_X1   g0667(.A1(new_n863), .A2(new_n865), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n795), .A2(G294), .B1(G97), .B2(new_n779), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT99), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n857), .A2(new_n861), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n852), .B1(new_n773), .B2(new_n871), .C1(new_n847), .C2(new_n825), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n850), .A2(new_n872), .ZN(G384));
  OR2_X1    g0673(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n874), .A2(G116), .A3(new_n216), .A4(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT36), .Z(new_n877));
  NAND4_X1  g0677(.A1(new_n221), .A2(G77), .A3(new_n389), .A4(new_n387), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n259), .A2(G68), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n205), .B(G13), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT16), .B1(new_n400), .B2(new_n401), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n405), .B1(new_n409), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n691), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n408), .B2(new_n426), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n419), .A2(new_n888), .A3(new_n406), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n415), .A2(new_n884), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n415), .A2(KEYINPUT102), .A3(new_n884), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n405), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n402), .A2(new_n252), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n394), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n897), .A2(new_n379), .B1(new_n883), .B2(new_n884), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n883), .A2(new_n418), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n888), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT103), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n894), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n892), .A2(new_n893), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n419), .A2(new_n888), .A3(new_n406), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n885), .A2(new_n899), .A3(new_n406), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT37), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT103), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(KEYINPUT38), .B(new_n887), .C1(new_n902), .C2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n901), .B1(new_n894), .B2(new_n900), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(KEYINPUT103), .A3(new_n907), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n913), .B2(new_n887), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT39), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n903), .A2(new_n406), .A3(new_n419), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n894), .B1(new_n917), .B2(KEYINPUT37), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n903), .B1(new_n407), .B2(new_n639), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n909), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n321), .A2(new_n694), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n283), .A2(new_n693), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n320), .A2(new_n325), .A3(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n283), .B(new_n693), .C1(new_n318), .C2(new_n319), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n840), .B2(new_n845), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT101), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n844), .B1(new_n727), .B2(new_n839), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT101), .B1(new_n935), .B2(new_n931), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n934), .B(new_n936), .C1(new_n910), .C2(new_n914), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n639), .A2(new_n884), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n926), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n438), .B1(new_n729), .B2(new_n733), .ZN(new_n941));
  INV_X1    g0741(.A(new_n647), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n940), .B(new_n943), .Z(new_n944));
  AOI21_X1  g0744(.A(new_n846), .B1(new_n928), .B2(new_n929), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n761), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n910), .B2(new_n914), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n909), .A2(new_n920), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n761), .A2(new_n945), .A3(KEYINPUT40), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n947), .A2(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n438), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(new_n761), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n953), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(G330), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n944), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n205), .B2(new_n766), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n944), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n881), .B1(new_n958), .B2(new_n959), .ZN(G367));
  OAI21_X1  g0760(.A(new_n827), .B1(new_n211), .B2(new_n354), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n819), .B2(new_n242), .ZN(new_n962));
  INV_X1    g0762(.A(G159), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n301), .B1(new_n802), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G50), .B2(new_n792), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n791), .A2(new_n855), .B1(new_n217), .B2(new_n799), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G77), .B2(new_n796), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n786), .A2(G137), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n795), .A2(G150), .B1(G68), .B2(new_n779), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n965), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT46), .B1(new_n798), .B2(G116), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n397), .B1(new_n793), .B2(new_n862), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(G294), .C2(new_n776), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n798), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  INV_X1    g0774(.A(G317), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n973), .B(new_n974), .C1(new_n975), .C2(new_n785), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n864), .A2(new_n458), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G303), .B2(new_n795), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n459), .B2(new_n778), .C1(new_n812), .C2(new_n791), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n970), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n833), .B(new_n962), .C1(new_n981), .C2(new_n772), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT111), .Z(new_n983));
  NAND3_X1  g0783(.A1(new_n657), .A2(new_n660), .A3(new_n693), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n694), .B1(new_n486), .B2(new_n487), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n678), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT105), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n983), .B1(new_n835), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n703), .B(new_n709), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(new_n712), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n764), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n649), .A2(new_n693), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n545), .A2(new_n539), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n693), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n994), .B1(new_n722), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n713), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n713), .A2(new_n998), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n710), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n993), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n764), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n715), .B(KEYINPUT41), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n768), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n709), .A2(new_n712), .A3(new_n998), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT42), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n667), .B1(new_n998), .B2(new_n680), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n693), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT106), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT106), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1011), .A2(KEYINPUT42), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT107), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT108), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1021), .B1(KEYINPUT109), .B2(new_n1022), .ZN(new_n1023));
  AND4_X1   g0823(.A1(new_n1005), .A2(new_n1019), .A3(new_n1023), .A4(new_n998), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1019), .A2(new_n1023), .B1(new_n1005), .B2(new_n998), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1022), .A2(KEYINPUT109), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n989), .B1(new_n1010), .B2(new_n1028), .ZN(G387));
  OR2_X1    g0829(.A1(new_n709), .A2(new_n835), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n239), .A2(G45), .A3(new_n397), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n460), .A2(G116), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n446), .B1(new_n218), .B2(new_n202), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n329), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1034), .A2(KEYINPUT50), .A3(new_n259), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT50), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n329), .B2(G50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1033), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1032), .B1(new_n1038), .B2(new_n301), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n212), .B1(new_n1031), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n827), .B1(new_n211), .B2(new_n459), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n301), .B1(new_n793), .B2(new_n218), .C1(new_n329), .C2(new_n802), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G150), .B2(new_n786), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n795), .A2(G50), .B1(new_n474), .B2(new_n779), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT112), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n799), .A2(new_n202), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n977), .B(new_n1047), .C1(new_n790), .C2(G159), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n798), .A2(G294), .B1(new_n779), .B2(G283), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G303), .A2(new_n792), .B1(new_n776), .B2(G311), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n975), .B2(new_n804), .C1(new_n805), .C2(new_n791), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT113), .Z(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(KEYINPUT49), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n301), .B1(new_n796), .B2(G116), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n808), .C2(new_n785), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT49), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n833), .B(new_n1042), .C1(new_n1061), .C2(new_n772), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n992), .A2(new_n768), .B1(new_n1030), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n993), .A2(new_n715), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n992), .A2(new_n764), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(G393));
  NOR2_X1   g0866(.A1(new_n820), .A2(new_n249), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n828), .B(new_n1067), .C1(G97), .C2(new_n212), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G150), .A2(new_n790), .B1(new_n795), .B2(G159), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT51), .Z(new_n1070));
  NOR2_X1   g0870(.A1(new_n778), .A2(new_n202), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1071), .B(new_n865), .C1(G68), .C2(new_n798), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n786), .A2(G143), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n301), .B1(new_n802), .B2(new_n259), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1034), .B2(new_n792), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G311), .A2(new_n795), .B1(new_n790), .B2(G317), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT52), .Z(new_n1078));
  OAI22_X1  g0878(.A1(new_n802), .A2(new_n608), .B1(new_n778), .B2(new_n596), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1079), .A2(KEYINPUT115), .B1(G294), .B2(new_n792), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(KEYINPUT115), .C2(new_n1079), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n301), .B1(new_n796), .B2(G107), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n862), .B2(new_n799), .C1(new_n785), .C2(new_n805), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT114), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1076), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n833), .B(new_n1068), .C1(new_n772), .C2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n998), .B2(new_n835), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1007), .A2(new_n715), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n993), .A2(new_n1006), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1087), .B1(new_n767), .B2(new_n1006), .C1(new_n1088), .C2(new_n1089), .ZN(G390));
  OAI21_X1  g0890(.A(KEYINPUT116), .B1(new_n932), .B2(new_n925), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT116), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n924), .C1(new_n935), .C2(new_n931), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1091), .A2(new_n915), .A3(new_n922), .A4(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n761), .A2(G330), .A3(new_n847), .A4(new_n930), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n694), .B(new_n843), .C1(new_n685), .C2(new_n731), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1096), .A2(new_n845), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n924), .B(new_n949), .C1(new_n1097), .C2(new_n931), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1094), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1095), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n768), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n833), .B1(new_n329), .B2(new_n851), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n864), .A2(new_n259), .B1(new_n963), .B2(new_n778), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n301), .B1(new_n793), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(G137), .C2(new_n776), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G128), .A2(new_n790), .B1(new_n795), .B2(G132), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT119), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n798), .A2(G150), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT53), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n786), .A2(G125), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n791), .A2(new_n862), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1071), .B(new_n1114), .C1(G116), .C2(new_n795), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n397), .B1(new_n793), .B2(new_n458), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G107), .B2(new_n776), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n786), .A2(G294), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n798), .A2(G87), .B1(new_n796), .B2(G68), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1113), .A2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1103), .B1(new_n773), .B2(new_n1121), .C1(new_n923), .C2(new_n825), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1102), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n759), .A2(new_n760), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n636), .A2(new_n550), .A3(new_n693), .ZN(new_n1125));
  OAI211_X1 g0925(.A(G330), .B(new_n847), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n931), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n1097), .A3(new_n1095), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT118), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT118), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(new_n1097), .A3(new_n1130), .A4(new_n1095), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1126), .A2(new_n1134), .A3(new_n931), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1095), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n935), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n762), .A2(new_n438), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n941), .A2(new_n1140), .A3(new_n942), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1100), .B2(new_n1099), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1095), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1094), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1146), .A2(new_n1147), .A3(new_n1141), .A4(new_n1139), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n715), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1123), .A2(new_n1149), .ZN(G378));
  AOI21_X1  g0950(.A(new_n830), .B1(new_n259), .B2(new_n851), .ZN(new_n1151));
  INV_X1    g0951(.A(G132), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n802), .A2(new_n1152), .B1(new_n793), .B2(new_n854), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n790), .A2(G125), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n795), .A2(G128), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n799), .C2(new_n1105), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1153), .B(new_n1156), .C1(G150), .C2(new_n779), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G33), .B(G41), .C1(new_n796), .C2(G159), .ZN(new_n1161));
  INV_X1    g0961(.A(G124), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n785), .B2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT120), .Z(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G41), .B(new_n301), .C1(new_n792), .C2(new_n474), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n458), .B2(new_n802), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1047), .B(new_n1167), .C1(G68), .C2(new_n779), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n862), .B2(new_n785), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n864), .A2(new_n217), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n804), .A2(new_n459), .B1(new_n791), .B2(new_n596), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1172), .A2(KEYINPUT58), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(KEYINPUT58), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n259), .B1(new_n395), .B2(G41), .ZN(new_n1175));
  AND4_X1   g0975(.A1(new_n1165), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n333), .A2(new_n884), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT55), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n646), .A2(new_n343), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n646), .B2(new_n343), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1178), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n646), .A2(new_n343), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1180), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n646), .A2(new_n343), .A3(new_n1180), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1177), .A3(new_n1187), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1183), .A2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1151), .B1(new_n773), .B2(new_n1176), .C1(new_n1189), .C2(new_n825), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1183), .A2(new_n1188), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n951), .B2(G330), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n950), .A2(new_n949), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n761), .A2(new_n945), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n887), .B1(new_n902), .B2(new_n908), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT38), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1194), .B1(new_n1197), .B2(new_n909), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G330), .B(new_n1193), .C1(new_n1198), .C2(KEYINPUT40), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(new_n1189), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n940), .B1(new_n1192), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1189), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n947), .A2(new_n948), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1203), .A2(new_n1191), .A3(G330), .A4(new_n1193), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n938), .B1(new_n923), .B2(new_n925), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n937), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1190), .B1(new_n1207), .B2(new_n767), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n715), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1201), .A2(KEYINPUT57), .A3(new_n1206), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1148), .A2(new_n1141), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1210), .B1(new_n1213), .B2(KEYINPUT122), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT122), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT123), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1140), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n647), .B(new_n1218), .C1(new_n734), .C2(new_n438), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1101), .B2(new_n1139), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1201), .A2(new_n1206), .A3(KEYINPUT57), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT122), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1222), .A2(new_n1216), .A3(KEYINPUT123), .A4(new_n715), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1220), .B2(new_n1207), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1209), .B1(new_n1217), .B2(new_n1226), .ZN(G375));
  NAND3_X1  g1027(.A1(new_n1219), .A2(new_n1138), .A3(new_n1132), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1142), .A3(new_n1009), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n930), .A2(new_n825), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT124), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n397), .B1(new_n793), .B2(new_n459), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G116), .B2(new_n776), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n791), .A2(new_n809), .B1(new_n458), .B2(new_n799), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G283), .B2(new_n795), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n786), .A2(G303), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n779), .A2(new_n474), .B1(new_n796), .B2(G77), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1233), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n791), .A2(new_n1152), .B1(new_n778), .B2(new_n259), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G137), .B2(new_n795), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n786), .A2(G128), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n792), .A2(G150), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n301), .C1(new_n802), .C2(new_n1105), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1170), .B1(G159), .B2(new_n798), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1240), .A2(new_n1241), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n773), .B1(new_n1238), .B2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1247), .B(new_n833), .C1(new_n218), .C2(new_n851), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1139), .A2(new_n768), .B1(new_n1231), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1229), .A2(new_n1249), .ZN(G381));
  OR2_X1    g1050(.A1(G387), .A2(G390), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G378), .A2(new_n1251), .A3(G375), .A4(new_n1252), .ZN(G407));
  INV_X1    g1053(.A(G378), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n692), .A2(G213), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G375), .C2(new_n1257), .ZN(G409));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1228), .A2(KEYINPUT125), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT60), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n715), .B(new_n1142), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1249), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n850), .A3(new_n872), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G384), .B(new_n1249), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G378), .B(new_n1209), .C1(new_n1217), .C2(new_n1226), .ZN(new_n1268));
  AND4_X1   g1068(.A1(new_n1009), .A2(new_n1212), .A3(new_n1206), .A4(new_n1201), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1254), .B1(new_n1269), .B2(new_n1208), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1256), .B(new_n1267), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1259), .B1(new_n1271), .B2(KEYINPUT127), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1255), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1255), .A2(KEYINPUT126), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1265), .A2(new_n1266), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1256), .A2(G2897), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1276), .B(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT61), .B1(new_n1274), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1267), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1273), .A2(new_n1255), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT127), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(KEYINPUT62), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1272), .A2(new_n1279), .A3(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(G393), .B(G396), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G387), .A2(G390), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1251), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1285), .B1(new_n1251), .B2(new_n1286), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1271), .A2(KEYINPUT63), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1271), .A2(KEYINPUT63), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .A4(new_n1279), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1290), .A2(new_n1294), .ZN(G405));
  XNOR2_X1  g1095(.A(G375), .B(G378), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1296), .A2(new_n1267), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1267), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1292), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1289), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(G402));
endmodule


