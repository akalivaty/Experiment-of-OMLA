//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT27), .Z(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  OR3_X1    g011(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n193), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n197), .B1(new_n200), .B2(new_n196), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n208), .A2(new_n209), .A3(G131), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n208), .B2(G131), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n204), .A2(new_n206), .A3(new_n213), .A4(new_n207), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n201), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n221), .A3(G128), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT69), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n193), .A3(new_n228), .A4(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n219), .B1(new_n225), .B2(new_n226), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n194), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n214), .B(KEYINPUT65), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n203), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n205), .A3(G134), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n238), .A3(new_n207), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n234), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(G116), .B(G119), .Z(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n217), .A2(new_n241), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT28), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n208), .A2(G131), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n208), .A2(new_n209), .A3(G131), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n235), .ZN(new_n254));
  INV_X1    g068(.A(new_n240), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n230), .B2(new_n233), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n254), .A2(new_n201), .B1(new_n256), .B2(new_n235), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n257), .B2(new_n245), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n217), .A2(new_n241), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n244), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n247), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n192), .B(new_n249), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n224), .A2(new_n229), .B1(new_n232), .B2(new_n194), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n216), .A2(new_n266), .A3(new_n255), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n198), .A2(new_n199), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n195), .B1(new_n268), .B2(new_n193), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n253), .A2(new_n235), .B1(new_n197), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT30), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n217), .A2(new_n241), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n247), .B1(new_n274), .B2(new_n244), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n265), .B1(new_n275), .B2(new_n192), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n217), .A2(new_n241), .A3(new_n272), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n272), .B1(new_n217), .B2(new_n241), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n244), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n246), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT72), .A3(new_n191), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n264), .A2(new_n276), .A3(new_n277), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n259), .A2(new_n244), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n246), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n259), .A2(KEYINPUT73), .A3(new_n244), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(KEYINPUT28), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n191), .A2(new_n277), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n249), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G472), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n260), .B1(new_n259), .B2(new_n244), .ZN(new_n297));
  AOI211_X1 g111(.A(KEYINPUT71), .B(new_n245), .C1(new_n217), .C2(new_n241), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n246), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT28), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n192), .B1(new_n300), .B2(new_n249), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n302));
  NAND4_X1  g116(.A1(new_n280), .A2(new_n192), .A3(new_n246), .A4(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n245), .B1(new_n271), .B2(new_n273), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n304), .A2(new_n191), .A3(new_n247), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n295), .B(new_n296), .C1(new_n301), .C2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n280), .A2(new_n192), .A3(new_n246), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT31), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n248), .B1(new_n299), .B2(KEYINPUT28), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n311), .B(new_n303), .C1(new_n312), .C2(new_n192), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n295), .B1(new_n313), .B2(new_n296), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n294), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(G234), .B2(new_n291), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(G125), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT75), .B(G125), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(new_n321), .ZN(new_n324));
  OR2_X1    g138(.A1(KEYINPUT75), .A2(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT75), .A2(G125), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n320), .A3(G140), .A4(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n319), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n323), .A2(new_n319), .A3(new_n321), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G146), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n330), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n218), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G128), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT23), .A3(G119), .ZN(new_n336));
  INV_X1    g150(.A(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G128), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(G128), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n336), .B(new_n338), .C1(new_n339), .C2(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G110), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT24), .B(G110), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n339), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n338), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n341), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n334), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n218), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n344), .A2(new_n345), .B1(new_n347), .B2(new_n338), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n340), .A2(G110), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n328), .A2(new_n218), .A3(new_n332), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G953), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(G221), .A3(G234), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT77), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G137), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n351), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n364), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n349), .B1(new_n331), .B2(new_n333), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(new_n358), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(new_n368), .A3(new_n291), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT25), .A4(new_n291), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n318), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n365), .A2(new_n368), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n317), .A2(G902), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n315), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n315), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G140), .ZN(new_n382));
  INV_X1    g196(.A(G227), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G953), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n382), .B(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G107), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n389), .A2(KEYINPUT3), .A3(G104), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n389), .B2(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT81), .A3(G101), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n394), .B(new_n388), .C1(new_n390), .C2(new_n391), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n392), .A2(KEYINPUT81), .A3(new_n397), .A4(G101), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n201), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n389), .B2(G104), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n389), .A2(G104), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n387), .A2(KEYINPUT82), .A3(G107), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n395), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT10), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n234), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n218), .A2(G143), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT1), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n193), .B2(G128), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n224), .B2(new_n229), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n407), .B1(new_n413), .B2(new_n406), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n399), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT83), .B1(new_n212), .B2(new_n216), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n253), .A2(new_n235), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n386), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT87), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n415), .A2(new_n254), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT87), .B(new_n386), .C1(new_n415), .C2(new_n419), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n415), .A2(new_n419), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n230), .A2(new_n406), .A3(new_n233), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n406), .B2(new_n413), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n429));
  XOR2_X1   g243(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n253), .B2(new_n235), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n429), .B1(new_n428), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n230), .A2(new_n406), .A3(new_n233), .ZN(new_n435));
  INV_X1    g249(.A(new_n412), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n406), .B1(new_n230), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT86), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n427), .B(new_n439), .C1(new_n406), .C2(new_n413), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n254), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT12), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n426), .B1(new_n434), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n385), .B(KEYINPUT80), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n425), .B(G469), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G469), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n420), .B1(new_n434), .B2(new_n443), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n415), .A2(new_n419), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n386), .B1(new_n449), .B2(new_n423), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n447), .B(new_n291), .C1(new_n448), .C2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n447), .A2(new_n291), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n446), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT9), .B(G234), .ZN(new_n455));
  OAI21_X1  g269(.A(G221), .B1(new_n455), .B2(G902), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT79), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT88), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n461), .A3(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n466));
  OAI21_X1  g280(.A(G131), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n468));
  INV_X1    g282(.A(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n360), .A3(G214), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n220), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n213), .A3(new_n464), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n464), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(KEYINPUT17), .A3(G131), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n331), .A2(new_n476), .A3(new_n333), .ZN(new_n477));
  NAND2_X1  g291(.A1(KEYINPUT18), .A2(G131), .ZN(new_n478));
  OR3_X1    g292(.A1(new_n474), .A2(KEYINPUT91), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n474), .B2(KEYINPUT91), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n324), .A2(G146), .A3(new_n327), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(new_n353), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G113), .B(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(new_n387), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT93), .Z(new_n486));
  NAND3_X1  g300(.A1(new_n477), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n328), .A2(new_n332), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n488), .A2(G146), .B1(new_n467), .B2(new_n472), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n324), .A2(KEYINPUT19), .A3(new_n327), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT19), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n352), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n324), .A2(new_n491), .A3(KEYINPUT19), .A4(new_n327), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n218), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n482), .B1(new_n489), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n487), .B1(new_n498), .B2(new_n485), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n500));
  NOR2_X1   g314(.A1(G475), .A2(G902), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT94), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n499), .A2(new_n504), .A3(new_n500), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n499), .A2(new_n501), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT20), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(G234), .A2(G237), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(G952), .A3(new_n360), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT21), .B(G898), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(G902), .A3(G953), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n220), .A2(G128), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n335), .A2(G143), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n203), .ZN(new_n518));
  XNOR2_X1  g332(.A(G116), .B(G122), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n389), .ZN(new_n520));
  INV_X1    g334(.A(G116), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT14), .A3(G122), .ZN(new_n522));
  INV_X1    g336(.A(new_n519), .ZN(new_n523));
  OAI211_X1 g337(.A(G107), .B(new_n522), .C1(new_n523), .C2(KEYINPUT14), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n515), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n526), .A2(KEYINPUT13), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n516), .B1(new_n526), .B2(KEYINPUT13), .ZN(new_n528));
  OAI21_X1  g342(.A(G134), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n517), .A2(new_n203), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n519), .B(new_n389), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n455), .A2(new_n316), .A3(G953), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n525), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n525), .B2(new_n532), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n291), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT15), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(G478), .ZN(new_n538));
  INV_X1    g352(.A(G478), .ZN(new_n539));
  OAI221_X1 g353(.A(new_n291), .B1(KEYINPUT15), .B2(new_n539), .C1(new_n534), .C2(new_n535), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n487), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n485), .B1(new_n477), .B2(new_n483), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n291), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G475), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n508), .A2(new_n514), .A3(new_n541), .A4(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT5), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n337), .A3(G116), .ZN(new_n552));
  OAI211_X1 g366(.A(G113), .B(new_n552), .C1(new_n242), .C2(new_n551), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n242), .A2(new_n243), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n555), .A2(new_n406), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n396), .A2(new_n244), .A3(new_n398), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G122), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT89), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(KEYINPUT6), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n201), .A2(new_n323), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n266), .B2(new_n323), .ZN(new_n566));
  INV_X1    g380(.A(G224), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n565), .B(new_n570), .C1(new_n266), .C2(new_n323), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT6), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n558), .A2(new_n573), .A3(new_n561), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n564), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n568), .A2(KEYINPUT7), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n569), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n560), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n561), .A2(KEYINPUT8), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n555), .A2(new_n406), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n553), .A2(new_n554), .B1(new_n405), .B2(new_n395), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n563), .B(new_n583), .C1(KEYINPUT7), .C2(new_n571), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n291), .B1(new_n577), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n550), .B1(new_n575), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n563), .A2(new_n583), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n571), .A2(KEYINPUT7), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n569), .A2(new_n571), .A3(new_n576), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n564), .A2(new_n572), .A3(new_n574), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n549), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G214), .B1(G237), .B2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT90), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n595), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n586), .B2(new_n593), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT90), .ZN(new_n601));
  AND4_X1   g415(.A1(new_n463), .A2(new_n548), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n381), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n394), .ZN(G3));
  INV_X1    g418(.A(new_n463), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n296), .B1(new_n301), .B2(new_n307), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n313), .B2(new_n291), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n376), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n605), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n508), .A2(new_n545), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n539), .A2(new_n291), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n536), .B2(G478), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n534), .A2(new_n535), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n618), .A2(KEYINPUT33), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(KEYINPUT33), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n621), .B2(G478), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n614), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n600), .A2(new_n514), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n613), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT96), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  INV_X1    g443(.A(new_n541), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n630), .B(new_n545), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n613), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n371), .A2(new_n372), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n317), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n367), .A2(new_n358), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n366), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n375), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n639), .A2(KEYINPUT97), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT97), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n373), .B2(new_n644), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n611), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n602), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT37), .B(G110), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  OAI21_X1  g467(.A(new_n510), .B1(new_n513), .B2(G900), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT98), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n633), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n646), .A2(new_n600), .A3(new_n648), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n463), .A2(new_n315), .A3(new_n656), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XOR2_X1   g474(.A(new_n655), .B(KEYINPUT39), .Z(new_n661));
  AND2_X1   g475(.A1(new_n463), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n606), .A2(KEYINPUT32), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n308), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n286), .A2(new_n191), .A3(new_n287), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(KEYINPUT99), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n310), .B1(new_n668), .B2(KEYINPUT99), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n291), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G472), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n594), .B(KEYINPUT38), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n639), .A2(new_n645), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n675), .A2(new_n541), .A3(new_n599), .ZN(new_n676));
  AND4_X1   g490(.A1(new_n614), .A2(new_n673), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n664), .A2(new_n665), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  INV_X1    g493(.A(new_n655), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n614), .A2(new_n622), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n463), .A2(new_n315), .A3(new_n658), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT100), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n657), .B1(new_n667), .B2(new_n294), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n463), .A4(new_n681), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  OR2_X1    g502(.A1(new_n448), .A2(new_n450), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n291), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(new_n456), .A3(new_n451), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n315), .A2(new_n625), .A3(new_n376), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT41), .B(G113), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  NAND4_X1  g509(.A1(new_n315), .A2(new_n376), .A3(new_n634), .A4(new_n692), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  NAND4_X1  g511(.A1(new_n548), .A2(new_n315), .A3(new_n658), .A4(new_n692), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT101), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  NAND3_X1  g514(.A1(new_n614), .A2(new_n630), .A3(new_n600), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(new_n514), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n192), .B1(new_n288), .B2(new_n249), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n307), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n609), .B1(new_n296), .B2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n706), .A3(new_n376), .A4(new_n692), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  AND4_X1   g522(.A1(new_n456), .A2(new_n691), .A3(new_n451), .A4(new_n600), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n706), .A3(new_n675), .A4(new_n681), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  OAI21_X1  g525(.A(KEYINPUT102), .B1(new_n309), .B2(new_n314), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n666), .A2(new_n713), .A3(new_n308), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n294), .A3(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n586), .A2(new_n595), .A3(new_n593), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n716), .A2(new_n454), .A3(new_n456), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n717), .A2(new_n681), .A3(KEYINPUT42), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(new_n718), .A3(new_n376), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n715), .A2(new_n718), .A3(new_n721), .A4(new_n376), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n315), .A2(new_n376), .A3(new_n681), .A4(new_n717), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n720), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT104), .B(G131), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G33));
  NAND4_X1  g542(.A1(new_n315), .A2(new_n376), .A3(new_n656), .A4(new_n717), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND3_X1  g548(.A1(new_n586), .A2(new_n595), .A3(new_n593), .ZN(new_n735));
  INV_X1    g549(.A(new_n614), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n622), .ZN(new_n737));
  XOR2_X1   g551(.A(new_n737), .B(KEYINPUT43), .Z(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n611), .A3(new_n675), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n740), .B2(new_n739), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n742), .A2(KEYINPUT107), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n425), .B1(new_n444), .B2(new_n445), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n447), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n452), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(KEYINPUT46), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n451), .B1(new_n748), .B2(KEYINPUT46), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n456), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n661), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n742), .A2(KEYINPUT107), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n743), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  OR2_X1    g571(.A1(new_n752), .A2(KEYINPUT47), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n752), .A2(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n681), .A2(new_n612), .A3(new_n716), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n315), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  AND2_X1   g578(.A1(new_n691), .A2(new_n451), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT49), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n622), .A2(new_n458), .A3(new_n595), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n674), .A2(new_n612), .A3(new_n614), .A4(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(new_n667), .A3(new_n672), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n598), .A2(new_n514), .A3(new_n601), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n508), .A2(new_n541), .A3(new_n545), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n736), .B2(new_n622), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n463), .A3(new_n376), .A4(new_n610), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n693), .A2(new_n774), .A3(new_n707), .A4(new_n696), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n602), .B1(new_n381), .B2(new_n650), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n699), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n538), .A2(new_n540), .A3(new_n680), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n545), .B(new_n779), .C1(new_n631), .C2(new_n632), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n778), .B1(new_n716), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n735), .A2(new_n780), .A3(KEYINPUT108), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n782), .A2(new_n649), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n463), .A3(new_n315), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n706), .A2(new_n681), .A3(new_n675), .A4(new_n717), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n731), .B2(new_n732), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n726), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n777), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n680), .A2(new_n456), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n454), .A2(new_n639), .A3(new_n645), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n701), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n673), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n659), .A2(new_n710), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n687), .A2(KEYINPUT110), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT110), .B1(new_n687), .B2(new_n795), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT52), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n687), .A2(new_n795), .A3(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT109), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n687), .A2(new_n795), .A3(new_n801), .A4(KEYINPUT52), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n790), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(KEYINPUT111), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n687), .A2(new_n795), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n687), .A2(new_n795), .A3(KEYINPUT110), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(KEYINPUT53), .B(new_n790), .C1(new_n798), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT111), .B1(new_n804), .B2(new_n805), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT54), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT112), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n737), .B(KEYINPUT43), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n510), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n692), .A2(new_n716), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n819), .A2(new_n675), .A3(new_n706), .A4(new_n821), .ZN(new_n822));
  OR4_X1    g636(.A1(new_n510), .A2(new_n820), .A3(new_n673), .A4(new_n612), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n614), .A2(new_n622), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n706), .A2(new_n376), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(new_n692), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n674), .A2(new_n595), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n819), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n825), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n765), .A2(new_n457), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n758), .A2(new_n759), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n826), .A3(new_n716), .A4(new_n819), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(KEYINPUT51), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT114), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n836), .B1(new_n833), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n715), .A2(new_n376), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n819), .A2(new_n844), .A3(new_n821), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT48), .ZN(new_n846));
  OAI211_X1 g660(.A(G952), .B(new_n360), .C1(new_n823), .C2(new_n623), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n819), .A2(new_n827), .A3(new_n600), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n838), .A2(new_n843), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n804), .A2(new_n805), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n798), .A2(new_n812), .ZN(new_n859));
  INV_X1    g673(.A(new_n790), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n857), .B(new_n858), .C1(KEYINPUT53), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n863), .B(KEYINPUT54), .C1(new_n814), .C2(new_n815), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n817), .A2(new_n856), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n865), .A2(new_n866), .B1(G952), .B2(G953), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n862), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n804), .A2(new_n805), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT111), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n813), .A3(new_n806), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n863), .B1(new_n872), .B2(KEYINPUT54), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT117), .B1(new_n874), .B2(new_n856), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n769), .B1(new_n867), .B2(new_n875), .ZN(G75));
  OAI21_X1  g690(.A(new_n857), .B1(KEYINPUT53), .B2(new_n861), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(G210), .A3(G902), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n564), .A2(new_n574), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT118), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n572), .B(KEYINPUT55), .Z(new_n881));
  XNOR2_X1  g695(.A(new_n880), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT120), .ZN(new_n883));
  XOR2_X1   g697(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n360), .A2(G952), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n877), .A2(G902), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT56), .B1(new_n891), .B2(G210), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n892), .B2(new_n882), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n888), .A2(new_n893), .ZN(G51));
  XNOR2_X1  g708(.A(new_n452), .B(KEYINPUT57), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(new_n862), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n689), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n891), .A2(new_n746), .A3(new_n747), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n889), .B1(new_n899), .B2(new_n900), .ZN(G54));
  NAND3_X1  g715(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n902));
  INV_X1    g716(.A(new_n499), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n904), .A2(new_n905), .A3(new_n889), .ZN(G60));
  INV_X1    g720(.A(new_n621), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n615), .B(KEYINPUT59), .Z(new_n908));
  OAI211_X1 g722(.A(new_n907), .B(new_n908), .C1(new_n896), .C2(new_n897), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n890), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n868), .B2(new_n873), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n621), .B2(new_n911), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT122), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n877), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n374), .B(KEYINPUT123), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n918), .B(new_n890), .C1(new_n642), .C2(new_n916), .ZN(new_n919));
  AND2_X1   g733(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n920));
  NOR2_X1   g734(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n919), .B2(new_n921), .ZN(G66));
  AOI21_X1  g737(.A(new_n360), .B1(new_n512), .B2(G224), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n777), .B2(new_n360), .ZN(new_n925));
  INV_X1    g739(.A(G898), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n880), .B1(new_n926), .B2(G953), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n925), .B(new_n927), .ZN(G69));
  AND3_X1   g742(.A1(new_n687), .A2(new_n659), .A3(new_n710), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n678), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n663), .A2(new_n735), .A3(new_n772), .ZN(new_n933));
  AOI22_X1  g747(.A1(new_n760), .A2(new_n762), .B1(new_n381), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n756), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n360), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n274), .B(new_n496), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT125), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n940));
  INV_X1    g754(.A(G900), .ZN(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n383), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n754), .A2(new_n702), .A3(new_n844), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n756), .A2(new_n943), .A3(new_n726), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n763), .A2(new_n733), .A3(new_n929), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(G953), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(G900), .A2(G953), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n937), .A2(new_n947), .ZN(new_n948));
  OAI221_X1 g762(.A(new_n939), .B1(new_n940), .B2(new_n942), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n942), .A2(new_n940), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G72));
  NOR2_X1   g765(.A1(new_n281), .A2(new_n192), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT127), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n944), .A2(new_n777), .A3(new_n945), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n953), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n935), .B2(new_n777), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n192), .A3(new_n281), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n960), .A3(new_n890), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n276), .A2(new_n282), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n957), .B1(new_n962), .B2(new_n310), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n961), .B1(new_n872), .B2(new_n963), .ZN(G57));
endmodule


