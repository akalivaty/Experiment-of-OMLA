//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  INV_X1    g001(.A(G234), .ZN(new_n188));
  OAI21_X1  g002(.A(G217), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT69), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G902), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(G125), .A2(G140), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n192), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n197), .ZN(new_n201));
  NOR2_X1   g015(.A1(G125), .A2(G140), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT16), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n199), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(G128), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT70), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(KEYINPUT70), .A3(G128), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT24), .B(G110), .Z(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n207), .B2(G128), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT23), .A3(G119), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n209), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT71), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT71), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n219), .A3(new_n222), .A4(new_n209), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G110), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n206), .B(new_n215), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n196), .A2(new_n197), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n192), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n213), .A2(new_n214), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n220), .A2(G110), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n205), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT73), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT73), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G137), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT72), .ZN(new_n237));
  INV_X1    g051(.A(G221), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n238), .A2(new_n188), .A3(G953), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n237), .B(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n233), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n240), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n242), .A2(new_n234), .A3(new_n226), .A4(new_n231), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n191), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n233), .A2(new_n235), .A3(new_n240), .ZN(new_n246));
  AOI21_X1  g060(.A(G902), .B1(new_n246), .B2(new_n243), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT25), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n190), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT74), .B(KEYINPUT25), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  AOI211_X1 g066(.A(G902), .B(new_n252), .C1(new_n246), .C2(new_n243), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n187), .B(new_n245), .C1(new_n250), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G902), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(new_n251), .C1(new_n241), .C2(new_n244), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n257), .B(new_n190), .C1(new_n249), .C2(new_n247), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n187), .B1(new_n258), .B2(new_n245), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(G116), .B(G119), .Z(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT2), .B(G113), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n261), .B(new_n262), .Z(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n192), .A2(G143), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n218), .A2(KEYINPUT0), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n218), .A2(KEYINPUT0), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n268), .B(KEYINPUT64), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  XNOR2_X1  g086(.A(G143), .B(G146), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT0), .B(G128), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT11), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(G137), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(G137), .ZN(new_n280));
  INV_X1    g094(.A(G137), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT11), .A3(G134), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G131), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n279), .A2(new_n282), .A3(new_n285), .A4(new_n280), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n288));
  NAND2_X1  g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n268), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n273), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n276), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n273), .A2(new_n294), .A3(G128), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n266), .B(G146), .C1(new_n218), .C2(KEYINPUT1), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n218), .A2(new_n192), .A3(G143), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n296), .A2(KEYINPUT66), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT66), .B1(new_n296), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n280), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n278), .A2(G137), .ZN(new_n302));
  OAI21_X1  g116(.A(G131), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n303), .A2(new_n286), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT30), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n293), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n293), .B2(new_n305), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n264), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n293), .A2(new_n305), .A3(new_n263), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(G101), .ZN(new_n313));
  NOR2_X1   g127(.A1(G237), .A2(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G210), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n313), .B(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n310), .A2(new_n311), .A3(new_n316), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n293), .A2(new_n305), .A3(new_n263), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n263), .B1(new_n293), .B2(new_n305), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n311), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n316), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n317), .B1(new_n323), .B2(KEYINPUT31), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT67), .B(KEYINPUT31), .Z(new_n325));
  NAND4_X1  g139(.A1(new_n310), .A2(new_n311), .A3(new_n316), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT68), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n293), .A2(new_n305), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT30), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n307), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n318), .B1(new_n330), .B2(new_n264), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n316), .A4(new_n325), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G472), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n256), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n334), .A2(new_n338), .A3(new_n335), .A4(new_n256), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n331), .A2(new_n316), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n320), .A2(new_n316), .A3(new_n322), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n256), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n342), .A2(new_n343), .ZN(new_n346));
  OAI21_X1  g160(.A(G472), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n260), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT96), .ZN(new_n349));
  INV_X1    g163(.A(G478), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(KEYINPUT15), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT95), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT14), .ZN(new_n356));
  INV_X1    g170(.A(G116), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(G122), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(G122), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G122), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G116), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n356), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(G116), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT92), .B(new_n364), .C1(new_n362), .C2(new_n356), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G107), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n266), .A2(G128), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n218), .A2(G143), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n373), .A3(new_n278), .ZN(new_n374));
  OAI21_X1  g188(.A(G134), .B1(new_n370), .B2(new_n372), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n359), .A2(new_n362), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n366), .A2(KEYINPUT93), .A3(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n369), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n383));
  OR3_X1    g197(.A1(new_n372), .A2(new_n383), .A3(KEYINPUT13), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n370), .B1(KEYINPUT13), .B2(new_n372), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n372), .B2(KEYINPUT13), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n377), .B(new_n378), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n374), .A3(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT9), .B(G234), .Z(new_n391));
  INV_X1    g205(.A(G953), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(G217), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n382), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(new_n382), .B2(new_n390), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n256), .B(new_n354), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n352), .A2(new_n353), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n349), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n397), .ZN(new_n401));
  AOI21_X1  g215(.A(G902), .B1(new_n401), .B2(new_n395), .ZN(new_n402));
  INV_X1    g216(.A(new_n399), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n402), .A2(KEYINPUT96), .A3(new_n403), .A4(new_n354), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT94), .B1(new_n402), .B2(new_n352), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n256), .B1(new_n396), .B2(new_n397), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT94), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n351), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G952), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G953), .ZN(new_n412));
  INV_X1    g226(.A(G237), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n188), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n256), .B(new_n392), .C1(G234), .C2(G237), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT21), .B(G898), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n415), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(new_n392), .A3(G214), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT84), .A3(G143), .ZN(new_n422));
  OR2_X1    g236(.A1(KEYINPUT84), .A2(G143), .ZN(new_n423));
  NAND2_X1  g237(.A1(KEYINPUT84), .A2(G143), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n423), .A2(G214), .A3(new_n314), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n285), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT17), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(new_n425), .A3(G131), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT87), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n429), .A2(new_n428), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(new_n206), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n427), .A2(new_n434), .A3(new_n428), .A4(new_n429), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT18), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n426), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n227), .B(new_n192), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n422), .A2(new_n425), .A3(KEYINPUT18), .A4(G131), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n438), .A2(new_n427), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G113), .B(G122), .ZN(new_n443));
  INV_X1    g257(.A(G104), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT90), .ZN(new_n447));
  AOI21_X1  g261(.A(G902), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n442), .B2(new_n447), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G475), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n405), .A2(new_n410), .A3(new_n420), .A4(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n427), .A2(new_n429), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT19), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n227), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n196), .A2(KEYINPUT19), .A3(new_n197), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n192), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n205), .A3(KEYINPUT85), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT85), .B1(new_n458), .B2(new_n205), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n441), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n205), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n454), .A3(new_n459), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT86), .B1(new_n468), .B2(new_n441), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n446), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n436), .A2(new_n445), .A3(new_n441), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n453), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n452), .B(KEYINPUT88), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n463), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n468), .A2(KEYINPUT86), .A3(new_n441), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n445), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n471), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n473), .B(new_n475), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n470), .A2(new_n471), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n473), .A4(new_n475), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n474), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n451), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G214), .B1(G237), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT3), .B1(new_n444), .B2(G107), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT77), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n444), .A2(G107), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n378), .A3(G104), .ZN(new_n494));
  OAI211_X1 g308(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n444), .C2(G107), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n491), .A2(new_n492), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT78), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n494), .A2(new_n492), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n499), .A2(KEYINPUT78), .A3(new_n491), .A4(new_n495), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(G101), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G101), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n499), .A2(new_n502), .A3(new_n491), .A4(new_n495), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n498), .A2(KEYINPUT4), .A3(G101), .A4(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n264), .ZN(new_n508));
  XOR2_X1   g322(.A(G110), .B(G122), .Z(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n492), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n444), .A2(G107), .ZN(new_n512));
  OAI21_X1  g326(.A(G101), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n207), .A3(G116), .ZN(new_n517));
  OAI211_X1 g331(.A(G113), .B(new_n517), .C1(new_n261), .C2(new_n516), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n261), .A2(new_n262), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n508), .A2(new_n510), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n263), .B1(new_n505), .B2(new_n506), .ZN(new_n523));
  INV_X1    g337(.A(new_n521), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n509), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(KEYINPUT6), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n509), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n296), .A2(new_n297), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT66), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n296), .A2(KEYINPUT66), .A3(new_n297), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n531), .A2(new_n532), .B1(new_n273), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n194), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n276), .A2(new_n292), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n537), .B2(new_n194), .ZN(new_n538));
  INV_X1    g352(.A(G224), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G953), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT82), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n538), .B(new_n541), .Z(new_n542));
  NAND3_X1  g356(.A1(new_n526), .A2(new_n528), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n538), .A2(KEYINPUT83), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT83), .B1(new_n538), .B2(new_n544), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n538), .A2(new_n544), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n509), .B(KEYINPUT8), .Z(new_n549));
  NOR2_X1   g363(.A1(new_n515), .A2(new_n520), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n524), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n547), .A2(new_n522), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n543), .A2(new_n256), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G210), .B1(G237), .B2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n543), .A2(new_n256), .A3(new_n552), .A4(new_n554), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n488), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n238), .B1(new_n391), .B2(new_n256), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT79), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n536), .B1(new_n505), .B2(new_n506), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n562), .A2(new_n503), .A3(new_n513), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n563), .A2(KEYINPUT10), .B1(new_n564), .B2(new_n514), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n561), .A2(new_n287), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n514), .A2(new_n534), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n562), .A2(new_n503), .A3(new_n513), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT12), .B1(new_n569), .B2(new_n287), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n571));
  INV_X1    g385(.A(new_n287), .ZN(new_n572));
  AOI211_X1 g386(.A(new_n571), .B(new_n572), .C1(new_n567), .C2(new_n568), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n560), .B1(new_n566), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n572), .B1(new_n567), .B2(new_n568), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT12), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n507), .A2(new_n537), .ZN(new_n578));
  INV_X1    g392(.A(new_n565), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n580), .A3(KEYINPUT79), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G140), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT76), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n392), .A2(G227), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n287), .B1(new_n561), .B2(new_n565), .ZN(new_n587));
  INV_X1    g401(.A(new_n585), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n580), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n589), .A3(G469), .ZN(new_n590));
  INV_X1    g404(.A(G469), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n256), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT80), .B1(new_n566), .B2(new_n585), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT80), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n580), .A2(new_n596), .A3(new_n588), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n597), .A3(new_n577), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT81), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n580), .A2(new_n587), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n585), .ZN(new_n601));
  AOI211_X1 g415(.A(KEYINPUT81), .B(new_n588), .C1(new_n580), .C2(new_n587), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(new_n591), .A3(new_n256), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n559), .B1(new_n594), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n348), .A2(new_n486), .A3(new_n558), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(new_n594), .A2(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n258), .A2(new_n245), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT75), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n254), .ZN(new_n611));
  INV_X1    g425(.A(new_n559), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n608), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n334), .A2(new_n256), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n335), .A2(KEYINPUT97), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT33), .B1(new_n396), .B2(new_n397), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n401), .A2(new_n619), .A3(new_n395), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(G478), .A3(new_n256), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT99), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n350), .B1(new_n618), .B2(new_n620), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n256), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT100), .B1(new_n402), .B2(G478), .ZN(new_n627));
  OR3_X1    g441(.A1(new_n402), .A2(KEYINPUT100), .A3(G478), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n623), .A2(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n481), .A2(new_n484), .ZN(new_n630));
  INV_X1    g444(.A(new_n474), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n630), .A2(new_n631), .B1(G475), .B2(new_n449), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n487), .B1(new_n556), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n556), .A2(new_n634), .A3(new_n557), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n633), .A2(new_n636), .A3(new_n420), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n617), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT34), .B(G104), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  XNOR2_X1  g455(.A(new_n419), .B(KEYINPUT102), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n472), .B2(new_n473), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n478), .A2(new_n479), .ZN(new_n646));
  OAI211_X1 g460(.A(KEYINPUT101), .B(KEYINPUT20), .C1(new_n646), .C2(new_n453), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n482), .A2(new_n473), .A3(new_n452), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n405), .A2(new_n410), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n649), .A2(new_n650), .A3(new_n450), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n636), .A2(new_n637), .A3(new_n643), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT103), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n556), .A2(new_n634), .A3(new_n557), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n635), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n643), .A4(new_n651), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n617), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT35), .B(G107), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NAND4_X1  g474(.A1(new_n605), .A2(new_n486), .A3(new_n616), .A4(new_n558), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n242), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n232), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n191), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n258), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT37), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G110), .ZN(G12));
  NAND2_X1  g483(.A1(new_n340), .A2(new_n347), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n605), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n636), .A2(new_n637), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n671), .A2(new_n672), .A3(new_n666), .ZN(new_n673));
  INV_X1    g487(.A(new_n416), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n414), .B1(new_n674), .B2(G900), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n651), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  INV_X1    g492(.A(new_n331), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n316), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n318), .A2(new_n319), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n256), .B1(new_n683), .B2(new_n316), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n340), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n650), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n632), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n556), .A2(new_n557), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT38), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n487), .A2(new_n687), .A3(new_n689), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n675), .B(KEYINPUT39), .Z(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n605), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n697), .A3(new_n666), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NAND3_X1  g513(.A1(new_n633), .A2(KEYINPUT104), .A3(new_n675), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n630), .A2(new_n631), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n450), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n628), .A2(new_n627), .ZN(new_n703));
  INV_X1    g517(.A(new_n626), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n625), .B1(new_n624), .B2(new_n256), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n702), .A2(new_n706), .A3(new_n675), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n673), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NAND2_X1  g526(.A1(new_n604), .A2(KEYINPUT105), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n591), .B1(new_n603), .B2(new_n256), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI211_X1 g529(.A(KEYINPUT105), .B(new_n591), .C1(new_n603), .C2(new_n256), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n612), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n670), .A2(new_n611), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n717), .A2(new_n638), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT41), .B(G113), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND2_X1  g535(.A1(new_n653), .A2(new_n657), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n603), .A2(new_n256), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(KEYINPUT105), .A3(new_n604), .ZN(new_n725));
  INV_X1    g539(.A(new_n716), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n559), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n722), .A2(new_n348), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  OAI211_X1 g543(.A(new_n655), .B(new_n612), .C1(new_n715), .C2(new_n716), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT106), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n727), .A2(new_n732), .A3(new_n655), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n451), .A2(new_n666), .A3(new_n485), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n731), .A2(new_n733), .A3(new_n670), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  INV_X1    g550(.A(new_n609), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n614), .A2(G472), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n738), .A2(new_n739), .A3(new_n336), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n614), .A2(new_n739), .A3(G472), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT108), .ZN(new_n743));
  INV_X1    g557(.A(new_n741), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n738), .A2(new_n739), .A3(new_n336), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n737), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n730), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n689), .A2(new_n643), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  AOI21_X1  g568(.A(new_n666), .B1(new_n744), .B2(new_n745), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n700), .A2(new_n709), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n731), .A2(new_n756), .A3(new_n733), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  NOR2_X1   g572(.A1(new_n690), .A2(new_n488), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n700), .A2(new_n709), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n670), .A2(new_n737), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n605), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n700), .A2(new_n709), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n670), .A2(new_n611), .A3(new_n605), .A4(new_n759), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G131), .ZN(G33));
  INV_X1    g583(.A(new_n766), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n676), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n278), .ZN(G36));
  NAND2_X1  g586(.A1(new_n586), .A2(new_n589), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n586), .A2(KEYINPUT45), .A3(new_n589), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(G469), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n593), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n593), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n604), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n612), .A3(new_n694), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n759), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n616), .A2(new_n666), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n703), .B(new_n788), .C1(new_n704), .C2(new_n705), .ZN(new_n789));
  NOR2_X1   g603(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n789), .B(new_n632), .C1(new_n629), .C2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n702), .C2(new_n629), .ZN(new_n792));
  OR2_X1    g606(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n787), .A2(new_n791), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n786), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n783), .A2(new_n784), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n785), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  AND3_X1   g614(.A1(new_n782), .A2(KEYINPUT112), .A3(new_n612), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT112), .B1(new_n782), .B2(new_n612), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n801), .A2(new_n802), .B1(KEYINPUT113), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n782), .A2(new_n612), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n808));
  NAND3_X1  g622(.A1(new_n782), .A2(KEYINPUT112), .A3(new_n612), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n765), .A2(new_n670), .A3(new_n786), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n804), .A2(new_n810), .A3(new_n260), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n415), .A2(new_n791), .A3(new_n792), .A4(new_n793), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n749), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT118), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n691), .A2(new_n487), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(new_n727), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n749), .A2(new_n727), .A3(new_n815), .ZN(new_n821));
  INV_X1    g635(.A(new_n819), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT118), .B(new_n817), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n717), .A2(new_n786), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n815), .ZN(new_n826));
  INV_X1    g640(.A(new_n755), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n717), .A2(new_n260), .A3(new_n786), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n686), .A2(new_n415), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n830), .A2(new_n632), .A3(new_n629), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n824), .A2(KEYINPUT117), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n816), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n804), .A2(new_n810), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n725), .A2(new_n726), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n559), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n786), .B(new_n835), .C1(new_n836), .C2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n824), .A2(new_n829), .A3(new_n833), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n814), .B(new_n834), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n833), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n828), .B(new_n842), .C1(new_n820), .C2(new_n823), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n836), .A2(new_n838), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n759), .A3(new_n816), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n843), .B(new_n845), .C1(KEYINPUT117), .C2(KEYINPUT51), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n826), .A2(KEYINPUT119), .A3(new_n761), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n826), .B2(new_n761), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(KEYINPUT48), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n816), .A2(new_n731), .A3(new_n733), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n830), .A2(new_n633), .A3(new_n832), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n412), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n849), .A2(KEYINPUT48), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n673), .B1(new_n710), .B2(new_n676), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n655), .A2(new_n689), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n686), .A2(new_n665), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n605), .A4(new_n675), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n757), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n757), .A2(new_n856), .A3(KEYINPUT52), .A4(new_n859), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n771), .B1(new_n764), .B2(new_n767), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n688), .A2(new_n450), .ZN(new_n866));
  INV_X1    g680(.A(new_n649), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n671), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n665), .A3(new_n675), .A4(new_n759), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n760), .A2(KEYINPUT116), .A3(new_n605), .A4(new_n755), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n700), .A2(new_n709), .A3(new_n605), .A4(new_n759), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n871), .B1(new_n872), .B2(new_n827), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n865), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n719), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n735), .A2(new_n753), .A3(new_n728), .A4(new_n876), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n488), .B(new_n642), .C1(new_n556), .C2(new_n557), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n605), .A2(new_n878), .A3(new_n611), .A4(new_n616), .ZN(new_n879));
  INV_X1    g693(.A(new_n633), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n608), .A2(new_n486), .A3(new_n558), .A4(new_n612), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n879), .A2(new_n880), .B1(new_n718), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n613), .A2(new_n616), .A3(new_n633), .A4(new_n878), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(KEYINPUT115), .A3(new_n606), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n632), .A2(new_n650), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n879), .A2(new_n888), .B1(new_n661), .B2(new_n666), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n877), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n864), .A2(new_n875), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n864), .A2(new_n875), .A3(new_n892), .A4(KEYINPUT53), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(KEYINPUT54), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT54), .B1(new_n895), .B2(new_n896), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n847), .B(new_n855), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n411), .A2(new_n392), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n837), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT49), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n702), .A2(new_n629), .A3(new_n559), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n737), .A3(new_n487), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT114), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n687), .B(new_n691), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OAI221_X1 g722(.A(new_n908), .B1(new_n907), .B2(new_n906), .C1(KEYINPUT49), .C2(new_n903), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n902), .A2(new_n909), .ZN(G75));
  NAND2_X1  g724(.A1(new_n526), .A2(new_n528), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n542), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  INV_X1    g727(.A(G210), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n914), .B(new_n256), .C1(new_n895), .C2(new_n896), .ZN(new_n915));
  NOR2_X1   g729(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n256), .B1(new_n895), .B2(new_n896), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G210), .ZN(new_n920));
  INV_X1    g734(.A(new_n913), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n392), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n918), .A2(new_n922), .A3(new_n924), .ZN(G51));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n889), .B1(new_n884), .B2(new_n886), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n730), .B1(new_n748), .B2(new_n743), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n719), .B1(new_n928), .B2(new_n752), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n927), .A2(new_n929), .A3(new_n728), .A4(new_n735), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n862), .B2(new_n863), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT53), .B1(new_n931), .B2(new_n875), .ZN(new_n932));
  INV_X1    g746(.A(new_n896), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n926), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n592), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n897), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n603), .ZN(new_n938));
  INV_X1    g752(.A(new_n777), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n919), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n923), .B1(new_n938), .B2(new_n940), .ZN(G54));
  NAND3_X1  g755(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n646), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n924), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n646), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(G60));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT59), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n934), .A2(new_n897), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n621), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n934), .A2(new_n621), .A3(new_n897), .A4(new_n948), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n924), .A3(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n932), .B2(new_n933), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n241), .A2(new_n244), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n923), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n663), .B(new_n956), .C1(new_n932), .C2(new_n933), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n959), .B(new_n960), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n961));
  INV_X1    g775(.A(new_n958), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n895), .B2(new_n896), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n960), .B(new_n924), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT61), .B1(new_n960), .B2(KEYINPUT122), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n961), .A2(new_n966), .ZN(G66));
  OAI21_X1  g781(.A(G953), .B1(new_n418), .B2(new_n539), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n892), .B2(G953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n911), .B1(G898), .B2(new_n392), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  AND2_X1   g785(.A1(new_n812), .A2(new_n799), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n757), .A2(new_n856), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(KEYINPUT62), .A3(new_n698), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n698), .A2(new_n757), .A3(new_n856), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n456), .A2(new_n457), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n330), .B(new_n979), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n880), .A2(new_n888), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT123), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n694), .A3(new_n770), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n972), .A2(new_n978), .A3(new_n981), .A4(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n812), .A2(new_n799), .A3(new_n865), .A4(new_n973), .ZN(new_n986));
  INV_X1    g800(.A(new_n761), .ZN(new_n987));
  AND4_X1   g801(.A1(new_n987), .A2(new_n785), .A3(new_n798), .A4(new_n857), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n980), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n985), .A2(new_n989), .A3(new_n392), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n981), .A2(G227), .A3(G900), .ZN(new_n991));
  OAI21_X1  g805(.A(G900), .B1(KEYINPUT124), .B2(G227), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n980), .B(new_n992), .C1(KEYINPUT124), .C2(G900), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(G953), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n990), .A2(new_n994), .ZN(G72));
  NAND4_X1  g809(.A1(new_n972), .A2(new_n978), .A3(new_n892), .A4(new_n984), .ZN(new_n996));
  XNOR2_X1  g810(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n335), .A2(new_n256), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n997), .B(new_n998), .Z(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n681), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1001), .A2(KEYINPUT126), .A3(new_n681), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n679), .A2(new_n316), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT127), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n986), .A2(new_n930), .A3(new_n988), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n999), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1004), .A2(new_n1005), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1006), .A2(new_n1000), .ZN(new_n1011));
  AOI211_X1 g825(.A(new_n681), .B(new_n1011), .C1(new_n895), .C2(new_n896), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1010), .A2(new_n923), .A3(new_n1012), .ZN(G57));
endmodule


