//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT2), .B(G113), .Z(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(KEYINPUT68), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  INV_X1    g007(.A(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n191), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n189), .B2(new_n188), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G143), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(KEYINPUT64), .A3(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n203), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n204), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G137), .ZN(new_n218));
  INV_X1    g032(.A(G137), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT11), .A3(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT66), .A4(new_n221), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n220), .A2(new_n221), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n218), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n218), .A2(new_n220), .A3(new_n229), .A4(new_n221), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n224), .A2(new_n226), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n202), .A2(new_n234), .A3(G128), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n208), .A2(G143), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n205), .A2(KEYINPUT64), .A3(G146), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT64), .B1(new_n205), .B2(G146), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G128), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT67), .B1(new_n211), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n236), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n219), .A2(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n221), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G131), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI22_X1  g068(.A1(new_n215), .A2(new_n233), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT30), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n241), .B1(new_n240), .B2(new_n243), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n211), .A2(KEYINPUT67), .A3(new_n246), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n235), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n230), .A2(new_n232), .B1(G131), .B2(new_n250), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n230), .A2(new_n232), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n224), .A2(G131), .A3(new_n225), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n240), .A2(new_n213), .B1(new_n202), .B2(new_n203), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n201), .B1(new_n256), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n261), .A2(new_n266), .A3(new_n201), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n271));
  NOR2_X1   g085(.A1(G237), .A2(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G210), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n271), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT31), .B1(new_n269), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n248), .A2(new_n254), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n215), .B1(new_n262), .B2(new_n263), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n200), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(new_n283), .B2(new_n270), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n270), .A2(new_n280), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n276), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n282), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n267), .B1(new_n261), .B2(new_n266), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n200), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  INV_X1    g104(.A(new_n278), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n279), .A2(new_n286), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n279), .A2(new_n286), .A3(new_n292), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n187), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n298), .ZN(new_n300));
  AOI211_X1 g114(.A(KEYINPUT32), .B(new_n300), .C1(new_n294), .C2(new_n296), .ZN(new_n301));
  INV_X1    g115(.A(new_n285), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n277), .A2(KEYINPUT29), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT71), .B1(new_n255), .B2(new_n200), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n283), .A2(new_n270), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(KEYINPUT71), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n302), .B(new_n303), .C1(new_n306), .C2(new_n280), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n277), .B1(new_n284), .B2(new_n285), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n289), .A2(new_n270), .A3(new_n276), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G472), .ZN(new_n316));
  OAI22_X1  g130(.A1(new_n299), .A2(new_n301), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(new_n208), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  AND4_X1   g138(.A1(new_n318), .A2(new_n322), .A3(new_n324), .A4(new_n208), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n322), .A2(KEYINPUT16), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(G146), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n245), .A2(G119), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n245), .A2(KEYINPUT23), .A3(G119), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n192), .A2(G128), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT74), .B(G110), .Z(new_n337));
  OR2_X1    g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n331), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT24), .B(G110), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n338), .A2(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n330), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n336), .A2(KEYINPUT73), .ZN(new_n346));
  OAI21_X1  g160(.A(G110), .B1(new_n336), .B2(KEYINPUT73), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n327), .A2(new_n328), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n208), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n329), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n341), .A2(new_n342), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT22), .B(G137), .ZN(new_n354));
  INV_X1    g168(.A(G221), .ZN(new_n355));
  INV_X1    g169(.A(G234), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n355), .A2(new_n356), .A3(G953), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n354), .B(new_n357), .Z(new_n358));
  NAND3_X1  g172(.A1(new_n345), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n358), .ZN(new_n360));
  INV_X1    g174(.A(new_n353), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(new_n344), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n362), .A3(new_n309), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n359), .A2(new_n362), .A3(KEYINPUT25), .A4(new_n309), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(G234), .B2(new_n309), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n359), .A2(new_n362), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(G902), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n367), .A2(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G469), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(new_n374), .B2(G107), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n376));
  INV_X1    g190(.A(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(G104), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT77), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n375), .A2(new_n378), .A3(KEYINPUT77), .A4(new_n379), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n265), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(G101), .A3(new_n383), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n375), .A2(new_n378), .A3(new_n384), .A4(new_n379), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(KEYINPUT4), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n374), .A2(G107), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n377), .A2(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT10), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n388), .A2(new_n392), .B1(new_n259), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT78), .B1(new_n246), .B2(new_n202), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n205), .A2(G146), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n237), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n243), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n235), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n396), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n400), .B1(new_n408), .B2(new_n397), .ZN(new_n409));
  AOI211_X1 g223(.A(KEYINPUT79), .B(KEYINPUT10), .C1(new_n406), .C2(new_n407), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n399), .B(new_n233), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G140), .ZN(new_n412));
  INV_X1    g226(.A(G953), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G227), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n412), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n235), .B(new_n396), .C1(new_n257), .C2(new_n258), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n408), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT12), .A3(new_n264), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT12), .B1(new_n418), .B2(new_n264), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n409), .A2(new_n410), .ZN(new_n424));
  INV_X1    g238(.A(new_n392), .ZN(new_n425));
  INV_X1    g239(.A(new_n398), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n425), .A2(new_n387), .B1(new_n248), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n264), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n415), .B1(new_n428), .B2(new_n411), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n373), .B(new_n309), .C1(new_n423), .C2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n373), .A2(new_n309), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n411), .A3(new_n415), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n424), .A2(new_n427), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n418), .A2(new_n264), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT12), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n434), .A2(new_n233), .B1(new_n419), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(G469), .B(new_n433), .C1(new_n438), .C2(new_n415), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n432), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT9), .B(G234), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n355), .B1(new_n442), .B2(new_n309), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n272), .A2(G143), .A3(G214), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(G143), .B1(new_n272), .B2(G214), .ZN(new_n448));
  OAI21_X1  g262(.A(G131), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  INV_X1    g264(.A(G237), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n413), .A3(G214), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n205), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n229), .A3(new_n446), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT17), .B(G131), .C1(new_n447), .C2(new_n448), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n350), .A3(new_n329), .A4(new_n456), .ZN(new_n457));
  OAI22_X1  g271(.A1(new_n320), .A2(new_n325), .B1(new_n208), .B2(new_n319), .ZN(new_n458));
  NAND2_X1  g272(.A1(KEYINPUT18), .A2(G131), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n446), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n453), .B2(new_n446), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n463));
  AOI211_X1 g277(.A(new_n463), .B(new_n459), .C1(new_n453), .C2(new_n446), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n458), .B(new_n460), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(G113), .B(G122), .Z(new_n466));
  XOR2_X1   g280(.A(KEYINPUT90), .B(G104), .Z(new_n467));
  XOR2_X1   g281(.A(new_n466), .B(new_n467), .Z(new_n468));
  NAND3_X1  g282(.A1(new_n457), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT91), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n457), .A2(new_n465), .A3(new_n471), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n457), .A2(new_n465), .ZN(new_n474));
  INV_X1    g288(.A(new_n468), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT93), .B(G475), .Z(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n449), .A2(new_n454), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT88), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n319), .A2(KEYINPUT89), .A3(KEYINPUT19), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT19), .B1(new_n319), .B2(KEYINPUT89), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n208), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n329), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n481), .A2(KEYINPUT88), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n465), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n475), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n480), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n470), .A2(new_n472), .B1(new_n488), .B2(new_n475), .ZN(new_n491));
  NOR2_X1   g305(.A1(G475), .A2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n490), .A2(KEYINPUT20), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n491), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(new_n480), .A3(new_n496), .A4(new_n492), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n479), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n205), .A2(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n245), .A2(G143), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(G134), .ZN(new_n502));
  INV_X1    g316(.A(G122), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G116), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n194), .A2(G122), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n504), .B2(new_n505), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n377), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n194), .A2(KEYINPUT14), .A3(G122), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n505), .ZN(new_n511));
  OAI211_X1 g325(.A(G107), .B(new_n510), .C1(new_n511), .C2(KEYINPUT14), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n502), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT95), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n205), .A2(G128), .ZN(new_n515));
  OAI21_X1  g329(.A(G134), .B1(new_n515), .B2(KEYINPUT13), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n501), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT13), .A4(G134), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n511), .A2(KEYINPUT94), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(G107), .A3(new_n520), .ZN(new_n521));
  AOI221_X4 g335(.A(new_n514), .B1(new_n517), .B2(new_n518), .C1(new_n509), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n509), .A2(new_n521), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n518), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT95), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n513), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n441), .A2(new_n368), .A3(G953), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT96), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n513), .B(new_n527), .C1(new_n522), .C2(new_n525), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(KEYINPUT96), .A3(new_n528), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n309), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n536), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n532), .A2(new_n309), .A3(new_n533), .A4(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(G902), .B(G953), .C1(new_n356), .C2(new_n451), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n541), .B(KEYINPUT97), .Z(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT21), .B(G898), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n413), .A2(G952), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n356), .B2(new_n451), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n498), .A2(new_n540), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT86), .Z(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G224), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(G953), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n215), .A2(G125), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT83), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT83), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n215), .A2(new_n557), .A3(G125), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(G125), .B(new_n236), .C1(new_n244), .C2(new_n247), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT7), .B(new_n554), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n560), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n554), .A2(KEYINPUT7), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n555), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g379(.A(G110), .B(G122), .Z(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT81), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT5), .ZN(new_n570));
  OR3_X1    g384(.A1(new_n194), .A2(KEYINPUT5), .A3(G119), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(G113), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n199), .A2(new_n407), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT80), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n198), .A2(new_n190), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT80), .A4(G113), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n407), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT85), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n572), .A2(new_n574), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n199), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n396), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT85), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n569), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n200), .A2(new_n392), .A3(new_n386), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n407), .A3(new_n576), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n567), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n565), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n309), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n562), .A2(new_n553), .A3(new_n556), .A4(new_n558), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n585), .A2(new_n586), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n567), .B(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n585), .A2(new_n586), .A3(new_n567), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT6), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n593), .A2(KEYINPUT6), .A3(new_n594), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n592), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n551), .B1(new_n589), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G214), .B1(G237), .B2(G902), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n587), .A2(KEYINPUT6), .B1(new_n593), .B2(new_n594), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n593), .A2(KEYINPUT6), .A3(new_n594), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n591), .B(new_n590), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(new_n309), .A3(new_n550), .A4(new_n588), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n445), .A2(new_n548), .A3(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n317), .A2(new_n372), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n384), .ZN(G3));
  NAND2_X1  g424(.A1(new_n297), .A2(new_n309), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n297), .A2(new_n298), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n440), .A2(new_n372), .A3(new_n444), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n494), .A2(new_n497), .ZN(new_n618));
  INV_X1    g432(.A(new_n479), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n535), .A2(G902), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n623));
  INV_X1    g437(.A(new_n513), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n507), .A2(new_n508), .A3(new_n377), .ZN(new_n625));
  AOI21_X1  g439(.A(G107), .B1(new_n519), .B2(new_n520), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n524), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n514), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n523), .A2(KEYINPUT95), .A3(new_n524), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n623), .B1(new_n630), .B2(new_n527), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n531), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n623), .A3(new_n527), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(KEYINPUT33), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n532), .A2(new_n636), .A3(new_n533), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n631), .B2(new_n531), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(KEYINPUT99), .A3(new_n633), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n622), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n534), .A2(new_n535), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n620), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n601), .A2(new_n606), .A3(new_n602), .A4(new_n547), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n617), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT98), .B1(new_n526), .B2(new_n528), .ZN(new_n647));
  INV_X1    g461(.A(new_n531), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT33), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n633), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n649), .A2(new_n635), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT99), .B1(new_n639), .B2(new_n633), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n637), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n642), .B1(new_n653), .B2(new_n622), .ZN(new_n654));
  INV_X1    g468(.A(new_n645), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n654), .A2(KEYINPUT100), .A3(new_n655), .A4(new_n620), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n646), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n616), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  OAI21_X1  g474(.A(KEYINPUT20), .B1(new_n491), .B2(new_n493), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n495), .A2(new_n496), .A3(new_n492), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n479), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n537), .A2(new_n539), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n547), .B(KEYINPUT101), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n607), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n663), .A2(KEYINPUT102), .A3(new_n664), .A4(new_n665), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n616), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  AND3_X1   g488(.A1(new_n498), .A2(new_n540), .A3(new_n547), .ZN(new_n675));
  AOI21_X1  g489(.A(G902), .B1(new_n294), .B2(new_n296), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n675), .B(new_n613), .C1(new_n316), .C2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n440), .A2(new_n444), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n345), .A2(new_n353), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n367), .A2(new_n369), .B1(new_n371), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n678), .A2(new_n669), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT37), .B(G110), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G12));
  NOR3_X1   g501(.A1(new_n445), .A2(new_n607), .A3(new_n682), .ZN(new_n688));
  INV_X1    g502(.A(new_n546), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n689), .B1(new_n542), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n663), .A2(new_n664), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n317), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  NAND2_X1  g509(.A1(new_n601), .A2(new_n606), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  INV_X1    g511(.A(new_n602), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n620), .A2(new_n664), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n697), .A2(new_n698), .A3(new_n683), .A4(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n691), .B(KEYINPUT39), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n678), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n306), .A2(new_n276), .ZN(new_n704));
  INV_X1    g518(.A(new_n270), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n277), .B1(new_n269), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n708));
  AOI21_X1  g522(.A(G902), .B1(new_n707), .B2(KEYINPUT103), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI22_X1  g524(.A1(new_n299), .A2(new_n301), .B1(new_n710), .B2(new_n316), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n700), .A2(new_n703), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  OAI211_X1 g528(.A(new_n620), .B(new_n692), .C1(new_n641), .C2(new_n643), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n317), .A2(new_n688), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  OAI21_X1  g532(.A(new_n309), .B1(new_n423), .B2(new_n429), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n444), .A3(new_n430), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n720), .A2(KEYINPUT104), .A3(new_n444), .A4(new_n430), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n723), .A2(new_n372), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n657), .A2(new_n317), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n671), .A3(new_n317), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT105), .B(G116), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G18));
  AND3_X1   g545(.A1(new_n723), .A2(new_n669), .A3(new_n724), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n317), .A3(new_n675), .A4(new_n683), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  INV_X1    g548(.A(new_n665), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n498), .A2(new_n540), .A3(new_n735), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n669), .A2(new_n723), .A3(new_n724), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n292), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT71), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n283), .B2(new_n270), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT28), .B1(new_n741), .B2(new_n304), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n302), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n739), .B1(new_n743), .B2(new_n276), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n738), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n277), .B1(new_n742), .B2(new_n302), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT106), .B1(new_n747), .B2(new_n739), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n300), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n372), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT107), .B(G472), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n297), .B2(new_n309), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n749), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n737), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT108), .B(G122), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G24));
  AND4_X1   g571(.A1(new_n669), .A2(new_n723), .A3(new_n683), .A4(new_n724), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n749), .A2(new_n715), .A3(new_n753), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  AOI21_X1  g575(.A(KEYINPUT109), .B1(new_n696), .B2(new_n602), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n763), .B(new_n698), .C1(new_n601), .C2(new_n606), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n762), .A2(new_n764), .A3(new_n445), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n317), .A2(new_n765), .A3(new_n372), .A4(new_n716), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n715), .A2(new_n762), .A3(new_n764), .A4(new_n445), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(KEYINPUT42), .A3(new_n317), .A4(new_n372), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NAND4_X1  g586(.A1(new_n317), .A2(new_n765), .A3(new_n372), .A4(new_n693), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  OAI21_X1  g588(.A(new_n433), .B1(new_n438), .B2(new_n415), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n373), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n432), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n430), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n444), .B(new_n701), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n654), .A2(new_n498), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT43), .Z(new_n789));
  AOI21_X1  g603(.A(new_n682), .B1(new_n612), .B2(new_n613), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT44), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(KEYINPUT44), .A3(new_n790), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n762), .A2(new_n764), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n787), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n219), .ZN(G39));
  OAI21_X1  g610(.A(new_n444), .B1(new_n785), .B2(new_n786), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT47), .B(new_n444), .C1(new_n785), .C2(new_n786), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n793), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n317), .A2(new_n802), .A3(new_n372), .A4(new_n715), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NAND2_X1  g619(.A1(new_n723), .A2(new_n724), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n793), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT113), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n546), .B1(new_n808), .B2(KEYINPUT113), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n711), .A2(new_n750), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n620), .A3(new_n654), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n789), .A2(new_n689), .A3(new_n754), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(new_n732), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n545), .B(new_n814), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n809), .A2(new_n789), .A3(new_n810), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT114), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n744), .A2(new_n745), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n748), .A3(new_n292), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n824), .A2(new_n298), .B1(new_n611), .B2(new_n751), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n683), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n807), .A2(new_n698), .A3(new_n697), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n815), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n815), .A2(KEYINPUT50), .A3(new_n827), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n654), .A2(new_n620), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n830), .A2(new_n831), .B1(new_n813), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n720), .A2(new_n430), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n443), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n799), .A2(new_n800), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n815), .A2(new_n793), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n820), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n317), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n750), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n822), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT48), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n826), .A2(new_n833), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n801), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n799), .A2(KEYINPUT112), .A3(new_n800), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n837), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n846), .B1(new_n850), .B2(new_n839), .ZN(new_n851));
  XNOR2_X1  g665(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n841), .B(new_n845), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n664), .A2(new_n691), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n683), .A2(new_n663), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n317), .A2(new_n765), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n765), .A2(new_n825), .A3(new_n683), .A4(new_n716), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n773), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n771), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n620), .B(new_n642), .C1(new_n653), .C2(new_n622), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n498), .A2(new_n540), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n669), .A3(new_n861), .A4(new_n665), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n615), .A2(new_n862), .B1(new_n677), .B2(new_n684), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n609), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n613), .A2(KEYINPUT32), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n297), .A2(new_n187), .A3(new_n298), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(G472), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n548), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n870), .A2(new_n758), .B1(new_n754), .B2(new_n737), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n317), .B(new_n725), .C1(new_n657), .C2(new_n671), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n859), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n620), .A2(new_n682), .A3(new_n664), .A4(new_n692), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n875), .A2(new_n445), .A3(new_n607), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n711), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n760), .A2(new_n694), .A3(new_n717), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n874), .A2(new_n880), .A3(KEYINPUT53), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n726), .A2(new_n733), .A3(new_n755), .A4(new_n729), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n771), .A3(new_n864), .A4(new_n858), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n684), .B1(new_n867), .B2(new_n869), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n885), .A2(new_n693), .B1(new_n758), .B2(new_n759), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n717), .A2(new_n877), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n879), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n723), .A2(new_n669), .A3(new_n683), .A4(new_n724), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n825), .A2(new_n716), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n694), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n717), .A2(new_n877), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT52), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n882), .B1(new_n884), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n881), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n853), .A2(new_n901), .B1(G952), .B2(G953), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n836), .B(KEYINPUT49), .Z(new_n903));
  NAND3_X1  g717(.A1(new_n697), .A2(new_n602), .A3(new_n444), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n903), .A2(new_n788), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n902), .B1(new_n812), .B2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n413), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n897), .A2(new_n309), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n909), .B2(new_n550), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n598), .A2(new_n599), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT116), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n592), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n908), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n910), .B2(new_n915), .ZN(G51));
  XNOR2_X1  g731(.A(new_n431), .B(KEYINPUT57), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n901), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n429), .B2(new_n423), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n909), .A2(new_n779), .A3(new_n780), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n907), .B1(new_n920), .B2(new_n921), .ZN(G54));
  NAND2_X1  g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT117), .Z(new_n924));
  AND3_X1   g738(.A1(new_n909), .A2(new_n495), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n495), .B1(new_n909), .B2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n907), .ZN(G60));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT59), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n898), .A2(new_n900), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(new_n653), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT118), .B1(new_n931), .B2(new_n908), .ZN(new_n932));
  OAI211_X1 g746(.A(KEYINPUT118), .B(new_n908), .C1(new_n930), .C2(new_n653), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n653), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n932), .A2(new_n935), .ZN(G63));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n368), .A2(new_n309), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT53), .B1(new_n874), .B2(new_n880), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n884), .A2(new_n894), .A3(new_n882), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n681), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  INV_X1    g758(.A(new_n940), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n881), .B2(new_n895), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n908), .B1(new_n946), .B2(new_n370), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n937), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n949));
  INV_X1    g763(.A(new_n370), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n907), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n946), .B2(new_n681), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(KEYINPUT121), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n946), .A2(KEYINPUT120), .A3(new_n681), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n943), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n951), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n952), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT122), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n955), .A2(new_n960), .A3(KEYINPUT122), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G66));
  OAI21_X1  g779(.A(G953), .B1(new_n543), .B2(new_n552), .ZN(new_n966));
  INV_X1    g780(.A(new_n873), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(G953), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n912), .B1(G898), .B2(new_n413), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G69));
  AOI21_X1  g784(.A(new_n795), .B1(new_n801), .B2(new_n803), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n891), .B1(new_n885), .B2(new_n716), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n771), .A3(new_n773), .ZN(new_n973));
  INV_X1    g787(.A(new_n787), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n842), .A2(new_n750), .A3(new_n607), .A4(new_n699), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n413), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n287), .A2(new_n288), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n483), .A2(new_n484), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(G900), .B2(G953), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n972), .A2(new_n713), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n802), .A2(new_n702), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n988), .A2(new_n861), .A3(new_n860), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n987), .B1(new_n843), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n971), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n413), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n981), .B(KEYINPUT123), .ZN(new_n993));
  AOI22_X1  g807(.A1(new_n978), .A2(new_n982), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n413), .B1(G227), .B2(G900), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n994), .B(new_n996), .ZN(G72));
  XOR2_X1   g811(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n998));
  NOR2_X1   g812(.A1(new_n316), .A2(new_n309), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n706), .A2(new_n313), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT127), .B1(new_n896), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n896), .A2(KEYINPUT127), .A3(new_n1003), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1000), .B1(new_n977), .B2(new_n967), .ZN(new_n1006));
  OAI221_X1 g820(.A(new_n908), .B1(new_n1004), .B2(new_n1005), .C1(new_n1006), .C2(new_n313), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n986), .A2(new_n971), .A3(new_n967), .A4(new_n990), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n706), .B1(new_n1008), .B2(new_n1001), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .ZN(G57));
endmodule


