//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1221,
    new_n1222, new_n1223;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT2), .B(G226), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G97), .B(G107), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  AND2_X1   g0040(.A1(KEYINPUT3), .A2(G33), .ZN(new_n241));
  NOR2_X1   g0041(.A1(KEYINPUT3), .A2(G33), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G1698), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g0045(.A1(new_n245), .A2(G223), .B1(G77), .B2(new_n243), .ZN(new_n246));
  INV_X1    g0046(.A(G222), .ZN(new_n247));
  OR2_X1    g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n244), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n246), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n205), .B(G274), .C1(G41), .C2(G45), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT64), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n253), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(G226), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT65), .A2(G179), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT65), .A2(G179), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g0068(.A(new_n268), .B(KEYINPUT66), .Z(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n214), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(new_n205), .B2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n274), .A2(new_n206), .A3(G1), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  XOR2_X1   g0083(.A(KEYINPUT8), .B(G58), .Z(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n271), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n273), .B1(G50), .B2(new_n276), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(new_n264), .B2(G169), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n269), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n264), .A2(G190), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT69), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n287), .A2(KEYINPUT9), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(KEYINPUT9), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(new_n293), .B1(G200), .B2(new_n263), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n264), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(KEYINPUT10), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n291), .A2(new_n300), .A3(new_n294), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n289), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT16), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n249), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT73), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n243), .A2(KEYINPUT73), .A3(KEYINPUT7), .A4(new_n206), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n248), .A2(new_n206), .A3(new_n249), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n304), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G58), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n304), .ZN(new_n315));
  OAI21_X1  g0115(.A(G20), .B1(new_n315), .B2(new_n201), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n279), .A2(G159), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n303), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n312), .A2(new_n305), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n320), .B2(G68), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n286), .B1(new_n321), .B2(KEYINPUT16), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n284), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n205), .B2(G20), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n275), .A2(new_n271), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n325), .A2(new_n326), .B1(new_n275), .B2(new_n324), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n256), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(G223), .A2(G1698), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n330), .B1(G226), .B2(new_n244), .C1(new_n241), .C2(new_n242), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n258), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n256), .A2(new_n328), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n297), .B1(new_n337), .B2(new_n333), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT17), .ZN(new_n341));
  AND4_X1   g0141(.A1(new_n323), .A2(new_n327), .A3(new_n339), .A4(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n343));
  INV_X1    g0143(.A(new_n327), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n319), .B2(new_n322), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n329), .B2(new_n334), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n337), .A2(new_n333), .A3(new_n267), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n243), .B2(new_n206), .ZN(new_n353));
  NOR4_X1   g0153(.A1(new_n241), .A2(new_n242), .A3(new_n311), .A4(G20), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n318), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(KEYINPUT16), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n271), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n353), .B1(new_n307), .B2(new_n308), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n356), .B1(new_n359), .B2(new_n304), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n303), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n348), .B(new_n352), .C1(new_n361), .C2(new_n344), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n350), .A2(new_n351), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT18), .B1(new_n345), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n347), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G77), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n275), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n272), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n367), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT67), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n283), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n284), .A2(new_n279), .B1(G20), .B2(G77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n370), .B1(new_n376), .B2(new_n271), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT68), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n377), .B(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n245), .A2(G238), .B1(G107), .B2(new_n243), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n250), .A2(G232), .A3(new_n244), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n253), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n257), .B1(G244), .B2(new_n261), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G200), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n335), .B2(new_n385), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n267), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n349), .B2(new_n385), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n379), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n302), .A2(new_n366), .A3(new_n388), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n250), .A2(G226), .A3(new_n244), .ZN(new_n394));
  OAI211_X1 g0194(.A(G232), .B(G1698), .C1(new_n241), .C2(new_n242), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT71), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n394), .A2(KEYINPUT71), .A3(new_n395), .A4(new_n396), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n253), .ZN(new_n401));
  INV_X1    g0201(.A(G238), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n256), .B1(new_n260), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n258), .B1(new_n397), .B2(new_n398), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n407), .B2(new_n400), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT13), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(G179), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n406), .A2(KEYINPUT72), .A3(new_n410), .ZN(new_n413));
  OR3_X1    g0213(.A1(new_n408), .A2(KEYINPUT72), .A3(new_n409), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(G169), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n413), .A2(KEYINPUT14), .A3(new_n414), .A4(G169), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n412), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n283), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n420), .A2(new_n367), .B1(new_n206), .B2(G68), .ZN(new_n421));
  INV_X1    g0221(.A(G50), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n280), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n271), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n276), .A2(KEYINPUT12), .A3(G68), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT12), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n275), .B2(new_n304), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n428), .A2(new_n430), .B1(new_n369), .B2(new_n304), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n426), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n419), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n413), .A2(G200), .A3(new_n414), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n335), .B1(new_n408), .B2(new_n409), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n406), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n393), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT78), .B(G116), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n206), .A3(G33), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT83), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n206), .A2(G107), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT23), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT83), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n441), .A2(new_n446), .A3(new_n206), .A4(G33), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n250), .A2(new_n206), .A3(G87), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT22), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT24), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n450), .B(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT24), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n271), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n205), .A2(G33), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n276), .A2(new_n286), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G107), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT25), .B1(new_n275), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n275), .A2(KEYINPUT25), .A3(new_n462), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n461), .A2(G107), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n458), .A2(new_n459), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n286), .B1(new_n453), .B2(new_n456), .ZN(new_n468));
  INV_X1    g0268(.A(new_n466), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT84), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n243), .A2(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G250), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n245), .A2(G257), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT85), .B(G294), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G33), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n205), .A2(G45), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n253), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n476), .A2(new_n253), .B1(G264), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n479), .A2(G274), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n258), .A3(new_n477), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G169), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(G179), .A3(new_n483), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n467), .A2(new_n470), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(G200), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(G190), .A3(new_n483), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n458), .A2(new_n489), .A3(new_n466), .A4(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n250), .A2(G244), .A3(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n441), .A2(G33), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n494), .C1(new_n251), .C2(new_n402), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n253), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n478), .A2(G250), .ZN(new_n497));
  OR3_X1    g0297(.A1(new_n253), .A2(new_n497), .A3(KEYINPUT77), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT77), .B1(new_n253), .B2(new_n497), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n482), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT79), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT79), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(G190), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT81), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(new_n504), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n502), .A2(KEYINPUT81), .A3(G190), .A4(new_n504), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT19), .ZN(new_n511));
  INV_X1    g0311(.A(G97), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n420), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n250), .A2(new_n206), .A3(G68), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n206), .B1(new_n396), .B2(new_n511), .ZN(new_n515));
  INV_X1    g0315(.A(G87), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n512), .A3(new_n462), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n371), .B(KEYINPUT67), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n519), .A2(new_n271), .B1(new_n520), .B2(new_n275), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n461), .A2(G87), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n507), .A2(new_n509), .A3(new_n510), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n508), .A2(new_n349), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n502), .A2(new_n267), .A3(new_n504), .ZN(new_n526));
  INV_X1    g0326(.A(new_n461), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n521), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT80), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n528), .A2(KEYINPUT80), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n525), .A2(new_n526), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(new_n206), .C1(G33), .C2(new_n512), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n271), .B(new_n534), .C1(new_n441), .C2(new_n206), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT20), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n441), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n461), .A2(G116), .B1(new_n275), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n471), .A2(G257), .B1(G303), .B2(new_n243), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n245), .A2(G264), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n253), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n480), .A2(G270), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(KEYINPUT82), .A3(new_n483), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT82), .B1(new_n545), .B2(new_n483), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n540), .B1(new_n549), .B2(G200), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n335), .B2(new_n549), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT21), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n545), .A2(new_n483), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT82), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n546), .B1(new_n253), .B2(new_n543), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n540), .A2(G169), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n549), .A2(KEYINPUT21), .A3(G169), .A4(new_n540), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(G179), .A3(new_n540), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n551), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n480), .A2(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n483), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  INV_X1    g0364(.A(G244), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n251), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n245), .A2(G250), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n244), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n533), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n563), .B1(new_n569), .B2(new_n253), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n349), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n267), .ZN(new_n573));
  XNOR2_X1  g0373(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n512), .A2(G107), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n237), .A2(new_n574), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(G20), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n279), .A2(G77), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(KEYINPUT76), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT76), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n359), .A2(new_n462), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n286), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n276), .A2(G97), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n461), .B2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n572), .B(new_n573), .C1(new_n585), .C2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n582), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(new_n584), .A3(new_n580), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n271), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n571), .A2(G200), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n570), .A2(G190), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n587), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n561), .A2(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n440), .A2(new_n492), .A3(new_n532), .A4(new_n597), .ZN(G372));
  OAI21_X1  g0398(.A(new_n573), .B1(G169), .B2(new_n570), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n592), .B2(new_n587), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n524), .A2(new_n600), .A3(new_n531), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT26), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n458), .A2(new_n466), .B1(new_n485), .B2(new_n486), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n589), .B(new_n595), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n501), .A2(G200), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n507), .A2(new_n510), .A3(new_n523), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n501), .A2(new_n349), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n530), .A2(new_n526), .A3(new_n529), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n491), .A3(new_n609), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n601), .A2(new_n602), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n600), .A3(new_n609), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n609), .B1(new_n612), .B2(KEYINPUT26), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n440), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n365), .ZN(new_n616));
  INV_X1    g0416(.A(new_n392), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n433), .B1(new_n438), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n618), .B2(new_n347), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n299), .A2(new_n301), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n289), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n615), .A2(new_n621), .ZN(G369));
  NAND3_X1  g0422(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n537), .B2(new_n539), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n604), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n561), .B2(new_n630), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT86), .ZN(new_n633));
  INV_X1    g0433(.A(G330), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n467), .A2(new_n470), .A3(new_n628), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n492), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n488), .A2(new_n629), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n603), .A2(new_n629), .ZN(new_n642));
  INV_X1    g0442(.A(new_n604), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n628), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n492), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n642), .A3(new_n645), .ZN(G399));
  OR2_X1    g0446(.A1(new_n517), .A2(G116), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT87), .ZN(new_n648));
  INV_X1    g0448(.A(new_n209), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G41), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n648), .A2(new_n650), .A3(new_n205), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n213), .B2(new_n650), .ZN(new_n652));
  XOR2_X1   g0452(.A(new_n652), .B(KEYINPUT28), .Z(new_n653));
  INV_X1    g0453(.A(KEYINPUT30), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n502), .A2(new_n481), .A3(new_n504), .A4(new_n570), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n544), .B(G179), .C1(new_n547), .C2(new_n548), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n504), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n503), .B1(new_n496), .B2(new_n500), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n656), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n570), .A2(new_n481), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(KEYINPUT30), .A4(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n389), .B1(new_n496), .B2(new_n500), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n571), .A2(new_n549), .A3(new_n484), .A4(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n657), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n666), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT31), .B1(new_n666), .B2(new_n628), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n597), .A2(new_n492), .A3(new_n532), .A4(new_n629), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n614), .A2(new_n629), .ZN(new_n674));
  XNOR2_X1  g0474(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n601), .A2(new_n602), .ZN(new_n677));
  INV_X1    g0477(.A(new_n609), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n612), .B2(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n596), .A2(KEYINPUT89), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT89), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n589), .A2(new_n595), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n488), .A2(new_n643), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n677), .B(new_n679), .C1(new_n684), .C2(new_n610), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(KEYINPUT29), .A3(new_n629), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n673), .B1(new_n676), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n653), .B1(new_n687), .B2(G1), .ZN(G364));
  INV_X1    g0488(.A(new_n635), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n633), .A2(new_n634), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n274), .A2(G20), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n205), .B1(new_n691), .B2(G45), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n650), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n689), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(G13), .A2(G33), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G20), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n633), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n214), .B1(G20), .B2(new_n349), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n209), .A2(new_n250), .ZN(new_n704));
  XNOR2_X1  g0504(.A(G355), .B(KEYINPUT90), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n704), .A2(new_n705), .B1(G116), .B2(new_n209), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n649), .A2(new_n250), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G45), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n213), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n236), .A2(new_n709), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n706), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n206), .A2(new_n335), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n297), .A2(G179), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n243), .B1(new_n716), .B2(G87), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n206), .A2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n714), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n389), .A2(G200), .A3(new_n718), .ZN(new_n720));
  OAI221_X1 g0520(.A(new_n717), .B1(new_n462), .B2(new_n719), .C1(new_n720), .C2(new_n304), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n335), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n206), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G97), .ZN(new_n725));
  INV_X1    g0525(.A(new_n713), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n297), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n389), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n726), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n389), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n725), .B1(new_n728), .B2(new_n422), .C1(new_n314), .C2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n389), .A2(new_n297), .A3(new_n718), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n721), .B(new_n731), .C1(G77), .C2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n718), .A2(new_n735), .A3(new_n297), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT91), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G159), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT32), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n243), .B1(new_n719), .B2(new_n744), .C1(new_n745), .C2(new_n715), .ZN(new_n746));
  INV_X1    g0546(.A(G329), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT33), .B(G317), .Z(new_n748));
  OAI22_X1  g0548(.A1(new_n740), .A2(new_n747), .B1(new_n720), .B2(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n746), .B(new_n749), .C1(G311), .C2(new_n733), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT92), .B(G326), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n728), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n730), .A2(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n752), .B(new_n754), .C1(new_n474), .C2(new_n724), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n734), .A2(new_n743), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n701), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n694), .B1(new_n703), .B2(new_n712), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT93), .Z(new_n759));
  NAND2_X1  g0559(.A1(new_n700), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n696), .A2(new_n760), .ZN(G396));
  NOR2_X1   g0561(.A1(new_n701), .A2(new_n697), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n695), .B1(new_n367), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n725), .B1(new_n728), .B2(new_n745), .C1(new_n764), .C2(new_n730), .ZN(new_n765));
  INV_X1    g0565(.A(G311), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n740), .A2(new_n766), .B1(new_n538), .B2(new_n732), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n720), .A2(new_n744), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n243), .B1(new_n719), .B2(new_n516), .C1(new_n462), .C2(new_n715), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n765), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n728), .ZN(new_n771));
  INV_X1    g0571(.A(new_n730), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G137), .A2(new_n771), .B1(new_n772), .B2(G143), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n773), .B1(new_n278), .B2(new_n720), .C1(new_n741), .C2(new_n732), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT34), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n243), .B1(new_n716), .B2(G50), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n776), .B1(new_n314), .B2(new_n723), .C1(new_n304), .C2(new_n719), .ZN(new_n777));
  INV_X1    g0577(.A(new_n740), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n777), .B1(G132), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n770), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n392), .A2(new_n628), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n379), .A2(new_n628), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n388), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n783), .B2(new_n392), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n763), .B1(new_n757), .B2(new_n780), .C1(new_n784), .C2(new_n698), .ZN(new_n785));
  INV_X1    g0585(.A(new_n784), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n674), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n629), .B(new_n784), .C1(new_n611), .C2(new_n613), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(KEYINPUT94), .A3(new_n672), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n790), .B(new_n695), .C1(new_n672), .C2(new_n789), .ZN(new_n791));
  AOI21_X1  g0591(.A(KEYINPUT94), .B1(new_n789), .B2(new_n672), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n785), .B1(new_n791), .B2(new_n792), .ZN(G384));
  INV_X1    g0593(.A(KEYINPUT100), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n347), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n342), .A2(new_n346), .A3(KEYINPUT100), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n795), .A2(new_n365), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n323), .A2(new_n327), .ZN(new_n798));
  INV_X1    g0598(.A(new_n626), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n352), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT37), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n345), .A2(new_n339), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n801), .A2(new_n800), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT99), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n801), .A2(new_n800), .A3(new_n803), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n804), .A2(KEYINPUT99), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n797), .A2(new_n800), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n355), .A2(new_n356), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n303), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n322), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n626), .B1(new_n814), .B2(new_n327), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n347), .B2(new_n365), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n345), .A2(new_n339), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n363), .A2(new_n626), .B1(new_n814), .B2(new_n327), .ZN(new_n818));
  OAI21_X1  g0618(.A(KEYINPUT37), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n816), .A2(KEYINPUT38), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n811), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n432), .A2(new_n629), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n438), .B(new_n824), .C1(new_n419), .C2(new_n432), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n417), .A2(new_n418), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n823), .B1(new_n826), .B2(new_n412), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n828), .A2(new_n671), .A3(new_n784), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n822), .A2(new_n829), .A3(KEYINPUT40), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT101), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n828), .A2(new_n671), .A3(new_n784), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT97), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n821), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n816), .A2(new_n820), .A3(KEYINPUT97), .A4(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n816), .A2(new_n820), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n810), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT98), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT38), .B1(new_n816), .B2(new_n820), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n834), .B2(new_n821), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n843), .A2(KEYINPUT98), .A3(new_n836), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n833), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n832), .B1(new_n845), .B2(KEYINPUT40), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT98), .B1(new_n843), .B2(new_n836), .ZN(new_n847));
  AND4_X1   g0647(.A1(KEYINPUT98), .A2(new_n835), .A3(new_n836), .A4(new_n838), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n829), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT40), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(KEYINPUT101), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n831), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n440), .A2(new_n671), .ZN(new_n854));
  OAI21_X1  g0654(.A(G330), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n811), .A2(new_n857), .A3(new_n821), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n434), .A2(new_n628), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n781), .B(KEYINPUT96), .Z(new_n863));
  NAND2_X1  g0663(.A1(new_n788), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n828), .B(new_n864), .C1(new_n847), .C2(new_n848), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n365), .A2(new_n626), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n440), .A2(new_n676), .A3(new_n686), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n621), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n867), .B(new_n869), .Z(new_n870));
  OR2_X1    g0670(.A1(new_n856), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n856), .A2(new_n870), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n871), .B(new_n872), .C1(new_n205), .C2(new_n691), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n576), .A2(KEYINPUT35), .A3(new_n577), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(G116), .A3(new_n215), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT35), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n576), .A2(new_n577), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n878), .A2(KEYINPUT36), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(KEYINPUT36), .ZN(new_n880));
  OAI21_X1  g0680(.A(G77), .B1(new_n314), .B2(new_n304), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n212), .A2(new_n881), .B1(G50), .B2(new_n304), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(G1), .A3(new_n274), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT95), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n873), .A2(new_n879), .A3(new_n880), .A4(new_n884), .ZN(G367));
  OAI221_X1 g0685(.A(new_n702), .B1(new_n209), .B2(new_n520), .C1(new_n708), .C2(new_n232), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n716), .A2(KEYINPUT46), .A3(G116), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n243), .C1(new_n512), .C2(new_n719), .ZN(new_n888));
  INV_X1    g0688(.A(new_n720), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n474), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n778), .A2(G317), .B1(G283), .B2(new_n733), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n772), .A2(G303), .B1(G107), .B2(new_n724), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT46), .B1(new_n716), .B2(new_n441), .ZN(new_n893));
  XOR2_X1   g0693(.A(KEYINPUT105), .B(G311), .Z(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n771), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n243), .B1(new_n716), .B2(G58), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n367), .B2(new_n719), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(G50), .B2(new_n733), .ZN(new_n899));
  INV_X1    g0699(.A(G137), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n899), .B1(new_n900), .B2(new_n740), .C1(new_n741), .C2(new_n720), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n724), .A2(G68), .ZN(new_n902));
  INV_X1    g0702(.A(G143), .ZN(new_n903));
  OAI221_X1 g0703(.A(new_n902), .B1(new_n728), .B2(new_n903), .C1(new_n278), .C2(new_n730), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n896), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT47), .Z(new_n906));
  OAI211_X1 g0706(.A(new_n694), .B(new_n886), .C1(new_n906), .C2(new_n757), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n523), .A2(new_n629), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n607), .B2(new_n609), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n609), .B2(new_n908), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT102), .Z(new_n911));
  AOI21_X1  g0711(.A(new_n907), .B1(new_n911), .B2(new_n699), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT104), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n628), .B1(new_n585), .B2(new_n588), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n680), .A2(new_n682), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n600), .B2(new_n628), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n645), .A2(new_n642), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT44), .Z(new_n920));
  NOR2_X1   g0720(.A1(new_n917), .A2(new_n918), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT45), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(new_n641), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n645), .B1(new_n640), .B2(new_n644), .C1(new_n635), .C2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n689), .A2(KEYINPUT103), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n687), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n687), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n650), .B(KEYINPUT41), .Z(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n913), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(KEYINPUT104), .B(new_n933), .C1(new_n931), .C2(new_n687), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n692), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n917), .A2(new_n645), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT42), .Z(new_n939));
  OAI21_X1  g0739(.A(new_n589), .B1(new_n915), .B2(new_n488), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n940), .A2(new_n629), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT43), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n939), .A2(new_n941), .B1(new_n942), .B2(new_n911), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n911), .A2(new_n942), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n943), .B(new_n944), .Z(new_n945));
  NOR2_X1   g0745(.A1(new_n641), .A2(new_n917), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n912), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT106), .ZN(G387));
  OR2_X1    g0749(.A1(new_n928), .A2(new_n687), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(new_n650), .A3(new_n929), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n639), .A2(new_n699), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n229), .A2(new_n709), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT108), .Z(new_n954));
  NAND2_X1  g0754(.A1(new_n284), .A2(new_n422), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT50), .Z(new_n956));
  AOI211_X1 g0756(.A(G45), .B(new_n648), .C1(G68), .C2(G77), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n708), .B(new_n954), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n648), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n959), .A2(new_n704), .B1(G107), .B2(new_n209), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT107), .Z(new_n961));
  OAI21_X1  g0761(.A(new_n702), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n694), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n250), .B1(new_n719), .B2(new_n512), .C1(new_n367), .C2(new_n715), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT109), .B(G150), .Z(new_n965));
  OAI22_X1  g0765(.A1(new_n740), .A2(new_n965), .B1(new_n720), .B2(new_n324), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n422), .A2(new_n730), .B1(new_n728), .B2(new_n741), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n520), .A2(new_n723), .B1(new_n732), .B2(new_n304), .ZN(new_n968));
  OR4_X1    g0768(.A1(new_n964), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n724), .A2(G283), .B1(new_n716), .B2(new_n474), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G317), .A2(new_n772), .B1(new_n771), .B2(G322), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n889), .A2(new_n894), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(new_n745), .C2(new_n732), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT48), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT110), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(KEYINPUT49), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n719), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n250), .B1(new_n979), .B2(new_n441), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n978), .B(new_n980), .C1(new_n751), .C2(new_n740), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT49), .B1(new_n976), .B2(new_n977), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n969), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n963), .B1(new_n983), .B2(new_n701), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n928), .A2(new_n693), .B1(new_n952), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n951), .A2(new_n985), .ZN(G393));
  INV_X1    g0786(.A(new_n650), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n924), .B2(new_n930), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n924), .B2(new_n930), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n917), .A2(new_n699), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G311), .A2(new_n772), .B1(new_n771), .B2(G317), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT52), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n250), .B1(new_n979), .B2(G107), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n744), .B2(new_n715), .C1(new_n740), .C2(new_n753), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT112), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n732), .A2(new_n764), .B1(new_n538), .B2(new_n723), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G303), .B2(new_n889), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n992), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n278), .A2(new_n728), .B1(new_n730), .B2(new_n741), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT51), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n250), .B1(new_n719), .B2(new_n516), .C1(new_n723), .C2(new_n367), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n720), .A2(new_n422), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n284), .C2(new_n733), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n740), .A2(new_n903), .B1(new_n304), .B2(new_n715), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT111), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1000), .A2(new_n1003), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n757), .B1(new_n998), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n708), .A2(new_n239), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n703), .B(new_n1010), .C1(G97), .C2(new_n649), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1009), .A2(new_n695), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n924), .A2(new_n693), .B1(new_n990), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n989), .A2(new_n1013), .ZN(G390));
  INV_X1    g0814(.A(new_n861), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n685), .A2(new_n629), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n783), .A2(new_n392), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n781), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n828), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1015), .B(new_n822), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n861), .B1(new_n864), .B2(new_n828), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n859), .B(new_n858), .C1(new_n1021), .C2(KEYINPUT113), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1021), .A2(KEYINPUT113), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n828), .A2(new_n784), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n672), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1026), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1020), .B(new_n1028), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n440), .A2(new_n673), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n868), .A2(new_n621), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1019), .B1(new_n672), .B2(new_n786), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n864), .B1(new_n1034), .B2(new_n1026), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1028), .A2(new_n1018), .A3(new_n1033), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n987), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1027), .A2(new_n1029), .A3(new_n1037), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(G132), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n250), .B1(new_n422), .B2(new_n719), .C1(new_n730), .C2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT54), .B(G143), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n733), .B2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n965), .A2(new_n715), .A3(KEYINPUT53), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT53), .B1(new_n965), .B2(new_n715), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n741), .B2(new_n723), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(G128), .C2(new_n771), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n778), .A2(G125), .B1(G137), .B2(new_n889), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1045), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n740), .A2(new_n764), .B1(new_n304), .B2(new_n719), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT114), .Z(new_n1053));
  AOI22_X1  g0853(.A1(G116), .A2(new_n772), .B1(new_n771), .B2(G283), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n243), .B1(new_n715), .B2(new_n516), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G77), .B2(new_n724), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G97), .A2(new_n733), .B1(new_n889), .B2(G107), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1051), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n701), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n695), .B1(new_n324), .B2(new_n762), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n860), .C2(new_n698), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n1030), .B2(new_n692), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1041), .A2(new_n1063), .ZN(G378));
  NAND2_X1  g0864(.A1(new_n846), .A2(new_n851), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n287), .A2(new_n799), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n302), .B(new_n1066), .Z(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  AND4_X1   g0869(.A1(G330), .A2(new_n1065), .A3(new_n830), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n852), .B2(G330), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n867), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1070), .A2(new_n1071), .B1(KEYINPUT119), .B2(new_n1072), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n845), .A2(new_n832), .A3(KEYINPUT40), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT101), .B1(new_n849), .B2(new_n850), .ZN(new_n1075));
  OAI211_X1 g0875(.A(G330), .B(new_n830), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1069), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n852), .A2(G330), .A3(new_n1069), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1072), .A2(KEYINPUT119), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1073), .A2(new_n693), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n695), .B1(new_n422), .B2(new_n762), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n778), .A2(G283), .B1(new_n373), .B2(new_n733), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n979), .A2(G58), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT115), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(new_n512), .C2(new_n720), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n772), .A2(G107), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT116), .ZN(new_n1089));
  AOI211_X1 g0889(.A(G41), .B(new_n250), .C1(new_n716), .C2(G77), .ZN(new_n1090));
  INV_X1    g0890(.A(G116), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n902), .C1(new_n1091), .C2(new_n728), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1087), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT117), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1094), .A2(KEYINPUT58), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G132), .A2(new_n889), .B1(new_n733), .B2(G137), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n771), .A2(G125), .B1(new_n716), .B2(new_n1044), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n772), .A2(G128), .B1(G150), .B2(new_n724), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT59), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(KEYINPUT59), .ZN(new_n1101));
  AOI211_X1 g0901(.A(G33), .B(G41), .C1(new_n979), .C2(G159), .ZN(new_n1102));
  INV_X1    g0902(.A(G124), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n740), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT118), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1100), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n422), .B1(new_n241), .B2(G41), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1095), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(KEYINPUT58), .B2(new_n1094), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1083), .B1(new_n757), .B2(new_n1109), .C1(new_n1069), .C2(new_n698), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1082), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1032), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1040), .A2(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1073), .A2(new_n1113), .A3(new_n1081), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n650), .B1(new_n1114), .B2(KEYINPUT57), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(KEYINPUT57), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n867), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT120), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1078), .A2(new_n1118), .A3(new_n1079), .A4(new_n1072), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1078), .A2(new_n1072), .A3(new_n1079), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT120), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1116), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1111), .B1(new_n1115), .B2(new_n1123), .ZN(G375));
  AOI21_X1  g0924(.A(new_n692), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1019), .A2(new_n697), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n771), .A2(G294), .B1(new_n733), .B2(G107), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n538), .B2(new_n720), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT122), .Z(new_n1129));
  AOI21_X1  g0929(.A(new_n250), .B1(new_n979), .B2(G77), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n512), .B2(new_n715), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n740), .A2(new_n745), .B1(new_n520), .B2(new_n723), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(G283), .C2(new_n772), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n250), .B1(new_n715), .B2(new_n741), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1042), .A2(new_n728), .B1(new_n730), .B2(new_n900), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(G50), .C2(new_n724), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n778), .A2(G128), .B1(new_n889), .B2(new_n1044), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n733), .A2(G150), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1086), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n757), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n695), .B(new_n1141), .C1(new_n304), .C2(new_n762), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1125), .B1(new_n1126), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1038), .A2(new_n934), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT121), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1032), .A2(new_n1035), .A3(KEYINPUT121), .A4(new_n1036), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1143), .B1(new_n1144), .B2(new_n1149), .ZN(G381));
  NOR2_X1   g0950(.A1(G375), .A2(G378), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(G393), .A2(G396), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OR4_X1    g0954(.A1(G384), .A2(new_n1154), .A3(G390), .A4(G381), .ZN(new_n1155));
  OR3_X1    g0955(.A1(G387), .A2(new_n1152), .A3(new_n1155), .ZN(G407));
  OAI211_X1 g0956(.A(G407), .B(G213), .C1(G343), .C2(new_n1152), .ZN(G409));
  NOR2_X1   g0957(.A1(new_n1041), .A2(new_n1063), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n692), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1073), .A2(new_n1113), .A3(new_n934), .A4(new_n1081), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1110), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1158), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT123), .ZN(new_n1163));
  OAI211_X1 g0963(.A(G378), .B(new_n1111), .C1(new_n1115), .C2(new_n1123), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT123), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1158), .B(new_n1165), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n627), .A2(G213), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT60), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1037), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1149), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1032), .A2(new_n1035), .A3(KEYINPUT60), .A4(new_n1036), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT124), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT125), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1171), .A2(new_n1174), .A3(new_n1175), .A4(new_n650), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n650), .B1(new_n1149), .B2(new_n1170), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT125), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT126), .ZN(new_n1180));
  OR2_X1    g0980(.A1(G384), .A2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1181), .A2(new_n1143), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(G384), .A2(new_n1180), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1184), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1179), .A2(new_n1182), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1167), .A2(new_n1168), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT62), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1167), .A2(KEYINPUT62), .A3(new_n1168), .A4(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1168), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1194), .A2(G2897), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1185), .A2(new_n1187), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT61), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1193), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT127), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT106), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(G393), .A2(G396), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1203), .B1(new_n1205), .B2(new_n1153), .ZN(new_n1206));
  INV_X1    g1006(.A(G390), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(G390), .B1(new_n1205), .B2(new_n1153), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(new_n948), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT127), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1193), .A2(new_n1212), .A3(new_n1200), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1202), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT63), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1189), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1211), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1189), .A2(new_n1215), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1216), .A2(new_n1200), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1214), .A2(new_n1219), .ZN(G405));
  XNOR2_X1  g1020(.A(new_n1211), .B(new_n1188), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(G375), .A2(new_n1158), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1164), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1221), .B(new_n1223), .ZN(G402));
endmodule


