

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n418), .B(n417), .ZN(n534) );
  XNOR2_X1 U325 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n417) );
  AND2_X1 U326 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  NAND2_X1 U327 ( .A1(n559), .A2(n578), .ZN(n411) );
  XNOR2_X1 U328 ( .A(n378), .B(n292), .ZN(n379) );
  XNOR2_X1 U329 ( .A(n380), .B(n379), .ZN(n383) );
  XNOR2_X1 U330 ( .A(n455), .B(n454), .ZN(n569) );
  XOR2_X1 U331 ( .A(n470), .B(KEYINPUT28), .Z(n539) );
  XNOR2_X1 U332 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U333 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(G155GAT), .B(KEYINPUT3), .Z(n294) );
  XNOR2_X1 U335 ( .A(KEYINPUT91), .B(KEYINPUT2), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n326) );
  XOR2_X1 U337 ( .A(n326), .B(G162GAT), .Z(n296) );
  NAND2_X1 U338 ( .A1(G225GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U340 ( .A(G29GAT), .B(n297), .ZN(n313) );
  XOR2_X1 U341 ( .A(G85GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U342 ( .A(G141GAT), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U344 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n301) );
  XNOR2_X1 U345 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U348 ( .A(KEYINPUT86), .B(G134GAT), .Z(n305) );
  XNOR2_X1 U349 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U351 ( .A(G113GAT), .B(n306), .Z(n448) );
  XOR2_X1 U352 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n308) );
  XNOR2_X1 U353 ( .A(KEYINPUT93), .B(G57GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n448), .B(n309), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n523) );
  INV_X1 U358 ( .A(n523), .ZN(n575) );
  XOR2_X1 U359 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n315) );
  NAND2_X1 U360 ( .A1(G228GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U362 ( .A(n316), .B(KEYINPUT22), .Z(n325) );
  XNOR2_X1 U363 ( .A(G148GAT), .B(KEYINPUT73), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n317), .B(KEYINPUT74), .ZN(n318) );
  XOR2_X1 U365 ( .A(n318), .B(G204GAT), .Z(n320) );
  XNOR2_X1 U366 ( .A(G78GAT), .B(G106GAT), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n385) );
  XOR2_X1 U368 ( .A(KEYINPUT90), .B(G218GAT), .Z(n322) );
  XNOR2_X1 U369 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U371 ( .A(G197GAT), .B(n323), .Z(n431) );
  XNOR2_X1 U372 ( .A(n385), .B(n431), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n327) );
  XOR2_X1 U374 ( .A(n327), .B(n326), .Z(n329) );
  XOR2_X1 U375 ( .A(G141GAT), .B(G22GAT), .Z(n395) );
  XOR2_X1 U376 ( .A(G50GAT), .B(G162GAT), .Z(n333) );
  XNOR2_X1 U377 ( .A(n395), .B(n333), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n470) );
  AND2_X1 U379 ( .A1(n575), .A2(n470), .ZN(n435) );
  XOR2_X1 U380 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n331) );
  XNOR2_X1 U381 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n350) );
  XOR2_X1 U383 ( .A(G99GAT), .B(G85GAT), .Z(n373) );
  XNOR2_X1 U384 ( .A(G36GAT), .B(G190GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n332), .B(KEYINPUT79), .ZN(n423) );
  XNOR2_X1 U386 ( .A(n333), .B(n423), .ZN(n337) );
  INV_X1 U387 ( .A(n337), .ZN(n335) );
  AND2_X1 U388 ( .A1(G232GAT), .A2(G233GAT), .ZN(n336) );
  INV_X1 U389 ( .A(n336), .ZN(n334) );
  NAND2_X1 U390 ( .A1(n335), .A2(n334), .ZN(n339) );
  NAND2_X1 U391 ( .A1(n337), .A2(n336), .ZN(n338) );
  NAND2_X1 U392 ( .A1(n339), .A2(n338), .ZN(n341) );
  INV_X1 U393 ( .A(G92GAT), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U395 ( .A(G29GAT), .B(G43GAT), .Z(n343) );
  XNOR2_X1 U396 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n399) );
  XNOR2_X1 U398 ( .A(n399), .B(G106GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U400 ( .A(n373), .B(n346), .Z(n348) );
  XNOR2_X1 U401 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n462) );
  XNOR2_X1 U404 ( .A(KEYINPUT36), .B(n462), .ZN(n489) );
  XOR2_X1 U405 ( .A(KEYINPUT83), .B(KEYINPUT12), .Z(n352) );
  XNOR2_X1 U406 ( .A(G64GAT), .B(KEYINPUT85), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U408 ( .A(G155GAT), .B(G211GAT), .Z(n354) );
  XNOR2_X1 U409 ( .A(G127GAT), .B(G71GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n370) );
  XOR2_X1 U412 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n358) );
  XNOR2_X1 U413 ( .A(KEYINPUT82), .B(KEYINPUT84), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U415 ( .A(G8GAT), .B(G183GAT), .Z(n420) );
  XOR2_X1 U416 ( .A(n420), .B(G78GAT), .Z(n360) );
  XOR2_X1 U417 ( .A(G15GAT), .B(G1GAT), .Z(n394) );
  XNOR2_X1 U418 ( .A(G22GAT), .B(n394), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U420 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U423 ( .A(n365), .B(KEYINPUT81), .Z(n368) );
  XNOR2_X1 U424 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n366), .B(KEYINPUT70), .ZN(n384) );
  XNOR2_X1 U426 ( .A(n384), .B(KEYINPUT14), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n585) );
  NAND2_X1 U429 ( .A1(n489), .A2(n585), .ZN(n372) );
  XOR2_X1 U430 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n408) );
  XOR2_X1 U432 ( .A(KEYINPUT76), .B(KEYINPUT71), .Z(n375) );
  XOR2_X1 U433 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U434 ( .A(n441), .B(n373), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U436 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n377) );
  XNOR2_X1 U437 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U439 ( .A(KEYINPUT75), .B(G64GAT), .Z(n382) );
  XNOR2_X1 U440 ( .A(G176GAT), .B(G92GAT), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n419) );
  XOR2_X1 U442 ( .A(n383), .B(n419), .Z(n387) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n460) );
  INV_X1 U445 ( .A(n460), .ZN(n581) );
  XOR2_X1 U446 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n389) );
  XNOR2_X1 U447 ( .A(G113GAT), .B(G8GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U449 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n391) );
  XNOR2_X1 U450 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n406) );
  XOR2_X1 U453 ( .A(G36GAT), .B(G50GAT), .Z(n397) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U456 ( .A(n398), .B(G197GAT), .Z(n404) );
  XOR2_X1 U457 ( .A(n399), .B(KEYINPUT69), .Z(n401) );
  NAND2_X1 U458 ( .A1(G229GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U460 ( .A(G169GAT), .B(n402), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n578) );
  NOR2_X1 U463 ( .A1(n581), .A2(n578), .ZN(n407) );
  AND2_X1 U464 ( .A1(n408), .A2(n407), .ZN(n410) );
  INV_X1 U465 ( .A(KEYINPUT111), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n416) );
  XNOR2_X1 U467 ( .A(KEYINPUT41), .B(n460), .ZN(n559) );
  XNOR2_X1 U468 ( .A(n411), .B(KEYINPUT46), .ZN(n412) );
  INV_X1 U469 ( .A(n585), .ZN(n464) );
  NAND2_X1 U470 ( .A1(n412), .A2(n464), .ZN(n413) );
  NOR2_X1 U471 ( .A1(n462), .A2(n413), .ZN(n414) );
  XOR2_X1 U472 ( .A(KEYINPUT47), .B(n414), .Z(n415) );
  NOR2_X1 U473 ( .A1(n416), .A2(n415), .ZN(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT94), .B(n419), .Z(n422) );
  XNOR2_X1 U475 ( .A(G204GAT), .B(n420), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U477 ( .A(n423), .B(KEYINPUT95), .Z(n425) );
  NAND2_X1 U478 ( .A1(G226GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U480 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U481 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n429) );
  XNOR2_X1 U482 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U484 ( .A(G169GAT), .B(n430), .Z(n452) );
  XNOR2_X1 U485 ( .A(n452), .B(n431), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n511) );
  NOR2_X1 U487 ( .A1(n534), .A2(n511), .ZN(n434) );
  XNOR2_X1 U488 ( .A(KEYINPUT54), .B(n434), .ZN(n574) );
  NAND2_X1 U489 ( .A1(n435), .A2(n574), .ZN(n437) );
  XOR2_X1 U490 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n453) );
  XOR2_X1 U492 ( .A(G183GAT), .B(G176GAT), .Z(n439) );
  XNOR2_X1 U493 ( .A(G15GAT), .B(G190GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U495 ( .A(n440), .B(G99GAT), .Z(n443) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U498 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n445) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U501 ( .A(n447), .B(n446), .Z(n450) );
  XNOR2_X1 U502 ( .A(n448), .B(KEYINPUT88), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n537) );
  NAND2_X1 U505 ( .A1(n453), .A2(n537), .ZN(n455) );
  INV_X1 U506 ( .A(KEYINPUT122), .ZN(n454) );
  NAND2_X1 U507 ( .A1(n569), .A2(n559), .ZN(n459) );
  XOR2_X1 U508 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n457) );
  XNOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n460), .A2(n578), .ZN(n461) );
  XNOR2_X1 U511 ( .A(n461), .B(KEYINPUT77), .ZN(n494) );
  INV_X1 U512 ( .A(n462), .ZN(n463) );
  INV_X1 U513 ( .A(n463), .ZN(n568) );
  NOR2_X1 U514 ( .A1(n568), .A2(n464), .ZN(n465) );
  XNOR2_X1 U515 ( .A(KEYINPUT16), .B(n465), .ZN(n478) );
  INV_X1 U516 ( .A(n537), .ZN(n513) );
  XOR2_X1 U517 ( .A(n511), .B(KEYINPUT27), .Z(n472) );
  NAND2_X1 U518 ( .A1(n523), .A2(n472), .ZN(n535) );
  NOR2_X1 U519 ( .A1(n539), .A2(n535), .ZN(n466) );
  NAND2_X1 U520 ( .A1(n513), .A2(n466), .ZN(n477) );
  INV_X1 U521 ( .A(n511), .ZN(n525) );
  NAND2_X1 U522 ( .A1(n537), .A2(n525), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n467), .A2(n470), .ZN(n468) );
  XNOR2_X1 U524 ( .A(n468), .B(KEYINPUT96), .ZN(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(n469), .Z(n474) );
  NOR2_X1 U526 ( .A1(n537), .A2(n470), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n471), .B(KEYINPUT26), .ZN(n576) );
  NAND2_X1 U528 ( .A1(n472), .A2(n576), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n475), .A2(n575), .ZN(n476) );
  NAND2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n490) );
  AND2_X1 U532 ( .A1(n478), .A2(n490), .ZN(n508) );
  NAND2_X1 U533 ( .A1(n494), .A2(n508), .ZN(n486) );
  NOR2_X1 U534 ( .A1(n575), .A2(n486), .ZN(n479) );
  XOR2_X1 U535 ( .A(KEYINPUT34), .B(n479), .Z(n480) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n511), .A2(n486), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1325GAT) );
  NOR2_X1 U540 ( .A1(n513), .A2(n486), .ZN(n484) );
  XNOR2_X1 U541 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  INV_X1 U544 ( .A(n539), .ZN(n516) );
  NOR2_X1 U545 ( .A1(n516), .A2(n486), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  NAND2_X1 U549 ( .A1(n489), .A2(n490), .ZN(n491) );
  NOR2_X1 U550 ( .A1(n585), .A2(n491), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT37), .B(n492), .Z(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT100), .B(n493), .ZN(n520) );
  NAND2_X1 U553 ( .A1(n520), .A2(n494), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n495), .B(KEYINPUT38), .ZN(n496) );
  XNOR2_X1 U555 ( .A(KEYINPUT101), .B(n496), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n523), .A2(n503), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n503), .A2(n525), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n501) );
  NAND2_X1 U561 ( .A1(n503), .A2(n537), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U563 ( .A(G43GAT), .B(n502), .Z(G1330GAT) );
  XOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT103), .Z(n505) );
  NAND2_X1 U565 ( .A1(n539), .A2(n503), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  INV_X1 U567 ( .A(n578), .ZN(n506) );
  NAND2_X1 U568 ( .A1(n559), .A2(n506), .ZN(n507) );
  XOR2_X1 U569 ( .A(KEYINPUT104), .B(n507), .Z(n521) );
  NAND2_X1 U570 ( .A1(n508), .A2(n521), .ZN(n515) );
  NOR2_X1 U571 ( .A1(n575), .A2(n515), .ZN(n509) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n511), .A2(n515), .ZN(n512) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n513), .A2(n515), .ZN(n514) );
  XOR2_X1 U577 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X1 U579 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n519), .Z(G1335GAT) );
  NAND2_X1 U582 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U583 ( .A(KEYINPUT106), .B(n522), .Z(n530) );
  NAND2_X1 U584 ( .A1(n523), .A2(n530), .ZN(n524) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  XOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT107), .Z(n527) );
  NAND2_X1 U587 ( .A1(n530), .A2(n525), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n527), .B(n526), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n530), .A2(n537), .ZN(n528) );
  XNOR2_X1 U590 ( .A(n528), .B(KEYINPUT108), .ZN(n529) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n532) );
  NAND2_X1 U593 ( .A1(n539), .A2(n530), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n536), .B(KEYINPUT112), .ZN(n552) );
  NAND2_X1 U598 ( .A1(n537), .A2(n552), .ZN(n538) );
  NOR2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n549) );
  NAND2_X1 U600 ( .A1(n549), .A2(n578), .ZN(n540) );
  XOR2_X1 U601 ( .A(KEYINPUT113), .B(n540), .Z(n541) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n543) );
  NAND2_X1 U604 ( .A1(n549), .A2(n559), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n546) );
  NAND2_X1 U609 ( .A1(n549), .A2(n585), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n548), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U613 ( .A1(n549), .A2(n568), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n552), .A2(n576), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n553), .B(KEYINPUT117), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n563), .A2(n578), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n557) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(n558), .Z(n561) );
  NAND2_X1 U624 ( .A1(n563), .A2(n559), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n563), .A2(n585), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n568), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U630 ( .A(G169GAT), .B(KEYINPUT123), .Z(n566) );
  NAND2_X1 U631 ( .A1(n578), .A2(n569), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n585), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n571) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(G190GAT), .ZN(G1351GAT) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(KEYINPUT59), .ZN(n580) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n577) );
  AND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n587), .A2(n578), .ZN(n579) );
  XOR2_X1 U644 ( .A(n580), .B(n579), .Z(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n583) );
  NAND2_X1 U646 ( .A1(n587), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n587), .A2(n585), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n489), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

