//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT71), .B(KEYINPUT1), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT70), .ZN(new_n205));
  AND2_X1   g004(.A1(G127gat), .A2(G134gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G127gat), .A2(G134gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  INV_X1    g008(.A(G134gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G127gat), .A2(G134gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT70), .A3(new_n212), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n203), .A2(new_n204), .A3(new_n208), .A4(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(new_n206), .B2(new_n207), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(KEYINPUT69), .A3(new_n212), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n216), .B(new_n217), .C1(KEYINPUT1), .C2(new_n202), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n222), .A2(KEYINPUT26), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n223), .A2(KEYINPUT26), .ZN(new_n227));
  OR3_X1    g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT28), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT27), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT27), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n233));
  OAI211_X1 g032(.A(KEYINPUT67), .B(G183gat), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G183gat), .ZN(new_n235));
  AOI21_X1  g034(.A(G190gat), .B1(new_n235), .B2(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(KEYINPUT27), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n229), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  INV_X1    g042(.A(new_n236), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n232), .A2(G183gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT28), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n243), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n236), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n228), .B1(new_n242), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252));
  INV_X1    g051(.A(new_n223), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n222), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(KEYINPUT64), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n255), .A2(new_n226), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n255), .B(new_n226), .C1(KEYINPUT64), .C2(KEYINPUT24), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260));
  INV_X1    g059(.A(G190gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n235), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT24), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT65), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n262), .A2(new_n264), .A3(new_n225), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n225), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n265), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n253), .A2(new_n252), .ZN(new_n268));
  INV_X1    g067(.A(new_n222), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n258), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n259), .A2(new_n260), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n219), .B1(new_n251), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G227gat), .ZN(new_n274));
  INV_X1    g073(.A(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n260), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n267), .A2(new_n271), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n214), .A2(new_n218), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n244), .B1(new_n240), .B2(KEYINPUT67), .ZN(new_n281));
  OAI21_X1  g080(.A(G183gat), .B1(new_n231), .B2(new_n233), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n249), .B1(new_n285), .B2(new_n229), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n279), .B(new_n280), .C1(new_n286), .C2(new_n228), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n273), .A2(new_n276), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT33), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G15gat), .B(G43gat), .Z(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n294), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n288), .B(KEYINPUT32), .C1(new_n290), .C2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n273), .A2(new_n287), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n274), .B2(new_n275), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT34), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n298), .B(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT36), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n295), .A2(new_n304), .A3(new_n297), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n295), .B2(new_n297), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(KEYINPUT73), .B(new_n301), .C1(new_n305), .C2(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n300), .B(KEYINPUT34), .Z(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n298), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n313), .A2(KEYINPUT36), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n303), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G78gat), .B(G106gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(G22gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G197gat), .B(G204gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT22), .ZN(new_n320));
  INV_X1    g119(.A(G211gat), .ZN(new_n321));
  INV_X1    g120(.A(G218gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n319), .A3(new_n323), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(KEYINPUT80), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n323), .B2(new_n319), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT29), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT3), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n334), .A2(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G155gat), .ZN(new_n339));
  INV_X1    g138(.A(G162gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT2), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G141gat), .B(G148gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n334), .B1(G155gat), .B2(G162gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n337), .B(new_n335), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n333), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n328), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT74), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n345), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n351), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n327), .B2(new_n328), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n349), .B1(new_n361), .B2(KEYINPUT3), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n359), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT31), .B(G50gat), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n360), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n364), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n358), .A2(new_n362), .ZN(new_n367));
  INV_X1    g166(.A(new_n359), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n358), .A3(new_n359), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n318), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n364), .B1(new_n360), .B2(new_n363), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n370), .A3(new_n366), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n317), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G1gat), .B(G29gat), .Z(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G57gat), .B(G85gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n355), .A3(new_n280), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n219), .A2(new_n350), .A3(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n214), .A2(new_n218), .A3(new_n345), .A4(new_n348), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n280), .A2(new_n349), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n387), .ZN(new_n393));
  INV_X1    g192(.A(new_n386), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n391), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n382), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n390), .A2(new_n397), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n390), .A2(new_n395), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n381), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n381), .B1(new_n400), .B2(new_n401), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n404), .A2(KEYINPUT79), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n399), .A2(new_n402), .A3(new_n408), .A4(new_n403), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G8gat), .B(G36gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n353), .ZN(new_n416));
  INV_X1    g215(.A(G226gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(new_n275), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n251), .A2(new_n272), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(KEYINPUT29), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n279), .B1(new_n286), .B2(new_n228), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n418), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n416), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n418), .B1(new_n422), .B2(new_n356), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n242), .A2(new_n250), .ZN(new_n426));
  INV_X1    g225(.A(new_n228), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n419), .B1(new_n428), .B2(new_n279), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n425), .A2(new_n429), .A3(new_n353), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n415), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n421), .A2(new_n416), .A3(new_n423), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n353), .B1(new_n425), .B2(new_n429), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n414), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n432), .A2(new_n433), .A3(new_n436), .A4(new_n414), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n376), .B1(new_n411), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n435), .A2(KEYINPUT81), .A3(new_n437), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT81), .B1(new_n435), .B2(new_n437), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT39), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n385), .A2(new_n389), .ZN(new_n444));
  INV_X1    g243(.A(new_n384), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n443), .B(new_n394), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n444), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n386), .B1(new_n447), .B2(new_n384), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT39), .B1(new_n393), .B2(new_n394), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n381), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n406), .B1(new_n451), .B2(KEYINPUT40), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(KEYINPUT82), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT82), .B1(new_n450), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n441), .A2(new_n442), .A3(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n372), .A2(new_n375), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n432), .A2(new_n433), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n414), .B1(new_n460), .B2(KEYINPUT37), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT38), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n432), .A2(new_n433), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n406), .A2(new_n405), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n404), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n467), .A3(new_n434), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n462), .B1(new_n461), .B2(new_n464), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n459), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n440), .B1(new_n458), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n315), .A2(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n376), .A2(new_n467), .A3(KEYINPUT35), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n302), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n441), .A2(new_n442), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n407), .A2(new_n409), .B1(new_n435), .B2(new_n437), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n376), .B1(new_n312), .B2(new_n298), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n295), .A2(new_n297), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT72), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n295), .A2(new_n304), .A3(new_n297), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT73), .B1(new_n482), .B2(new_n301), .ZN(new_n483));
  INV_X1    g282(.A(new_n310), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n477), .B(new_n478), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n476), .B1(new_n486), .B2(KEYINPUT83), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n459), .A2(new_n313), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n309), .B2(new_n310), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n490), .B2(new_n477), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n472), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G113gat), .B(G141gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT85), .ZN(new_n496));
  XOR2_X1   g295(.A(G169gat), .B(G197gat), .Z(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n500), .B(KEYINPUT12), .Z(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT14), .B(G29gat), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G29gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(KEYINPUT86), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n508), .B2(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n507), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n504), .A2(new_n506), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT87), .B1(new_n508), .B2(KEYINPUT15), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n517), .A2(new_n518), .B1(new_n509), .B2(new_n511), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT16), .ZN(new_n523));
  AOI21_X1  g322(.A(G1gat), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n522), .B(new_n525), .C1(new_n523), .C2(G1gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT90), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n521), .A2(new_n529), .B1(new_n530), .B2(G8gat), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n529), .A2(new_n521), .A3(G8gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n520), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n521), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(G8gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n529), .A2(new_n521), .A3(G8gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n518), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n512), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n509), .A2(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n507), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n533), .A2(new_n542), .A3(KEYINPUT92), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT13), .Z(new_n545));
  NOR2_X1   g344(.A1(new_n531), .A2(new_n532), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n541), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n543), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT93), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n543), .A2(new_n548), .A3(new_n551), .A4(new_n545), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n539), .B(new_n554), .C1(new_n507), .C2(new_n540), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n556), .B(KEYINPUT17), .C1(new_n516), .C2(new_n519), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n541), .B2(KEYINPUT17), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n546), .B(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n544), .A3(new_n533), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT91), .B1(new_n520), .B2(new_n554), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n557), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n536), .A2(new_n555), .A3(new_n537), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n536), .A2(new_n537), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n565), .A2(new_n566), .B1(new_n520), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(KEYINPUT18), .A3(new_n544), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n501), .B1(new_n553), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n550), .A2(new_n552), .ZN(new_n572));
  INV_X1    g371(.A(new_n501), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n563), .A4(new_n569), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n494), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n339), .ZN(new_n578));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n578), .B(new_n579), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n582));
  XNOR2_X1  g381(.A(G71gat), .B(G78gat), .ZN(new_n583));
  INV_X1    g382(.A(G64gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n585));
  XOR2_X1   g384(.A(G57gat), .B(G64gat), .Z(new_n586));
  OAI211_X1 g385(.A(new_n583), .B(new_n585), .C1(new_n586), .C2(KEYINPUT96), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT95), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT97), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n588), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n587), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  OR3_X1    g394(.A1(KEYINPUT94), .A2(G71gat), .A3(G78gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n589), .B2(new_n586), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n582), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n586), .A2(KEYINPUT96), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n585), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n592), .A2(new_n593), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n588), .A2(new_n591), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT97), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n604), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n600), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(KEYINPUT98), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n601), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(G231gat), .A3(G233gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n601), .A2(new_n611), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(G127gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n595), .A2(new_n582), .A3(new_n600), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT98), .B1(new_n609), .B2(new_n610), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n601), .A2(new_n611), .A3(KEYINPUT99), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(KEYINPUT21), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n546), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n614), .A2(new_n209), .A3(new_n616), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n618), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n618), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n581), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n618), .A2(new_n626), .ZN(new_n630));
  INV_X1    g429(.A(new_n625), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n618), .A2(new_n625), .A3(new_n626), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n580), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT7), .ZN(new_n639));
  INV_X1    g438(.A(G85gat), .ZN(new_n640));
  OAI21_X1  g439(.A(G92gat), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G92gat), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n641), .A2(new_n643), .B1(new_n639), .B2(new_n640), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT8), .ZN(new_n645));
  NAND2_X1  g444(.A1(G99gat), .A2(G106gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(G99gat), .B(G106gat), .Z(new_n651));
  OAI21_X1  g450(.A(new_n638), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n644), .A2(new_n653), .A3(new_n649), .A4(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT102), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n644), .B2(new_n649), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n541), .ZN(new_n662));
  AND2_X1   g461(.A1(G232gat), .A2(G233gat), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(KEYINPUT41), .B2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n555), .B(new_n661), .C1(new_n558), .C2(new_n559), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n637), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n665), .A3(new_n637), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n663), .A2(KEYINPUT41), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G134gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n340), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n672), .B1(new_n666), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n667), .A2(new_n673), .A3(new_n668), .A4(new_n672), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT10), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n622), .A2(new_n623), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n661), .A2(new_n601), .A3(new_n611), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n650), .A2(new_n651), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n658), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n656), .A2(KEYINPUT104), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n684), .A2(new_n609), .A3(new_n610), .A4(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n681), .A2(new_n686), .A3(new_n678), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(G230gat), .A2(G233gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n681), .B2(new_n686), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(G120gat), .B(G148gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT105), .ZN(new_n694));
  XNOR2_X1  g493(.A(G176gat), .B(G204gat), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n694), .B(new_n695), .Z(new_n696));
  NAND3_X1  g495(.A1(new_n690), .A2(new_n692), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n696), .ZN(new_n698));
  INV_X1    g497(.A(new_n689), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n680), .B2(new_n687), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n700), .B2(new_n691), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT106), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n697), .A2(KEYINPUT106), .A3(new_n701), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n635), .A2(new_n677), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n576), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n411), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g509(.A(KEYINPUT16), .B(G8gat), .Z(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n475), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n475), .ZN(new_n713));
  OAI21_X1  g512(.A(G8gat), .B1(new_n707), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  MUX2_X1   g514(.A(new_n712), .B(new_n715), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g515(.A(new_n315), .ZN(new_n717));
  OAI21_X1  g516(.A(G15gat), .B1(new_n707), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n302), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(G15gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n707), .B2(new_n720), .ZN(G1326gat));
  NOR3_X1   g520(.A1(new_n494), .A2(new_n575), .A3(new_n459), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n706), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT107), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT43), .B(G22gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  NAND2_X1  g525(.A1(new_n703), .A2(new_n704), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(new_n635), .A3(new_n677), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n576), .A2(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(G29gat), .A3(new_n410), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n494), .B2(new_n677), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n458), .A2(new_n470), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n311), .A2(new_n314), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n735), .B(new_n440), .C1(new_n303), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n713), .A2(new_n302), .A3(new_n473), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n491), .B2(new_n492), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n677), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(KEYINPUT44), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n727), .B(KEYINPUT109), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n575), .A3(new_n635), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n734), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G29gat), .B1(new_n747), .B2(new_n410), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n748), .ZN(G1328gat));
  OAI21_X1  g548(.A(G36gat), .B1(new_n747), .B2(new_n713), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n576), .A2(new_n503), .A3(new_n475), .A4(new_n728), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n750), .B(new_n754), .C1(new_n752), .C2(new_n751), .ZN(G1329gat));
  NOR2_X1   g554(.A1(new_n729), .A2(new_n719), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n315), .A2(G43gat), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n756), .A2(G43gat), .B1(new_n747), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g558(.A1(new_n734), .A2(new_n743), .A3(new_n376), .A4(new_n746), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT111), .B1(new_n760), .B2(G50gat), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n727), .A2(new_n635), .A3(new_n677), .A4(G50gat), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n760), .A2(G50gat), .B1(new_n722), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n763), .B(new_n765), .ZN(G1331gat));
  NAND2_X1  g565(.A1(new_n571), .A2(new_n574), .ZN(new_n767));
  INV_X1    g566(.A(new_n635), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n744), .A2(new_n767), .A3(new_n742), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n741), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n410), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g571(.A(new_n770), .B(KEYINPUT112), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n713), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT113), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n773), .A2(new_n777), .A3(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n584), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n776), .A2(new_n780), .A3(new_n584), .A4(new_n778), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1333gat));
  NAND3_X1  g583(.A1(new_n773), .A2(G71gat), .A3(new_n315), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n719), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(G71gat), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n376), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G78gat), .ZN(G1335gat));
  AND3_X1   g589(.A1(new_n697), .A2(KEYINPUT106), .A3(new_n701), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n702), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n487), .A2(new_n493), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n677), .B1(new_n793), .B2(new_n737), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n767), .A2(new_n635), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT51), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AND4_X1   g596(.A1(KEYINPUT51), .A2(new_n741), .A3(new_n742), .A4(new_n795), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n792), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n640), .A3(new_n411), .ZN(new_n801));
  INV_X1    g600(.A(new_n795), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n792), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n734), .A2(new_n743), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT114), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n734), .A2(new_n743), .A3(new_n806), .A4(new_n803), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n805), .A2(new_n411), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n801), .B1(new_n808), .B2(new_n640), .ZN(G1336gat));
  OAI21_X1  g608(.A(G92gat), .B1(new_n804), .B2(new_n713), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n713), .A2(G92gat), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n745), .B(new_n811), .C1(new_n796), .C2(new_n798), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n805), .A2(new_n475), .A3(new_n807), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(G92gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n812), .A2(KEYINPUT115), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(G92gat), .B2(new_n815), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n818), .B2(new_n820), .ZN(G1337gat));
  INV_X1    g620(.A(G99gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n800), .A2(new_n822), .A3(new_n302), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n805), .A2(new_n315), .A3(new_n807), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n822), .ZN(G1338gat));
  NAND3_X1  g624(.A1(new_n805), .A2(new_n376), .A3(new_n807), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n744), .B1(new_n797), .B2(new_n799), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n459), .A2(G106gat), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n826), .A2(G106gat), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n804), .A2(new_n459), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(G106gat), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n745), .B(new_n828), .C1(new_n796), .C2(new_n798), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n830), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n829), .A2(new_n830), .B1(new_n832), .B2(new_n834), .ZN(G1339gat));
  NAND3_X1  g634(.A1(new_n680), .A2(new_n687), .A3(new_n699), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n690), .A2(KEYINPUT54), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n838));
  AOI21_X1  g637(.A(new_n696), .B1(new_n700), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(KEYINPUT55), .A3(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n697), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n680), .A2(new_n699), .A3(new_n687), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n843), .A2(new_n700), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n688), .A2(new_n689), .A3(new_n838), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n698), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n842), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n767), .A2(new_n841), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n568), .A2(new_n544), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n545), .B1(new_n543), .B2(new_n548), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n500), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n574), .B(new_n852), .C1(new_n791), .C2(new_n702), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n742), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n848), .A2(new_n697), .A3(new_n840), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n574), .A2(new_n675), .A3(new_n676), .A4(new_n852), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n768), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT116), .B1(new_n705), .B2(new_n767), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n629), .A2(new_n634), .B1(new_n675), .B2(new_n676), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n575), .A2(new_n860), .A3(new_n861), .A4(new_n792), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n410), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n864), .A2(new_n713), .A3(new_n490), .ZN(new_n865));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865), .B2(new_n767), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n853), .B1(new_n575), .B2(new_n855), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n857), .B1(new_n867), .B2(new_n677), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n868), .B2(new_n635), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT118), .B1(new_n869), .B2(new_n459), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n719), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n475), .A2(new_n410), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n459), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n767), .A2(G113gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n866), .B1(new_n875), .B2(new_n876), .ZN(G1340gat));
  OAI21_X1  g676(.A(G120gat), .B1(new_n874), .B2(new_n744), .ZN(new_n878));
  INV_X1    g677(.A(G120gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n865), .A2(new_n879), .A3(new_n727), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n881), .B(new_n882), .ZN(G1341gat));
  OAI21_X1  g682(.A(G127gat), .B1(new_n874), .B2(new_n768), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n865), .A2(new_n209), .A3(new_n635), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(G1342gat));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n210), .A3(new_n742), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT56), .Z(new_n890));
  OAI21_X1  g689(.A(G134gat), .B1(new_n874), .B2(new_n677), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1343gat));
  NAND2_X1  g691(.A1(new_n717), .A2(new_n872), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n869), .A2(new_n376), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n459), .B1(new_n858), .B2(new_n863), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n893), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G141gat), .B1(new_n900), .B2(new_n575), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n315), .A2(new_n459), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n713), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n864), .A2(new_n905), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n906), .A2(G141gat), .A3(new_n575), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n902), .A2(new_n908), .A3(KEYINPUT58), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n901), .B(new_n907), .C1(KEYINPUT121), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1344gat));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G148gat), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(new_n899), .B2(new_n727), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n917), .A2(new_n869), .A3(KEYINPUT57), .A4(new_n376), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n705), .A2(new_n767), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n459), .B1(new_n858), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n921), .B2(KEYINPUT57), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n918), .B1(new_n922), .B2(new_n898), .ZN(new_n923));
  INV_X1    g722(.A(new_n893), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n727), .ZN(new_n925));
  OAI21_X1  g724(.A(G148gat), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n916), .B1(new_n926), .B2(KEYINPUT59), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n906), .A2(G148gat), .A3(new_n792), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n913), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n928), .ZN(new_n930));
  INV_X1    g729(.A(new_n925), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n848), .A2(new_n697), .A3(new_n840), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n574), .A2(new_n852), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n932), .A2(new_n767), .B1(new_n727), .B2(new_n933), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n934), .A2(new_n742), .B1(new_n855), .B2(new_n856), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n919), .B1(new_n935), .B2(new_n768), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n895), .B1(new_n936), .B2(new_n459), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n937), .A2(new_n917), .B1(KEYINPUT57), .B2(new_n897), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n931), .B1(new_n938), .B2(new_n918), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n914), .B1(new_n939), .B2(G148gat), .ZN(new_n940));
  OAI211_X1 g739(.A(KEYINPUT123), .B(new_n930), .C1(new_n940), .C2(new_n916), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n929), .A2(new_n941), .ZN(G1345gat));
  OAI21_X1  g741(.A(G155gat), .B1(new_n900), .B2(new_n768), .ZN(new_n943));
  INV_X1    g742(.A(new_n906), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n339), .A3(new_n635), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1346gat));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n340), .A3(new_n742), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT124), .ZN(new_n948));
  OAI21_X1  g747(.A(G162gat), .B1(new_n900), .B2(new_n677), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(KEYINPUT125), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1347gat));
  NOR2_X1   g753(.A1(new_n713), .A2(new_n411), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n871), .A2(new_n873), .A3(new_n955), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n956), .A2(new_n220), .A3(new_n575), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n411), .B1(new_n858), .B2(new_n863), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(new_n475), .A3(new_n490), .ZN(new_n959));
  AOI21_X1  g758(.A(G169gat), .B1(new_n959), .B2(new_n767), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n957), .A2(new_n960), .ZN(G1348gat));
  OAI21_X1  g760(.A(G176gat), .B1(new_n956), .B2(new_n744), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(new_n221), .A3(new_n727), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n964), .B(new_n965), .ZN(G1349gat));
  OAI21_X1  g765(.A(G183gat), .B1(new_n956), .B2(new_n768), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n235), .A2(KEYINPUT27), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n959), .A2(new_n968), .A3(new_n245), .A4(new_n635), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g770(.A1(new_n959), .A2(new_n261), .A3(new_n742), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n956), .A2(new_n677), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n973), .A2(new_n974), .A3(G190gat), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n973), .B2(G190gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(G1351gat));
  AND3_X1   g776(.A1(new_n958), .A2(new_n475), .A3(new_n903), .ZN(new_n978));
  AOI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n767), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n717), .A2(new_n955), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n923), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n767), .A2(G197gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1352gat));
  INV_X1    g782(.A(new_n981), .ZN(new_n984));
  OAI21_X1  g783(.A(G204gat), .B1(new_n984), .B2(new_n744), .ZN(new_n985));
  INV_X1    g784(.A(G204gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n978), .A2(new_n986), .A3(new_n727), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT62), .Z(new_n988));
  NAND2_X1  g787(.A1(new_n985), .A2(new_n988), .ZN(G1353gat));
  NAND3_X1  g788(.A1(new_n978), .A2(new_n321), .A3(new_n635), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT63), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n991), .A2(KEYINPUT127), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n981), .A2(new_n635), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n321), .B1(KEYINPUT127), .B2(new_n991), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(new_n992), .ZN(new_n996));
  INV_X1    g795(.A(new_n994), .ZN(new_n997));
  AOI211_X1 g796(.A(new_n996), .B(new_n997), .C1(new_n981), .C2(new_n635), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n990), .B1(new_n995), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n984), .B2(new_n677), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n978), .A2(new_n322), .A3(new_n742), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


