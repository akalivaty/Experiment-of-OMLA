//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT85), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(KEYINPUT81), .B(KEYINPUT1), .C1(new_n194), .C2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT81), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n193), .A2(new_n195), .A3(new_n201), .A4(G128), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n205), .A2(KEYINPUT80), .A3(new_n201), .A4(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n208), .A2(new_n213), .A3(new_n209), .A4(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n209), .A2(G104), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n212), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G107), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n219), .B2(new_n215), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n207), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n207), .B2(new_n221), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n191), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G134), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G137), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n228), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT11), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(KEYINPUT11), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n227), .A2(G134), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n226), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n233), .A2(new_n226), .A3(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n217), .A2(new_n220), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n202), .B1(new_n246), .B2(new_n205), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT10), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n244), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G101), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT79), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n255), .A3(G101), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n193), .A2(new_n195), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n193), .A2(new_n195), .A3(new_n259), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n215), .B1(new_n210), .B2(KEYINPUT3), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n212), .B1(new_n264), .B2(new_n214), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n250), .B1(new_n257), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n225), .A2(new_n243), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G227), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT77), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n243), .B1(new_n225), .B2(new_n267), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n268), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n207), .A2(new_n221), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT82), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n207), .A2(new_n221), .A3(new_n222), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n281), .A2(new_n282), .B1(new_n248), .B2(new_n244), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n279), .B1(new_n283), .B2(new_n243), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n244), .A2(new_n248), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n223), .B2(new_n224), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT84), .A3(KEYINPUT12), .A4(new_n242), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(KEYINPUT12), .A3(new_n242), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n278), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n190), .B(new_n277), .C1(new_n292), .C2(new_n273), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n284), .A3(new_n287), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n273), .B1(new_n294), .B2(new_n268), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT85), .B1(new_n295), .B2(new_n276), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n296), .A3(G469), .ZN(new_n297));
  INV_X1    g111(.A(G469), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT86), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n274), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n268), .A2(KEYINPUT86), .A3(new_n273), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n294), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n275), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n273), .B1(new_n305), .B2(new_n268), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n300), .B1(new_n308), .B2(new_n298), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n189), .B1(new_n297), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G125), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n247), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n314), .B2(new_n262), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n269), .A2(G224), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G110), .B(G122), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(KEYINPUT2), .A2(G113), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT2), .A2(G113), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(KEYINPUT68), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(KEYINPUT68), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G116), .B(G119), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n322), .B(KEYINPUT68), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n321), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n251), .A2(new_n263), .A3(G101), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n255), .B2(new_n265), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n335), .B2(new_n253), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n326), .A2(KEYINPUT5), .ZN(new_n337));
  INV_X1    g151(.A(G113), .ZN(new_n338));
  INV_X1    g152(.A(G116), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G119), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  AND4_X1   g157(.A1(new_n330), .A2(new_n343), .A3(new_n217), .A4(new_n220), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n320), .B1(new_n336), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n263), .A2(new_n265), .B1(new_n328), .B2(new_n330), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n257), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n319), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(KEYINPUT6), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n257), .A2(new_n346), .ZN(new_n351));
  INV_X1    g165(.A(new_n344), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n319), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR4_X1   g169(.A1(new_n347), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n319), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n318), .B(new_n349), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n317), .A2(KEYINPUT7), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n316), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT89), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n316), .A2(new_n358), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT89), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n316), .A2(new_n362), .A3(new_n358), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n319), .B(KEYINPUT8), .Z(new_n365));
  NAND2_X1  g179(.A1(new_n342), .A2(KEYINPUT88), .ZN(new_n366));
  INV_X1    g180(.A(G119), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G116), .ZN(new_n368));
  OAI21_X1  g182(.A(G113), .B1(new_n368), .B2(KEYINPUT5), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n337), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n244), .B1(new_n330), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n330), .A2(new_n343), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n365), .B(new_n373), .C1(new_n244), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n364), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(G902), .B1(new_n376), .B2(new_n348), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n357), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G210), .B1(G237), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n357), .A2(new_n377), .A3(new_n379), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n313), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n269), .A2(G952), .ZN(new_n384));
  NAND2_X1  g198(.A1(G234), .A2(G237), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(G902), .A3(G953), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT21), .B(G898), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n194), .A2(G128), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n245), .A2(G143), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n393), .A2(new_n394), .A3(new_n229), .ZN(new_n395));
  INV_X1    g209(.A(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G116), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n339), .A2(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n398), .A3(new_n209), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n393), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n394), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n393), .A2(new_n403), .ZN(new_n406));
  OAI21_X1  g220(.A(G134), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n339), .A2(KEYINPUT14), .A3(G122), .ZN(new_n409));
  OAI211_X1 g223(.A(G107), .B(new_n409), .C1(new_n399), .C2(KEYINPUT14), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n229), .B1(new_n393), .B2(new_n394), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n410), .B(new_n401), .C1(new_n395), .C2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G217), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n187), .A2(new_n413), .A3(G953), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n408), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(new_n408), .B2(new_n412), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT93), .B1(new_n417), .B2(G902), .ZN(new_n418));
  INV_X1    g232(.A(G478), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(KEYINPUT15), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n408), .A2(new_n412), .ZN(new_n421));
  INV_X1    g235(.A(new_n414), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n408), .A2(new_n412), .A3(new_n414), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT93), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n299), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n420), .A3(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n425), .B(new_n299), .C1(KEYINPUT15), .C2(new_n419), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT94), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n430), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n194), .A2(KEYINPUT90), .ZN(new_n434));
  NOR2_X1   g248(.A1(G237), .A2(G953), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(G214), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT90), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G143), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n439), .A2(new_n434), .B1(new_n435), .B2(G214), .ZN(new_n440));
  OAI211_X1 g254(.A(KEYINPUT18), .B(G131), .C1(new_n437), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT18), .A2(G131), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT90), .B(G143), .ZN(new_n443));
  INV_X1    g257(.A(G214), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n444), .A2(G237), .A3(G953), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n436), .B(new_n442), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G125), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n314), .A2(G140), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G146), .ZN(new_n451));
  XNOR2_X1  g265(.A(G125), .B(G140), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n192), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n441), .A2(new_n446), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G131), .B1(new_n437), .B2(new_n440), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT17), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n436), .B(new_n226), .C1(new_n443), .C2(new_n445), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(KEYINPUT17), .B(G131), .C1(new_n437), .C2(new_n440), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT16), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n447), .A3(G125), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n450), .B2(new_n461), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n192), .ZN(new_n464));
  OAI211_X1 g278(.A(G146), .B(new_n462), .C1(new_n450), .C2(new_n461), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n460), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n455), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(G113), .B(G122), .Z(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT91), .B(G104), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT92), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n299), .B1(new_n467), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g289(.A(G475), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n452), .B(KEYINPUT19), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n192), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n456), .A2(new_n458), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n465), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n454), .A2(new_n446), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n470), .B1(new_n481), .B2(new_n441), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n467), .A2(new_n470), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n476), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n433), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n383), .A2(new_n392), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n311), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n413), .B1(G234), .B2(new_n299), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT75), .B1(new_n367), .B2(G128), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n493), .A2(KEYINPUT23), .B1(new_n367), .B2(G128), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(KEYINPUT23), .B2(new_n493), .ZN(new_n495));
  XNOR2_X1  g309(.A(G119), .B(G128), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT24), .B(G110), .Z(new_n497));
  OAI22_X1  g311(.A1(new_n495), .A2(G110), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n465), .A3(new_n453), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n464), .A2(new_n465), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(G110), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n496), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT76), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n499), .A2(KEYINPUT76), .A3(new_n503), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT22), .B(G137), .Z(new_n507));
  AND3_X1   g321(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  AOI211_X1 g325(.A(KEYINPUT76), .B(new_n510), .C1(new_n499), .C2(new_n503), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT25), .B1(new_n514), .B2(new_n299), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n516), .B(G902), .C1(new_n511), .C2(new_n513), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n492), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n492), .A2(G902), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(G472), .A2(G902), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n241), .A2(new_n247), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT66), .B1(new_n227), .B2(G134), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT66), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n229), .A3(G137), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n527), .A3(new_n237), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G131), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(KEYINPUT67), .A3(G131), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n524), .A2(KEYINPUT69), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n241), .A2(new_n532), .A3(new_n247), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT67), .B1(new_n528), .B2(G131), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n331), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n258), .A2(new_n259), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n196), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n205), .A2(new_n259), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n232), .B1(new_n230), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n229), .A2(G137), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n237), .B2(new_n235), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n544), .A2(new_n546), .A3(G131), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n542), .B1(new_n547), .B2(new_n239), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n533), .A2(new_n537), .A3(new_n538), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(G101), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n435), .A2(G210), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT71), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n551), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n551), .A3(new_n556), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n550), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  INV_X1    g375(.A(new_n550), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n561), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n549), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT64), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n260), .B2(new_n261), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT64), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(new_n547), .C2(new_n239), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n531), .A2(new_n532), .A3(new_n247), .A4(new_n241), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n533), .A2(new_n537), .A3(new_n548), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(KEYINPUT30), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n565), .B(new_n566), .C1(new_n575), .C2(new_n538), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT72), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n548), .B1(new_n572), .B2(new_n534), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n241), .A2(new_n532), .A3(new_n247), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT69), .B1(new_n580), .B2(new_n531), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT30), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n573), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n331), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(KEYINPUT72), .A3(new_n566), .A4(new_n565), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT28), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n570), .A2(new_n572), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n331), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n549), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n331), .B1(new_n242), .B2(new_n542), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT28), .B1(new_n592), .B2(new_n572), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n564), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n565), .B1(new_n575), .B2(new_n538), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(KEYINPUT31), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n523), .B1(new_n587), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT73), .B1(new_n598), .B2(KEYINPUT32), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT73), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT32), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n595), .B1(new_n591), .B2(new_n593), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n549), .A2(new_n564), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n584), .B2(new_n331), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n602), .B1(new_n604), .B2(new_n566), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n578), .B2(new_n586), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n600), .B(new_n601), .C1(new_n606), .C2(new_n523), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n523), .A2(new_n601), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT74), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n587), .A2(new_n597), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT74), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(new_n609), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n574), .A2(new_n331), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n549), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n593), .B1(new_n616), .B2(KEYINPUT28), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT29), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n595), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n575), .A2(new_n538), .ZN(new_n621));
  INV_X1    g435(.A(new_n549), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n595), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n618), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n594), .A2(new_n595), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n620), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G472), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n611), .A2(new_n614), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n521), .B1(new_n608), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n491), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT95), .B(G101), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G3));
  INV_X1    g446(.A(G472), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n612), .B2(new_n299), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n598), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G472), .B1(new_n606), .B2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n311), .A2(new_n639), .A3(new_n521), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n383), .A2(new_n392), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n418), .A2(new_n419), .A3(new_n427), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT33), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n423), .B2(new_n424), .ZN(new_n645));
  OAI211_X1 g459(.A(G478), .B(new_n299), .C1(new_n643), .C2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n488), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n640), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT97), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  INV_X1    g468(.A(G475), .ZN(new_n655));
  INV_X1    g469(.A(new_n475), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(new_n473), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n431), .A2(new_n432), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(KEYINPUT98), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n486), .A2(new_n487), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n660), .B1(new_n661), .B2(KEYINPUT98), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n658), .A2(new_n392), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n381), .A2(new_n382), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n312), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n640), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT100), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT35), .B(G107), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NAND2_X1  g487(.A1(new_n506), .A2(new_n510), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n504), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n299), .B1(new_n675), .B2(new_n512), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n516), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n514), .A2(KEYINPUT25), .A3(new_n299), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n499), .A2(new_n503), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n679), .A2(new_n492), .B1(new_n519), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n490), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n310), .A3(new_n638), .A4(new_n636), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G12));
  NAND2_X1  g501(.A1(new_n682), .A2(new_n519), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n518), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n599), .A2(new_n607), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n611), .A2(new_n614), .A3(new_n627), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n386), .B1(G900), .B2(new_n388), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n433), .A2(new_n662), .A3(new_n476), .A4(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n668), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n310), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n245), .ZN(G30));
  XNOR2_X1  g512(.A(new_n693), .B(KEYINPUT39), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n310), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n667), .B(new_n702), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n518), .A2(new_n433), .A3(new_n488), .A4(new_n688), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n703), .A2(new_n312), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT40), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n310), .A2(new_n706), .A3(new_n699), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n613), .B1(new_n612), .B2(new_n609), .ZN(new_n708));
  AOI211_X1 g522(.A(KEYINPUT74), .B(new_n610), .C1(new_n587), .C2(new_n597), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n621), .A2(new_n622), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n595), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n299), .B1(new_n616), .B2(new_n564), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n710), .A2(new_n599), .A3(new_n607), .A4(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n701), .A2(new_n705), .A3(new_n707), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  AND3_X1   g531(.A1(new_n488), .A2(new_n647), .A3(new_n693), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n357), .A2(new_n377), .A3(new_n379), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n379), .B1(new_n357), .B2(new_n377), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n718), .B(new_n312), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n667), .A2(KEYINPUT102), .A3(new_n312), .A4(new_n718), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n310), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n692), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n192), .ZN(G48));
  AND3_X1   g542(.A1(new_n268), .A2(KEYINPUT86), .A3(new_n273), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT86), .B1(new_n268), .B2(new_n273), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n306), .B1(new_n731), .B2(new_n294), .ZN(new_n732));
  OAI21_X1  g546(.A(G469), .B1(new_n732), .B2(G902), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n304), .A2(new_n307), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n298), .A3(new_n299), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n188), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n629), .A2(new_n650), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND3_X1  g554(.A1(new_n629), .A2(new_n669), .A3(new_n737), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT103), .B(G116), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G18));
  OR2_X1    g557(.A1(new_n736), .A2(new_n490), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n692), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  XNOR2_X1  g560(.A(KEYINPUT104), .B(G472), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n606), .B2(G902), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n535), .A2(new_n536), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n749), .A2(KEYINPUT69), .B1(new_n242), .B2(new_n542), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n538), .B1(new_n750), .B2(new_n537), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT28), .B1(new_n751), .B2(new_n622), .ZN(new_n752));
  INV_X1    g566(.A(new_n593), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n754), .A2(new_n595), .B1(KEYINPUT31), .B2(new_n596), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n587), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n522), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n521), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n736), .A2(new_n391), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n383), .A2(new_n433), .A3(new_n488), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G122), .ZN(G24));
  INV_X1    g578(.A(new_n747), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n612), .B2(new_n299), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n523), .B1(new_n587), .B2(new_n755), .ZN(new_n767));
  INV_X1    g581(.A(new_n718), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n766), .A2(new_n683), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n383), .A2(new_n733), .A3(new_n188), .A4(new_n735), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G125), .ZN(G27));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  OAI211_X1 g587(.A(G469), .B(new_n277), .C1(new_n292), .C2(new_n273), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n300), .B(KEYINPUT105), .Z(new_n775));
  NAND3_X1  g589(.A1(new_n735), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n719), .A2(new_n720), .A3(new_n313), .A4(new_n189), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n773), .A2(new_n776), .A3(new_n718), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n710), .A2(new_n599), .A3(new_n607), .A4(new_n627), .ZN(new_n779));
  INV_X1    g593(.A(new_n521), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n627), .B1(new_n606), .B2(new_n610), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n598), .A2(KEYINPUT32), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n776), .A2(new_n718), .A3(new_n777), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT42), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n226), .ZN(G33));
  NAND2_X1  g602(.A1(new_n694), .A2(KEYINPUT106), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT106), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n658), .A2(new_n790), .A3(new_n662), .A4(new_n693), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n776), .A2(new_n789), .A3(new_n777), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n779), .A2(new_n792), .A3(new_n780), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  NAND3_X1  g608(.A1(new_n381), .A2(new_n312), .A3(new_n382), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT109), .Z(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n647), .B(new_n476), .C1(new_n487), .C2(new_n486), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n689), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n639), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n797), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n801), .B1(new_n636), .B2(new_n638), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT44), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n807), .B1(new_n806), .B2(KEYINPUT44), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n293), .B2(new_n296), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n277), .B1(new_n292), .B2(new_n273), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n814));
  OAI21_X1  g628(.A(G469), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n775), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT46), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(KEYINPUT46), .B(new_n775), .C1(new_n812), .C2(new_n815), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n735), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n188), .A3(new_n699), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT107), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n735), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n816), .B2(new_n817), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n189), .B1(new_n825), .B2(new_n819), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(KEYINPUT107), .A3(new_n699), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n811), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(KEYINPUT110), .B(G137), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(G39));
  NOR4_X1   g644(.A1(new_n779), .A2(new_n780), .A3(new_n768), .A4(new_n795), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n826), .A2(KEYINPUT47), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n820), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g648(.A(KEYINPUT111), .B(G140), .Z(new_n835));
  XNOR2_X1  g649(.A(new_n834), .B(new_n835), .ZN(G42));
  NAND2_X1  g650(.A1(new_n188), .A2(new_n312), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n703), .A2(new_n521), .A3(new_n798), .A4(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n733), .A2(new_n735), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT49), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n611), .A2(new_n614), .A3(new_n714), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n690), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT112), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n693), .A2(new_n188), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n776), .A2(new_n704), .A3(new_n383), .A4(new_n846), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n692), .A2(new_n726), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n771), .B1(new_n692), .B2(new_n696), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT52), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n781), .A2(new_n793), .A3(new_n786), .ZN(new_n851));
  INV_X1    g665(.A(new_n795), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n428), .A2(new_n429), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n853), .A2(new_n476), .A3(new_n693), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n852), .A2(new_n662), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n779), .A2(new_n310), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n785), .A2(new_n758), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n689), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n850), .A2(new_n851), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n630), .A2(new_n745), .A3(new_n685), .A4(new_n763), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n629), .B(new_n737), .C1(new_n650), .C2(new_n669), .ZN(new_n862));
  INV_X1    g676(.A(new_n639), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n853), .A2(new_n488), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n648), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n641), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n863), .A2(new_n780), .A3(new_n310), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n683), .B1(new_n608), .B2(new_n628), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n310), .A2(new_n725), .ZN(new_n871));
  INV_X1    g685(.A(new_n847), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n870), .A2(new_n871), .B1(new_n715), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n748), .A2(new_n689), .A3(new_n757), .A4(new_n718), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n874), .A2(new_n668), .A3(new_n736), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n310), .A2(new_n695), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n869), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n850), .A3(new_n851), .A4(new_n859), .ZN(new_n882));
  INV_X1    g696(.A(new_n763), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n629), .B2(new_n491), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n685), .B1(new_n692), .B2(new_n744), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n884), .A2(new_n886), .A3(new_n862), .A4(new_n867), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n881), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  MUX2_X1   g703(.A(new_n845), .B(KEYINPUT54), .S(new_n889), .Z(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n737), .A2(new_n852), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT115), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n780), .A3(new_n387), .A4(new_n842), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n894), .A2(new_n488), .A3(new_n647), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT114), .ZN(new_n896));
  OR3_X1    g710(.A1(new_n703), .A2(new_n312), .A3(new_n736), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n800), .A2(new_n387), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n759), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT50), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n893), .A2(new_n898), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n902), .A2(KEYINPUT116), .A3(new_n683), .A4(new_n758), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n904));
  INV_X1    g718(.A(new_n902), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n758), .A2(new_n683), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n895), .B(new_n901), .C1(new_n903), .C2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n832), .A2(new_n833), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n839), .A2(new_n189), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n899), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n796), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n891), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n895), .A2(new_n901), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n907), .A2(new_n903), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT51), .A4(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n770), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n384), .B(new_n919), .C1(new_n894), .C2(new_n649), .ZN(new_n920));
  INV_X1    g734(.A(new_n784), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(KEYINPUT48), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(KEYINPUT48), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n915), .A2(new_n918), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n890), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(G952), .A2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n844), .B1(new_n927), .B2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n269), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(G210), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n932), .B(new_n299), .C1(new_n880), .C2(new_n888), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n349), .B1(new_n355), .B2(new_n356), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n318), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT55), .Z(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(KEYINPUT56), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n931), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n889), .A2(G902), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT117), .B1(new_n939), .B2(new_n932), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT117), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT56), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n944), .B2(new_n936), .ZN(G51));
  XNOR2_X1  g759(.A(new_n775), .B(KEYINPUT118), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT57), .Z(new_n947));
  AND3_X1   g761(.A1(new_n880), .A2(new_n888), .A3(new_n845), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n845), .B1(new_n880), .B2(new_n888), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n734), .ZN(new_n951));
  OR3_X1    g765(.A1(new_n939), .A2(new_n812), .A3(new_n815), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n930), .B1(new_n951), .B2(new_n952), .ZN(G54));
  INV_X1    g767(.A(new_n483), .ZN(new_n954));
  NAND2_X1  g768(.A1(KEYINPUT58), .A2(G475), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n939), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n931), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n939), .A2(new_n954), .A3(new_n955), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(G60));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT59), .ZN(new_n961));
  OAI221_X1 g775(.A(new_n961), .B1(new_n645), .B2(new_n643), .C1(new_n948), .C2(new_n949), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n931), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n890), .A2(new_n961), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n643), .A2(new_n645), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(G63));
  XNOR2_X1  g780(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n889), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n514), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT120), .B1(new_n973), .B2(new_n931), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n969), .B1(new_n880), .B2(new_n888), .ZN(new_n975));
  OAI211_X1 g789(.A(KEYINPUT120), .B(new_n931), .C1(new_n975), .C2(new_n514), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n682), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n967), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n973), .A2(KEYINPUT61), .A3(new_n931), .A4(new_n977), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(G66));
  NAND2_X1  g795(.A1(new_n887), .A2(new_n269), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT121), .ZN(new_n983));
  INV_X1    g797(.A(G224), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n390), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT122), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n934), .B1(G898), .B2(new_n269), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  XNOR2_X1  g803(.A(new_n575), .B(new_n477), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n849), .A2(new_n727), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n716), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n992), .A2(KEYINPUT62), .A3(new_n716), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n796), .B1(new_n806), .B2(KEYINPUT44), .ZN(new_n998));
  INV_X1    g812(.A(new_n810), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(new_n808), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n821), .A2(new_n822), .ZN(new_n1001));
  AOI21_X1  g815(.A(KEYINPUT107), .B1(new_n826), .B2(new_n699), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n795), .A2(new_n865), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n629), .A2(new_n310), .A3(new_n699), .A4(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT123), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n997), .A2(new_n1003), .A3(new_n834), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n991), .B1(new_n1007), .B2(new_n269), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT126), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1003), .A2(new_n1009), .A3(new_n992), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n921), .A2(new_n762), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(new_n823), .B2(new_n827), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n1014), .B(new_n1011), .C1(new_n823), .C2(new_n827), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1010), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n992), .ZN(new_n1017));
  OAI21_X1  g831(.A(KEYINPUT126), .B1(new_n828), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n834), .A2(new_n851), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n269), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(G900), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(G953), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT125), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1008), .B1(new_n1025), .B2(new_n991), .ZN(new_n1026));
  INV_X1    g840(.A(G227), .ZN(new_n1027));
  OAI21_X1  g841(.A(G953), .B1(new_n1027), .B2(new_n1022), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n990), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1007), .A2(new_n269), .ZN(new_n1030));
  AOI21_X1  g844(.A(KEYINPUT124), .B1(new_n1030), .B2(new_n990), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT124), .ZN(new_n1032));
  AOI211_X1 g846(.A(new_n1032), .B(new_n991), .C1(new_n1007), .C2(new_n269), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1028), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g848(.A1(new_n1026), .A2(new_n1028), .B1(new_n1029), .B2(new_n1034), .ZN(G72));
  NAND2_X1  g849(.A1(new_n711), .A2(new_n595), .ZN(new_n1036));
  OR3_X1    g850(.A1(new_n1016), .A2(new_n1020), .A3(new_n887), .ZN(new_n1037));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT63), .Z(new_n1039));
  AOI21_X1  g853(.A(new_n1036), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1039), .B1(new_n1007), .B2(new_n887), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n712), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1039), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1043), .B1(new_n623), .B2(new_n596), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n930), .B1(new_n889), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1040), .A2(new_n1046), .ZN(G57));
endmodule


