//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n205), .A2(KEYINPUT25), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT24), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n205), .A2(new_n208), .A3(new_n207), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n210), .B(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n214), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n216), .B1(new_n221), .B2(KEYINPUT25), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT26), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT65), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(new_n204), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n204), .A2(new_n223), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(KEYINPUT66), .A3(new_n211), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT28), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT27), .B(G183gat), .ZN(new_n234));
  INV_X1    g033(.A(G190gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  AND4_X1   g039(.A1(new_n233), .A2(new_n238), .A3(new_n240), .A4(new_n235), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n232), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT66), .B1(new_n231), .B2(new_n211), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n222), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n203), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n211), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n232), .A3(new_n242), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n202), .B1(new_n251), .B2(new_n222), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT73), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT73), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT29), .B1(new_n251), .B2(new_n222), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(new_n203), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(KEYINPUT22), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G211gat), .B(G218gat), .Z(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n203), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n255), .B2(new_n203), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n264), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  NAND4_X1  g072(.A1(new_n265), .A2(KEYINPUT30), .A3(new_n270), .A4(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n273), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n269), .B1(new_n253), .B2(new_n256), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n267), .A2(new_n264), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT74), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n245), .A2(new_n246), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT73), .B1(new_n280), .B2(new_n202), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(KEYINPUT73), .B2(new_n267), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n270), .B1(new_n282), .B2(new_n269), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT74), .B1(new_n283), .B2(new_n275), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT75), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n277), .B1(new_n257), .B2(new_n264), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(new_n273), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n274), .A4(new_n278), .ZN(new_n290));
  NAND2_X1  g089(.A1(G225gat), .A2(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n293), .B1(new_n296), .B2(KEYINPUT2), .ZN(new_n297));
  XOR2_X1   g096(.A(G141gat), .B(G148gat), .Z(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT77), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G141gat), .ZN(new_n304));
  INV_X1    g103(.A(G148gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n311), .A3(new_n307), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n296), .A2(new_n293), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  INV_X1    g115(.A(G120gat), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n317), .A2(G113gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(G113gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G127gat), .B(G134gat), .Z(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT67), .B(G120gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G113gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n321), .A2(KEYINPUT1), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n303), .A2(new_n315), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n301), .A3(new_n302), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n322), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n292), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n315), .A2(new_n335), .A3(new_n301), .A4(new_n302), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n332), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n303), .B2(new_n315), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n291), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n327), .A2(new_n316), .A3(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n341), .A2(new_n326), .B1(new_n320), .B2(new_n321), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n303), .A4(new_n315), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n331), .B2(new_n332), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n334), .B(KEYINPUT5), .C1(new_n339), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n344), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n342), .A2(new_n315), .A3(new_n303), .A4(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(new_n331), .B2(new_n332), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n336), .A2(new_n332), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n292), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT0), .ZN(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n357), .A3(new_n362), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n358), .A2(KEYINPUT6), .A3(new_n363), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n265), .A2(new_n270), .A3(new_n273), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n367), .A2(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n285), .A2(new_n290), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT69), .B(G71gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(G99gat), .ZN(new_n374));
  XOR2_X1   g173(.A(G15gat), .B(G43gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n245), .A2(new_n342), .ZN(new_n377));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n332), .B(new_n222), .C1(new_n243), .C2(new_n244), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n376), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(KEYINPUT32), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n381), .B(KEYINPUT32), .C1(new_n382), .C2(new_n376), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n379), .A2(KEYINPUT34), .ZN(new_n388));
  INV_X1    g187(.A(new_n380), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n332), .B1(new_n251), .B2(new_n222), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT72), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n380), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT72), .A3(new_n388), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT34), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n379), .B1(new_n394), .B2(KEYINPUT70), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT70), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n399), .A3(new_n380), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n396), .B1(new_n401), .B2(KEYINPUT71), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT70), .B1(new_n389), .B2(new_n390), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n378), .A3(new_n400), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n404), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n387), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n393), .A2(new_n395), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(KEYINPUT34), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT71), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n385), .A2(new_n386), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n401), .A2(KEYINPUT71), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n335), .B1(new_n264), .B2(KEYINPUT29), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n331), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n336), .A2(new_n246), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n264), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n418), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G22gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT31), .B(G50gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  MUX2_X1   g225(.A(G22gat), .B(new_n423), .S(new_n426), .Z(new_n427));
  AND2_X1   g226(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n421), .A2(new_n427), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n406), .A2(new_n413), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT35), .B1(new_n372), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n367), .A2(new_n368), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT35), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n369), .A2(new_n370), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n436), .A2(new_n288), .A3(new_n274), .A4(new_n278), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n274), .A2(new_n278), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n440), .A2(KEYINPUT81), .A3(new_n288), .A4(new_n436), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n433), .A2(new_n435), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n430), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n402), .A2(new_n387), .A3(new_n405), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n411), .B1(new_n410), .B2(new_n412), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n406), .A2(KEYINPUT36), .A3(new_n413), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n372), .A2(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT38), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT37), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n452), .B(new_n270), .C1(new_n282), .C2(new_n269), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n287), .A2(new_n455), .A3(new_n452), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n273), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n283), .A2(KEYINPUT37), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n451), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n257), .A2(new_n269), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n452), .B1(new_n268), .B2(new_n264), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT38), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n455), .B1(new_n287), .B2(new_n452), .ZN(new_n463));
  NOR4_X1   g262(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT83), .A4(KEYINPUT37), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n275), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n430), .B1(new_n459), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n330), .A2(new_n333), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n291), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT39), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(KEYINPUT82), .A3(KEYINPUT39), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n349), .A2(new_n351), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n337), .A2(new_n338), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n292), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n477), .A2(KEYINPUT39), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n362), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n478), .A2(KEYINPUT40), .A3(new_n362), .A4(new_n479), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n364), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n439), .B2(new_n441), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n450), .A2(KEYINPUT80), .B1(new_n468), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n372), .A2(new_n444), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n448), .A2(new_n449), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n487), .A2(KEYINPUT80), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n443), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G57gat), .B(G64gat), .Z(new_n491));
  NAND2_X1  g290(.A1(G71gat), .A2(G78gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT9), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(KEYINPUT94), .A3(new_n493), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR3_X1   g299(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n492), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n492), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n506));
  INV_X1    g305(.A(G71gat), .ZN(new_n507));
  INV_X1    g306(.A(G78gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n505), .B1(new_n509), .B2(new_n499), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT93), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n498), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n513));
  NOR2_X1   g312(.A1(G71gat), .A2(G78gat), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n513), .A2(new_n505), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT20), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(G1gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT16), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n522), .A2(G1gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G8gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n516), .B2(new_n517), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT97), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n521), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT96), .ZN(new_n533));
  XOR2_X1   g332(.A(G127gat), .B(G155gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G183gat), .B(G211gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n531), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NOR2_X1   g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n541), .B1(KEYINPUT8), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G99gat), .B(G106gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(new_n545), .A3(new_n543), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(KEYINPUT98), .A3(new_n548), .ZN(new_n549));
  AOI211_X1 g348(.A(KEYINPUT98), .B(new_n545), .C1(new_n540), .C2(new_n543), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G43gat), .B(G50gat), .Z(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G29gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT14), .B(G29gat), .Z(new_n558));
  OAI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(G36gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT85), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n553), .A2(new_n554), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n559), .B(new_n562), .C1(new_n555), .C2(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT41), .ZN(new_n567));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568));
  OAI22_X1  g367(.A1(new_n552), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT86), .B1(new_n566), .B2(KEYINPUT17), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n564), .A2(new_n571), .A3(new_n572), .A4(new_n565), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n549), .A2(new_n551), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n566), .B2(KEYINPUT17), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n569), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT99), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n577), .A2(new_n579), .ZN(new_n581));
  XOR2_X1   g380(.A(G134gat), .B(G162gat), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n568), .A2(new_n567), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OR3_X1    g384(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n580), .B2(new_n581), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n538), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G8gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n527), .B(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n566), .B2(KEYINPUT17), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n565), .A3(new_n564), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n593), .A2(KEYINPUT18), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(KEYINPUT88), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(new_n598), .A3(new_n565), .A4(new_n564), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n566), .A2(new_n528), .A3(KEYINPUT89), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT89), .B1(new_n566), .B2(new_n528), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n597), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT87), .B(KEYINPUT13), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n594), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT90), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n596), .A2(new_n605), .A3(KEYINPUT90), .ZN(new_n609));
  INV_X1    g408(.A(new_n595), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n574), .B2(new_n592), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n594), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT18), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G197gat), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT11), .B(G169gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n596), .A2(new_n605), .A3(new_n621), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n614), .A2(KEYINPUT91), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT18), .B1(new_n611), .B2(new_n594), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT91), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n513), .A2(new_n505), .A3(new_n514), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n502), .A2(new_n503), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n510), .A2(KEYINPUT93), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n513), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n575), .A2(new_n641), .A3(KEYINPUT10), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n547), .A2(KEYINPUT100), .A3(new_n548), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n544), .A2(new_n644), .A3(new_n546), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n643), .B(new_n645), .C1(new_n512), .C2(new_n515), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n552), .B2(new_n641), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n647), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n636), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n647), .A2(new_n648), .ZN(new_n659));
  INV_X1    g458(.A(new_n642), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n650), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n653), .A2(KEYINPUT101), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n636), .B1(new_n653), .B2(KEYINPUT101), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(KEYINPUT102), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n658), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n589), .A2(new_n632), .A3(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n490), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n434), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g473(.A1(new_n439), .A2(new_n441), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(new_n677), .B2(new_n590), .ZN(new_n680));
  MUX2_X1   g479(.A(new_n679), .B(new_n680), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g480(.A(G15gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n406), .A2(new_n413), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n672), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n488), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n672), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n687), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n444), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NOR3_X1   g490(.A1(new_n538), .A2(new_n632), .A3(new_n670), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n450), .B1(new_n468), .B2(new_n485), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n693), .A2(new_n694), .A3(new_n443), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n693), .B2(new_n443), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n588), .A2(KEYINPUT44), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  INV_X1    g499(.A(new_n588), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n490), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n692), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT106), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n705), .B(new_n692), .C1(new_n699), .C2(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n434), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n490), .A2(new_n701), .A3(new_n692), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n556), .A3(new_n434), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(G1328gat));
  INV_X1    g513(.A(new_n675), .ZN(new_n715));
  OAI21_X1  g514(.A(G36gat), .B1(new_n707), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(G36gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n710), .A2(new_n717), .A3(new_n675), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT46), .Z(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n683), .A2(G43gat), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n710), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n703), .A2(new_n488), .ZN(new_n724));
  AOI211_X1 g523(.A(new_n721), .B(new_n723), .C1(new_n724), .C2(G43gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n704), .A2(new_n686), .A3(new_n706), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n723), .B1(new_n729), .B2(G43gat), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n727), .A2(new_n728), .B1(KEYINPUT47), .B2(new_n730), .ZN(G1330gat));
  OAI21_X1  g530(.A(G50gat), .B1(new_n703), .B2(new_n430), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n430), .A2(G50gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n710), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n704), .A2(new_n444), .A3(new_n706), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n736), .A2(new_n737), .A3(G50gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n736), .B2(G50gat), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n710), .A2(new_n733), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n735), .B1(new_n741), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n632), .A2(new_n670), .ZN(new_n743));
  NOR4_X1   g542(.A1(new_n695), .A2(new_n696), .A3(new_n589), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n434), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n675), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  NAND3_X1  g549(.A1(new_n744), .A2(new_n507), .A3(new_n684), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n744), .A2(new_n686), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n507), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n444), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT109), .B(G78gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1335gat));
  AOI22_X1  g556(.A1(new_n656), .A2(new_n657), .B1(new_n667), .B2(new_n668), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n758), .A2(new_n708), .A3(G85gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n588), .B1(new_n693), .B2(new_n443), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n538), .A2(new_n631), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(KEYINPUT111), .A3(new_n768), .ZN(new_n769));
  OR3_X1    g568(.A1(new_n765), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n769), .A2(new_n770), .A3(KEYINPUT112), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT112), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n759), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n699), .A2(new_n702), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n774), .A2(new_n538), .A3(new_n743), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n434), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G85gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n777), .ZN(G1336gat));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n675), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n766), .A2(new_n768), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n715), .A2(G92gat), .A3(new_n758), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT52), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n782), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n787), .A3(new_n780), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1337gat));
  NOR3_X1   g588(.A1(new_n758), .A2(new_n683), .A3(G99gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n771), .B2(new_n772), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n686), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G99gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1338gat));
  NAND2_X1  g593(.A1(new_n775), .A2(new_n444), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n758), .A2(G106gat), .A3(new_n430), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n781), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n769), .A2(new_n770), .A3(new_n797), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n796), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1339gat));
  NOR3_X1   g603(.A1(new_n589), .A2(new_n631), .A3(new_n670), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n611), .A2(new_n594), .B1(new_n602), .B2(new_n604), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT115), .B1(new_n806), .B2(new_n619), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n619), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n630), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n667), .A2(new_n668), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n635), .B1(new_n652), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT113), .B1(new_n649), .B2(new_n651), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n516), .A2(new_n575), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT10), .B1(new_n819), .B2(new_n646), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  NOR4_X1   g620(.A1(new_n820), .A2(new_n642), .A3(new_n821), .A4(new_n650), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n662), .A2(KEYINPUT54), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n817), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n814), .B1(new_n661), .B2(new_n650), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n826), .B(KEYINPUT114), .C1(new_n818), .C2(new_n822), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n816), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n813), .B1(new_n828), .B2(KEYINPUT55), .ZN(new_n829));
  INV_X1    g628(.A(new_n827), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n659), .A2(new_n651), .A3(new_n660), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n821), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n649), .A2(KEYINPUT113), .A3(new_n651), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT114), .B1(new_n834), .B2(new_n826), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n815), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n812), .A2(new_n829), .A3(new_n701), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n811), .A2(new_n758), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n623), .A2(new_n630), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n829), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n842), .B2(new_n701), .ZN(new_n843));
  INV_X1    g642(.A(new_n538), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n805), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n444), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n846), .A2(new_n434), .A3(new_n684), .A4(new_n715), .ZN(new_n847));
  OAI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n632), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n847), .B(KEYINPUT116), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n632), .A2(G113gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  OAI21_X1  g650(.A(G120gat), .B1(new_n847), .B2(new_n758), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n670), .A2(new_n323), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT117), .Z(new_n854));
  OAI21_X1  g653(.A(new_n852), .B1(new_n849), .B2(new_n854), .ZN(G1341gat));
  NOR2_X1   g654(.A1(new_n847), .A2(new_n844), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(G127gat), .Z(G1342gat));
  NOR3_X1   g656(.A1(new_n708), .A2(new_n683), .A3(new_n588), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n846), .A2(new_n715), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(G134gat), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT56), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(G134gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n686), .A2(new_n430), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n434), .B(new_n715), .C1(new_n864), .C2(KEYINPUT119), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n865), .B(new_n845), .C1(KEYINPUT119), .C2(new_n864), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n304), .A3(new_n631), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n845), .A2(new_n871), .A3(new_n430), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n829), .A2(new_n631), .A3(new_n838), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n810), .A2(new_n807), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n670), .A2(new_n874), .A3(new_n630), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n701), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n839), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n844), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n805), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n430), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT118), .B1(new_n880), .B2(KEYINPUT57), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n882), .B(new_n871), .C1(new_n845), .C2(new_n430), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n872), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n686), .A2(new_n708), .A3(new_n675), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n884), .A2(new_n632), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(KEYINPUT122), .ZN(new_n888));
  OAI21_X1  g687(.A(G141gat), .B1(new_n887), .B2(KEYINPUT122), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n870), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n872), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n627), .B1(new_n606), .B2(new_n607), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n621), .B1(new_n892), .B2(new_n609), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n893), .A2(new_n894), .B1(new_n828), .B2(KEYINPUT55), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n669), .B1(new_n836), .B2(new_n837), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n875), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n588), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n538), .B1(new_n898), .B2(new_n839), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n444), .B1(new_n899), .B2(new_n805), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n882), .B1(new_n900), .B2(new_n871), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n880), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n631), .A3(new_n885), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n868), .B1(new_n904), .B2(G141gat), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n867), .B1(new_n887), .B2(new_n304), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT120), .B1(new_n909), .B2(KEYINPUT58), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n890), .B1(new_n908), .B2(new_n910), .ZN(G1344gat));
  NAND3_X1  g710(.A1(new_n866), .A2(new_n305), .A3(new_n670), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n884), .A2(new_n758), .A3(new_n886), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(KEYINPUT59), .A3(new_n305), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n829), .A2(new_n701), .A3(new_n838), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n811), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(new_n917), .B2(new_n916), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n538), .B1(new_n919), .B2(new_n898), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n444), .B1(new_n920), .B2(new_n805), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n871), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n891), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n670), .A3(new_n885), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n915), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n912), .B1(new_n914), .B2(new_n925), .ZN(G1345gat));
  NAND3_X1  g725(.A1(new_n866), .A2(new_n294), .A3(new_n538), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n884), .A2(new_n844), .A3(new_n886), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n294), .ZN(G1346gat));
  NAND3_X1  g728(.A1(new_n866), .A2(new_n295), .A3(new_n701), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n884), .A2(new_n588), .A3(new_n886), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n295), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n845), .A2(new_n434), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n715), .A2(new_n431), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n632), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n934), .B(KEYINPUT124), .Z(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n632), .A2(G169gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT125), .Z(G1348gat));
  OAI21_X1  g740(.A(G176gat), .B1(new_n935), .B2(new_n758), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n758), .A2(G176gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT126), .ZN(G1349gat));
  OAI21_X1  g744(.A(G183gat), .B1(new_n935), .B2(new_n844), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n538), .A2(new_n234), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n938), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n935), .B2(new_n588), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n701), .A2(new_n235), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n938), .B2(new_n952), .ZN(G1351gat));
  AND3_X1   g752(.A1(new_n933), .A2(new_n675), .A3(new_n864), .ZN(new_n954));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n631), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n488), .A2(new_n675), .A3(new_n708), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n956), .B1(new_n922), .B2(new_n891), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n631), .A2(G197gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1352gat));
  INV_X1    g758(.A(G204gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n954), .A2(new_n960), .A3(new_n670), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT62), .Z(new_n962));
  AND2_X1   g761(.A1(new_n957), .A2(new_n670), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n960), .ZN(G1353gat));
  NAND3_X1  g763(.A1(new_n954), .A2(new_n259), .A3(new_n538), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n259), .B1(new_n957), .B2(new_n538), .ZN(new_n966));
  NOR2_X1   g765(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n966), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n965), .B1(new_n969), .B2(new_n971), .ZN(G1354gat));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n260), .A3(new_n701), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n957), .A2(new_n701), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n974), .B2(new_n260), .ZN(G1355gat));
endmodule


