

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n589), .A2(n553), .ZN(n804) );
  AND2_X1 U550 ( .A1(n711), .A2(n526), .ZN(n713) );
  AND2_X1 U551 ( .A1(n704), .A2(n703), .ZN(n705) );
  OR2_X1 U552 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U553 ( .A1(n650), .A2(n649), .ZN(n652) );
  NOR2_X1 U554 ( .A1(n657), .A2(n656), .ZN(n660) );
  XNOR2_X1 U555 ( .A(n658), .B(KEYINPUT29), .ZN(n659) );
  NOR2_X1 U556 ( .A1(n534), .A2(G2104), .ZN(n535) );
  AND2_X2 U557 ( .A1(n528), .A2(G2104), .ZN(n893) );
  INV_X1 U558 ( .A(KEYINPUT33), .ZN(n706) );
  BUF_X1 U559 ( .A(n665), .Z(n676) );
  INV_X1 U560 ( .A(KEYINPUT102), .ZN(n658) );
  INV_X1 U561 ( .A(n722), .ZN(n703) );
  INV_X1 U562 ( .A(KEYINPUT107), .ZN(n712) );
  INV_X1 U563 ( .A(n927), .ZN(n714) );
  XNOR2_X1 U564 ( .A(KEYINPUT93), .B(n622), .ZN(n744) );
  XNOR2_X1 U565 ( .A(n530), .B(n529), .ZN(n532) );
  NOR2_X1 U566 ( .A1(n748), .A2(n521), .ZN(n759) );
  BUF_X1 U567 ( .A(n620), .Z(G164) );
  BUF_X1 U568 ( .A(n621), .Z(G160) );
  XOR2_X1 U569 ( .A(KEYINPUT15), .B(n619), .Z(n519) );
  XNOR2_X1 U570 ( .A(n632), .B(n631), .ZN(n520) );
  XNOR2_X2 U571 ( .A(n624), .B(n623), .ZN(n666) );
  AND2_X1 U572 ( .A1(n932), .A2(n770), .ZN(n521) );
  AND2_X1 U573 ( .A1(n759), .A2(n766), .ZN(n522) );
  AND2_X1 U574 ( .A1(G8), .A2(n692), .ZN(n523) );
  OR2_X1 U575 ( .A1(n722), .A2(n721), .ZN(n524) );
  AND2_X1 U576 ( .A1(n723), .A2(n524), .ZN(n525) );
  OR2_X1 U577 ( .A1(n722), .A2(n710), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n523), .A2(n693), .ZN(n527) );
  AND2_X1 U579 ( .A1(n638), .A2(n637), .ZN(n639) );
  AND2_X1 U580 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U581 ( .A1(n667), .A2(n666), .ZN(n668) );
  INV_X1 U582 ( .A(KEYINPUT101), .ZN(n651) );
  INV_X1 U583 ( .A(KEYINPUT103), .ZN(n695) );
  NAND2_X1 U584 ( .A1(n746), .A2(n744), .ZN(n624) );
  INV_X1 U585 ( .A(n666), .ZN(n665) );
  INV_X1 U586 ( .A(G2105), .ZN(n534) );
  XNOR2_X1 U587 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n529) );
  INV_X1 U588 ( .A(G651), .ZN(n553) );
  BUF_X1 U589 ( .A(n728), .Z(n898) );
  NOR2_X1 U590 ( .A1(G651), .A2(n589), .ZN(n808) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n803) );
  NOR2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n621) );
  XNOR2_X1 U593 ( .A(KEYINPUT71), .B(n569), .ZN(G171) );
  INV_X1 U594 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U595 ( .A1(G101), .A2(n893), .ZN(n530) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U597 ( .A1(G113), .A2(n897), .ZN(n531) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n540) );
  NOR2_X1 U599 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XOR2_X1 U600 ( .A(KEYINPUT17), .B(n533), .Z(n727) );
  NAND2_X1 U601 ( .A1(n727), .A2(G137), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n535), .B(KEYINPUT66), .ZN(n543) );
  INV_X1 U603 ( .A(n543), .ZN(n536) );
  INV_X1 U604 ( .A(n536), .ZN(n728) );
  NAND2_X1 U605 ( .A1(G125), .A2(n728), .ZN(n537) );
  NAND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U607 ( .A1(G102), .A2(n893), .ZN(n542) );
  NAND2_X1 U608 ( .A1(G138), .A2(n727), .ZN(n541) );
  NAND2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n543), .A2(G126), .ZN(n545) );
  NAND2_X1 U611 ( .A1(G114), .A2(n897), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n547) );
  INV_X1 U613 ( .A(KEYINPUT91), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT92), .ZN(n620) );
  NAND2_X1 U617 ( .A1(G91), .A2(n803), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT0), .B(G543), .Z(n589) );
  NAND2_X1 U619 ( .A1(G78), .A2(n804), .ZN(n551) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n808), .A2(G53), .ZN(n557) );
  NOR2_X1 U622 ( .A1(G543), .A2(n553), .ZN(n554) );
  XOR2_X1 U623 ( .A(KEYINPUT68), .B(n554), .Z(n555) );
  XNOR2_X2 U624 ( .A(KEYINPUT1), .B(n555), .ZN(n809) );
  NAND2_X1 U625 ( .A1(G65), .A2(n809), .ZN(n556) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n558) );
  OR2_X1 U627 ( .A1(n559), .A2(n558), .ZN(G299) );
  NAND2_X1 U628 ( .A1(n808), .A2(G52), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G64), .A2(n809), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(KEYINPUT69), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G90), .A2(n803), .ZN(n564) );
  NAND2_X1 U634 ( .A1(G77), .A2(n804), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U636 ( .A(n566), .B(n565), .ZN(n567) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n569) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G89), .A2(n803), .ZN(n570) );
  XOR2_X1 U640 ( .A(KEYINPUT4), .B(n570), .Z(n571) );
  XNOR2_X1 U641 ( .A(n571), .B(KEYINPUT79), .ZN(n573) );
  NAND2_X1 U642 ( .A1(G76), .A2(n804), .ZN(n572) );
  NAND2_X1 U643 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT5), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n808), .A2(G51), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G63), .A2(n809), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U648 ( .A(KEYINPUT6), .B(n577), .Z(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U651 ( .A1(n808), .A2(G50), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G62), .A2(n809), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U654 ( .A(KEYINPUT88), .B(n583), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G75), .A2(n804), .ZN(n584) );
  XNOR2_X1 U656 ( .A(KEYINPUT89), .B(n584), .ZN(n585) );
  NOR2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n803), .A2(G88), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(G303) );
  XOR2_X1 U660 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U661 ( .A1(G87), .A2(n589), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G49), .A2(n808), .ZN(n591) );
  NAND2_X1 U663 ( .A1(G74), .A2(G651), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U665 ( .A1(n809), .A2(n592), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT83), .B(n593), .Z(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n596), .B(KEYINPUT84), .ZN(G288) );
  NAND2_X1 U669 ( .A1(n804), .A2(G73), .ZN(n598) );
  XNOR2_X1 U670 ( .A(KEYINPUT2), .B(KEYINPUT86), .ZN(n597) );
  XNOR2_X1 U671 ( .A(n598), .B(n597), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G86), .A2(n803), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G48), .A2(n808), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G61), .A2(n809), .ZN(n601) );
  XNOR2_X1 U676 ( .A(KEYINPUT85), .B(n601), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U679 ( .A(KEYINPUT87), .B(n606), .Z(G305) );
  NAND2_X1 U680 ( .A1(G85), .A2(n803), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G60), .A2(n809), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G72), .A2(n804), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G47), .A2(n808), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  OR2_X1 U686 ( .A1(n612), .A2(n611), .ZN(G290) );
  NAND2_X1 U687 ( .A1(G92), .A2(n803), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G79), .A2(n804), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n808), .A2(G54), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G66), .A2(n809), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(KEYINPUT77), .B(n519), .ZN(n785) );
  NOR2_X2 U695 ( .A1(n620), .A2(G1384), .ZN(n746) );
  NAND2_X1 U696 ( .A1(G40), .A2(n621), .ZN(n622) );
  INV_X1 U697 ( .A(KEYINPUT64), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G2067), .A2(n666), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n665), .A2(G1348), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n643) );
  NOR2_X1 U701 ( .A1(n785), .A2(n643), .ZN(n642) );
  NAND2_X1 U702 ( .A1(n666), .A2(G1996), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(KEYINPUT26), .ZN(n640) );
  NAND2_X1 U704 ( .A1(n665), .A2(G1341), .ZN(n638) );
  NAND2_X1 U705 ( .A1(n803), .A2(G81), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT12), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G68), .A2(n804), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT13), .B(KEYINPUT76), .Z(n631) );
  NAND2_X1 U710 ( .A1(G56), .A2(n809), .ZN(n633) );
  XOR2_X1 U711 ( .A(KEYINPUT14), .B(n633), .Z(n634) );
  NOR2_X1 U712 ( .A1(n520), .A2(n634), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n808), .A2(G43), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n935) );
  INV_X1 U715 ( .A(n935), .ZN(n637) );
  NOR2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n645) );
  AND2_X1 U717 ( .A1(n785), .A2(n643), .ZN(n644) );
  NOR2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n650) );
  NAND2_X1 U719 ( .A1(G2072), .A2(n666), .ZN(n646) );
  XOR2_X1 U720 ( .A(KEYINPUT27), .B(n646), .Z(n648) );
  NAND2_X1 U721 ( .A1(n676), .A2(G1956), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n653) );
  NOR2_X1 U723 ( .A1(n653), .A2(G299), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n657) );
  NAND2_X1 U725 ( .A1(G299), .A2(n653), .ZN(n655) );
  XOR2_X1 U726 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n654) );
  XNOR2_X1 U727 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n660), .B(n659), .ZN(n664) );
  NOR2_X1 U729 ( .A1(G1961), .A2(n666), .ZN(n662) );
  XOR2_X1 U730 ( .A(G2078), .B(KEYINPUT25), .Z(n985) );
  NOR2_X1 U731 ( .A1(n676), .A2(n985), .ZN(n661) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n672) );
  NOR2_X1 U733 ( .A1(G301), .A2(n672), .ZN(n663) );
  NOR2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n690) );
  INV_X1 U735 ( .A(n690), .ZN(n683) );
  NAND2_X1 U736 ( .A1(n665), .A2(G8), .ZN(n722) );
  NOR2_X1 U737 ( .A1(G1966), .A2(n722), .ZN(n693) );
  INV_X1 U738 ( .A(G2084), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(KEYINPUT99), .ZN(n691) );
  NAND2_X1 U740 ( .A1(G8), .A2(n691), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n693), .A2(n669), .ZN(n670) );
  XOR2_X1 U742 ( .A(KEYINPUT30), .B(n670), .Z(n671) );
  NOR2_X1 U743 ( .A1(G168), .A2(n671), .ZN(n674) );
  AND2_X1 U744 ( .A1(G301), .A2(n672), .ZN(n673) );
  NOR2_X1 U745 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n675), .B(KEYINPUT31), .ZN(n689) );
  INV_X1 U747 ( .A(G8), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n676), .A2(G2090), .ZN(n678) );
  NOR2_X1 U749 ( .A1(G1971), .A2(n722), .ZN(n677) );
  NOR2_X1 U750 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n679), .A2(G303), .ZN(n680) );
  NOR2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n689), .A2(n685), .ZN(n682) );
  NAND2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n687) );
  AND2_X1 U755 ( .A1(G286), .A2(G8), .ZN(n684) );
  OR2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U758 ( .A(n688), .B(KEYINPUT32), .ZN(n698) );
  INV_X1 U759 ( .A(n691), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n694), .A2(n527), .ZN(n696) );
  XNOR2_X1 U761 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n716) );
  NOR2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n708) );
  NOR2_X1 U764 ( .A1(G1971), .A2(G303), .ZN(n699) );
  NOR2_X1 U765 ( .A1(n708), .A2(n699), .ZN(n941) );
  NAND2_X1 U766 ( .A1(n716), .A2(n941), .ZN(n701) );
  NAND2_X1 U767 ( .A1(G288), .A2(G1976), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n700), .B(KEYINPUT104), .ZN(n942) );
  NAND2_X1 U769 ( .A1(n701), .A2(n942), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(KEYINPUT105), .ZN(n704) );
  XNOR2_X1 U771 ( .A(n705), .B(KEYINPUT65), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U773 ( .A1(KEYINPUT33), .A2(n708), .ZN(n709) );
  XNOR2_X1 U774 ( .A(KEYINPUT106), .B(n709), .ZN(n710) );
  XNOR2_X1 U775 ( .A(n713), .B(n712), .ZN(n715) );
  XNOR2_X1 U776 ( .A(G1981), .B(G305), .ZN(n927) );
  NAND2_X1 U777 ( .A1(n715), .A2(n714), .ZN(n724) );
  NOR2_X1 U778 ( .A1(G2090), .A2(G303), .ZN(n717) );
  NAND2_X1 U779 ( .A1(G8), .A2(n717), .ZN(n718) );
  NAND2_X1 U780 ( .A1(n716), .A2(n718), .ZN(n719) );
  NAND2_X1 U781 ( .A1(n719), .A2(n722), .ZN(n723) );
  NOR2_X1 U782 ( .A1(G1981), .A2(G305), .ZN(n720) );
  XOR2_X1 U783 ( .A(n720), .B(KEYINPUT24), .Z(n721) );
  NAND2_X1 U784 ( .A1(n724), .A2(n525), .ZN(n760) );
  NAND2_X1 U785 ( .A1(G107), .A2(n897), .ZN(n726) );
  NAND2_X1 U786 ( .A1(G95), .A2(n893), .ZN(n725) );
  NAND2_X1 U787 ( .A1(n726), .A2(n725), .ZN(n732) );
  BUF_X1 U788 ( .A(n727), .Z(n894) );
  NAND2_X1 U789 ( .A1(n894), .A2(G131), .ZN(n730) );
  NAND2_X1 U790 ( .A1(G119), .A2(n898), .ZN(n729) );
  NAND2_X1 U791 ( .A1(n730), .A2(n729), .ZN(n731) );
  OR2_X1 U792 ( .A1(n732), .A2(n731), .ZN(n888) );
  NAND2_X1 U793 ( .A1(G1991), .A2(n888), .ZN(n743) );
  NAND2_X1 U794 ( .A1(G117), .A2(n897), .ZN(n734) );
  NAND2_X1 U795 ( .A1(G129), .A2(n898), .ZN(n733) );
  NAND2_X1 U796 ( .A1(n734), .A2(n733), .ZN(n737) );
  NAND2_X1 U797 ( .A1(n893), .A2(G105), .ZN(n735) );
  XOR2_X1 U798 ( .A(KEYINPUT38), .B(n735), .Z(n736) );
  NOR2_X1 U799 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U800 ( .A(KEYINPUT95), .B(n738), .Z(n740) );
  NAND2_X1 U801 ( .A1(n894), .A2(G141), .ZN(n739) );
  NAND2_X1 U802 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U803 ( .A(KEYINPUT96), .B(n741), .ZN(n908) );
  NAND2_X1 U804 ( .A1(G1996), .A2(n908), .ZN(n742) );
  NAND2_X1 U805 ( .A1(n743), .A2(n742), .ZN(n1024) );
  INV_X1 U806 ( .A(n744), .ZN(n745) );
  NOR2_X1 U807 ( .A1(n746), .A2(n745), .ZN(n770) );
  NAND2_X1 U808 ( .A1(n1024), .A2(n770), .ZN(n747) );
  XNOR2_X1 U809 ( .A(n747), .B(KEYINPUT97), .ZN(n763) );
  XNOR2_X1 U810 ( .A(KEYINPUT98), .B(n763), .ZN(n748) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n932) );
  NAND2_X1 U812 ( .A1(n893), .A2(G104), .ZN(n749) );
  XNOR2_X1 U813 ( .A(n749), .B(KEYINPUT94), .ZN(n751) );
  NAND2_X1 U814 ( .A1(G140), .A2(n894), .ZN(n750) );
  NAND2_X1 U815 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U816 ( .A(KEYINPUT34), .B(n752), .ZN(n757) );
  NAND2_X1 U817 ( .A1(G116), .A2(n897), .ZN(n754) );
  NAND2_X1 U818 ( .A1(G128), .A2(n898), .ZN(n753) );
  NAND2_X1 U819 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U820 ( .A(KEYINPUT35), .B(n755), .Z(n756) );
  NOR2_X1 U821 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U822 ( .A(KEYINPUT36), .B(n758), .ZN(n911) );
  XNOR2_X1 U823 ( .A(KEYINPUT37), .B(G2067), .ZN(n768) );
  NOR2_X1 U824 ( .A1(n911), .A2(n768), .ZN(n1009) );
  NAND2_X1 U825 ( .A1(n770), .A2(n1009), .ZN(n766) );
  NAND2_X1 U826 ( .A1(n760), .A2(n522), .ZN(n773) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n908), .ZN(n1013) );
  NOR2_X1 U828 ( .A1(G1986), .A2(G290), .ZN(n761) );
  NOR2_X1 U829 ( .A1(G1991), .A2(n888), .ZN(n1006) );
  NOR2_X1 U830 ( .A1(n761), .A2(n1006), .ZN(n762) );
  NOR2_X1 U831 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U832 ( .A1(n1013), .A2(n764), .ZN(n765) );
  XNOR2_X1 U833 ( .A(n765), .B(KEYINPUT39), .ZN(n767) );
  NAND2_X1 U834 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U835 ( .A1(n911), .A2(n768), .ZN(n1010) );
  NAND2_X1 U836 ( .A1(n769), .A2(n1010), .ZN(n771) );
  NAND2_X1 U837 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U838 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U839 ( .A(n774), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U841 ( .A(G57), .ZN(G237) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  XOR2_X1 U843 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n776) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U845 ( .A(n776), .B(n775), .ZN(G223) );
  XOR2_X1 U846 ( .A(G223), .B(KEYINPUT74), .Z(n839) );
  NAND2_X1 U847 ( .A1(n839), .A2(G567), .ZN(n777) );
  XNOR2_X1 U848 ( .A(n777), .B(KEYINPUT75), .ZN(n778) );
  XNOR2_X1 U849 ( .A(KEYINPUT11), .B(n778), .ZN(G234) );
  INV_X1 U850 ( .A(G860), .ZN(n784) );
  OR2_X1 U851 ( .A1(n935), .A2(n784), .ZN(G153) );
  NOR2_X1 U852 ( .A1(G868), .A2(n785), .ZN(n780) );
  INV_X1 U853 ( .A(G868), .ZN(n824) );
  NOR2_X1 U854 ( .A1(n824), .A2(G301), .ZN(n779) );
  NOR2_X1 U855 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U856 ( .A(KEYINPUT78), .B(n781), .ZN(G284) );
  NOR2_X1 U857 ( .A1(G286), .A2(n824), .ZN(n783) );
  NOR2_X1 U858 ( .A1(G868), .A2(G299), .ZN(n782) );
  NOR2_X1 U859 ( .A1(n783), .A2(n782), .ZN(G297) );
  NAND2_X1 U860 ( .A1(n784), .A2(G559), .ZN(n786) );
  INV_X1 U861 ( .A(n785), .ZN(n930) );
  NAND2_X1 U862 ( .A1(n786), .A2(n930), .ZN(n787) );
  XNOR2_X1 U863 ( .A(n787), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U864 ( .A1(n930), .A2(G868), .ZN(n788) );
  NOR2_X1 U865 ( .A1(G559), .A2(n788), .ZN(n789) );
  XNOR2_X1 U866 ( .A(n789), .B(KEYINPUT80), .ZN(n791) );
  NOR2_X1 U867 ( .A1(n935), .A2(G868), .ZN(n790) );
  NOR2_X1 U868 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U869 ( .A1(G111), .A2(n897), .ZN(n793) );
  NAND2_X1 U870 ( .A1(G99), .A2(n893), .ZN(n792) );
  NAND2_X1 U871 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U872 ( .A1(n898), .A2(G123), .ZN(n794) );
  XOR2_X1 U873 ( .A(KEYINPUT18), .B(n794), .Z(n795) );
  NOR2_X1 U874 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U875 ( .A1(n894), .A2(G135), .ZN(n797) );
  NAND2_X1 U876 ( .A1(n798), .A2(n797), .ZN(n1003) );
  XNOR2_X1 U877 ( .A(n1003), .B(G2096), .ZN(n799) );
  XNOR2_X1 U878 ( .A(n799), .B(KEYINPUT81), .ZN(n801) );
  INV_X1 U879 ( .A(G2100), .ZN(n800) );
  NAND2_X1 U880 ( .A1(n801), .A2(n800), .ZN(G156) );
  NAND2_X1 U881 ( .A1(G559), .A2(n930), .ZN(n802) );
  XNOR2_X1 U882 ( .A(n802), .B(n935), .ZN(n820) );
  NOR2_X1 U883 ( .A1(n820), .A2(G860), .ZN(n814) );
  NAND2_X1 U884 ( .A1(G93), .A2(n803), .ZN(n806) );
  NAND2_X1 U885 ( .A1(G80), .A2(n804), .ZN(n805) );
  NAND2_X1 U886 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U887 ( .A(KEYINPUT82), .B(n807), .ZN(n813) );
  NAND2_X1 U888 ( .A1(n808), .A2(G55), .ZN(n811) );
  NAND2_X1 U889 ( .A1(G67), .A2(n809), .ZN(n810) );
  NAND2_X1 U890 ( .A1(n811), .A2(n810), .ZN(n812) );
  OR2_X1 U891 ( .A1(n813), .A2(n812), .ZN(n823) );
  XOR2_X1 U892 ( .A(n814), .B(n823), .Z(G145) );
  INV_X1 U893 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U894 ( .A(G288), .B(KEYINPUT19), .ZN(n816) );
  XNOR2_X1 U895 ( .A(G290), .B(G166), .ZN(n815) );
  XNOR2_X1 U896 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U897 ( .A(n823), .B(n817), .ZN(n818) );
  XNOR2_X1 U898 ( .A(G299), .B(n818), .ZN(n819) );
  XNOR2_X1 U899 ( .A(n819), .B(G305), .ZN(n914) );
  XNOR2_X1 U900 ( .A(n914), .B(n820), .ZN(n821) );
  NAND2_X1 U901 ( .A1(n821), .A2(G868), .ZN(n822) );
  XNOR2_X1 U902 ( .A(n822), .B(KEYINPUT90), .ZN(n826) );
  NAND2_X1 U903 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U904 ( .A1(n826), .A2(n825), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2078), .A2(G2084), .ZN(n827) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n827), .Z(n828) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n828), .ZN(n829) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n829), .ZN(n830) );
  NAND2_X1 U909 ( .A1(n830), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U911 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NOR2_X1 U912 ( .A1(G219), .A2(G220), .ZN(n831) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n831), .Z(n832) );
  NOR2_X1 U914 ( .A1(G218), .A2(n832), .ZN(n833) );
  NAND2_X1 U915 ( .A1(G96), .A2(n833), .ZN(n843) );
  NAND2_X1 U916 ( .A1(n843), .A2(G2106), .ZN(n837) );
  NAND2_X1 U917 ( .A1(G69), .A2(G120), .ZN(n834) );
  NOR2_X1 U918 ( .A1(G237), .A2(n834), .ZN(n835) );
  NAND2_X1 U919 ( .A1(G108), .A2(n835), .ZN(n844) );
  NAND2_X1 U920 ( .A1(n844), .A2(G567), .ZN(n836) );
  NAND2_X1 U921 ( .A1(n837), .A2(n836), .ZN(n925) );
  NAND2_X1 U922 ( .A1(G483), .A2(G661), .ZN(n838) );
  NOR2_X1 U923 ( .A1(n925), .A2(n838), .ZN(n842) );
  NAND2_X1 U924 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U927 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U929 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U936 ( .A(G1348), .B(G2454), .ZN(n845) );
  XNOR2_X1 U937 ( .A(n845), .B(G2430), .ZN(n846) );
  XNOR2_X1 U938 ( .A(n846), .B(G1341), .ZN(n852) );
  XOR2_X1 U939 ( .A(G2443), .B(G2427), .Z(n848) );
  XNOR2_X1 U940 ( .A(G2438), .B(G2446), .ZN(n847) );
  XNOR2_X1 U941 ( .A(n848), .B(n847), .ZN(n850) );
  XOR2_X1 U942 ( .A(G2451), .B(G2435), .Z(n849) );
  XNOR2_X1 U943 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U944 ( .A(n852), .B(n851), .ZN(n853) );
  NAND2_X1 U945 ( .A1(n853), .A2(G14), .ZN(n854) );
  XOR2_X1 U946 ( .A(KEYINPUT108), .B(n854), .Z(G401) );
  XOR2_X1 U947 ( .A(G2100), .B(G2096), .Z(n856) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n855) );
  XNOR2_X1 U949 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2090), .Z(n858) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U952 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U953 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n861) );
  XNOR2_X1 U955 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U956 ( .A(G2474), .B(G1971), .Z(n864) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U958 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U959 ( .A(n865), .B(KEYINPUT109), .Z(n867) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1956), .ZN(n866) );
  XNOR2_X1 U961 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U962 ( .A(G1976), .B(G1981), .Z(n869) );
  XNOR2_X1 U963 ( .A(G1966), .B(G1961), .ZN(n868) );
  XNOR2_X1 U964 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U965 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n872) );
  XNOR2_X1 U967 ( .A(n873), .B(n872), .ZN(G229) );
  NAND2_X1 U968 ( .A1(G112), .A2(n897), .ZN(n875) );
  NAND2_X1 U969 ( .A1(G100), .A2(n893), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U971 ( .A1(G124), .A2(n898), .ZN(n876) );
  XNOR2_X1 U972 ( .A(n876), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G136), .A2(n894), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U975 ( .A1(n880), .A2(n879), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G118), .A2(n897), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G130), .A2(n898), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n887) );
  NAND2_X1 U979 ( .A1(G106), .A2(n893), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G142), .A2(n894), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U985 ( .A(KEYINPUT48), .B(n890), .ZN(n892) );
  XNOR2_X1 U986 ( .A(G164), .B(KEYINPUT46), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n907) );
  NAND2_X1 U988 ( .A1(G103), .A2(n893), .ZN(n896) );
  NAND2_X1 U989 ( .A1(G139), .A2(n894), .ZN(n895) );
  NAND2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n904) );
  NAND2_X1 U991 ( .A1(G115), .A2(n897), .ZN(n900) );
  NAND2_X1 U992 ( .A1(G127), .A2(n898), .ZN(n899) );
  NAND2_X1 U993 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(KEYINPUT111), .B(n901), .ZN(n902) );
  XNOR2_X1 U995 ( .A(KEYINPUT47), .B(n902), .ZN(n903) );
  NOR2_X1 U996 ( .A1(n904), .A2(n903), .ZN(n1018) );
  XOR2_X1 U997 ( .A(G162), .B(n1018), .Z(n905) );
  XNOR2_X1 U998 ( .A(n1003), .B(n905), .ZN(n906) );
  XOR2_X1 U999 ( .A(n907), .B(n906), .Z(n910) );
  XNOR2_X1 U1000 ( .A(G160), .B(n908), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n910), .B(n909), .ZN(n912) );
  XOR2_X1 U1002 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n913), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(n914), .B(KEYINPUT112), .ZN(n916) );
  XNOR2_X1 U1005 ( .A(n935), .B(n930), .ZN(n915) );
  XNOR2_X1 U1006 ( .A(n916), .B(n915), .ZN(n918) );
  XOR2_X1 U1007 ( .A(G286), .B(G171), .Z(n917) );
  XNOR2_X1 U1008 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n919), .ZN(G397) );
  OR2_X1 U1010 ( .A1(n925), .A2(G401), .ZN(n922) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n920) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1013 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n925), .ZN(G319) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1019 ( .A(G16), .B(KEYINPUT56), .ZN(n951) );
  XOR2_X1 U1020 ( .A(G168), .B(G1966), .Z(n926) );
  NOR2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1022 ( .A(KEYINPUT57), .B(n928), .Z(n949) );
  XNOR2_X1 U1023 ( .A(G1961), .B(G171), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(n929), .B(KEYINPUT118), .ZN(n940) );
  XNOR2_X1 U1025 ( .A(n930), .B(G1348), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(G1956), .B(G299), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n938) );
  XNOR2_X1 U1029 ( .A(G1341), .B(n935), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(KEYINPUT120), .B(n936), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n947) );
  AND2_X1 U1033 ( .A1(G303), .A2(G1971), .ZN(n944) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(KEYINPUT119), .B(n945), .ZN(n946) );
  NOR2_X1 U1037 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1038 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1039 ( .A1(n951), .A2(n950), .ZN(n980) );
  INV_X1 U1040 ( .A(G16), .ZN(n978) );
  XNOR2_X1 U1041 ( .A(G1986), .B(G24), .ZN(n956) );
  XNOR2_X1 U1042 ( .A(G1971), .B(G22), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G23), .B(G1976), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(KEYINPUT125), .B(n954), .ZN(n955) );
  NOR2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(KEYINPUT58), .B(n957), .ZN(n972) );
  XNOR2_X1 U1048 ( .A(KEYINPUT121), .B(G1981), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(n958), .B(G6), .ZN(n965) );
  XOR2_X1 U1050 ( .A(KEYINPUT123), .B(G4), .Z(n960) );
  XNOR2_X1 U1051 ( .A(G1348), .B(KEYINPUT59), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n960), .B(n959), .ZN(n961) );
  XOR2_X1 U1053 ( .A(KEYINPUT122), .B(n961), .Z(n963) );
  XNOR2_X1 U1054 ( .A(G1341), .B(G19), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(G20), .B(G1956), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1059 ( .A(KEYINPUT60), .B(n968), .Z(n970) );
  XNOR2_X1 U1060 ( .A(G1961), .B(G5), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1063 ( .A(KEYINPUT124), .B(G1966), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G21), .B(n973), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(KEYINPUT61), .B(n976), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1069 ( .A(KEYINPUT126), .B(n981), .Z(n1002) );
  XOR2_X1 U1070 ( .A(G1991), .B(G25), .Z(n982) );
  NAND2_X1 U1071 ( .A1(n982), .A2(G28), .ZN(n991) );
  XNOR2_X1 U1072 ( .A(G1996), .B(G32), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G33), .B(G2072), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n989) );
  XNOR2_X1 U1075 ( .A(G2067), .B(G26), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G27), .B(n985), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1080 ( .A(KEYINPUT53), .B(n992), .Z(n995) );
  XOR2_X1 U1081 ( .A(KEYINPUT54), .B(G34), .Z(n993) );
  XNOR2_X1 U1082 ( .A(G2084), .B(n993), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(G35), .B(G2090), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1086 ( .A(KEYINPUT55), .B(n998), .Z(n999) );
  NOR2_X1 U1087 ( .A1(G29), .A2(n999), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(KEYINPUT117), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1034) );
  INV_X1 U1090 ( .A(KEYINPUT55), .ZN(n1030) );
  XNOR2_X1 U1091 ( .A(G160), .B(G2084), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(KEYINPUT113), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(KEYINPUT114), .B(n1014), .Z(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT51), .B(n1015), .Z(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1026) );
  XNOR2_X1 U1102 ( .A(G2072), .B(n1018), .ZN(n1021) );
  XOR2_X1 U1103 ( .A(G2078), .B(KEYINPUT115), .Z(n1019) );
  XNOR2_X1 U1104 ( .A(G164), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(n1022), .B(KEYINPUT50), .ZN(n1023) );
  NOR2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(KEYINPUT116), .B(n1027), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(KEYINPUT52), .B(n1028), .Z(n1029) );
  NAND2_X1 U1111 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1112 ( .A1(n1031), .A2(G29), .ZN(n1032) );
  NAND2_X1 U1113 ( .A1(n1032), .A2(G11), .ZN(n1033) );
  NOR2_X1 U1114 ( .A1(n1034), .A2(n1033), .ZN(n1036) );
  XOR2_X1 U1115 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n1035) );
  XNOR2_X1 U1116 ( .A(n1036), .B(n1035), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

