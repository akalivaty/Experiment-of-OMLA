

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U558 ( .A1(n543), .A2(G2104), .ZN(n871) );
  OR2_X2 U559 ( .A1(n824), .A2(n823), .ZN(n825) );
  BUF_X1 U560 ( .A(n742), .Z(n699) );
  XNOR2_X1 U561 ( .A(KEYINPUT93), .B(n742), .ZN(n735) );
  NOR2_X2 U562 ( .A1(G2104), .A2(n543), .ZN(n874) );
  NOR2_X1 U563 ( .A1(n716), .A2(n715), .ZN(n710) );
  OR2_X1 U564 ( .A1(n729), .A2(G299), .ZN(n726) );
  XNOR2_X1 U565 ( .A(n589), .B(KEYINPUT13), .ZN(n522) );
  AND2_X1 U566 ( .A1(G1976), .A2(G288), .ZN(n523) );
  NOR2_X1 U567 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U568 ( .A1(n732), .A2(n731), .ZN(n734) );
  INV_X1 U569 ( .A(KEYINPUT103), .ZN(n759) );
  NOR2_X1 U570 ( .A1(n775), .A2(n523), .ZN(n776) );
  AND2_X1 U571 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U572 ( .A1(G164), .A2(G1384), .ZN(n782) );
  INV_X1 U573 ( .A(KEYINPUT17), .ZN(n538) );
  NAND2_X1 U574 ( .A1(n870), .A2(G138), .ZN(n540) );
  NOR2_X1 U575 ( .A1(G651), .A2(n654), .ZN(n662) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n654) );
  NAND2_X1 U577 ( .A1(G51), .A2(n662), .ZN(n526) );
  INV_X1 U578 ( .A(G651), .ZN(n529) );
  NOR2_X1 U579 ( .A1(G543), .A2(n529), .ZN(n524) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n524), .Z(n663) );
  NAND2_X1 U581 ( .A1(G63), .A2(n663), .ZN(n525) );
  NAND2_X1 U582 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(n527), .ZN(n536) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n657) );
  NAND2_X1 U585 ( .A1(n657), .A2(G89), .ZN(n528) );
  XNOR2_X1 U586 ( .A(n528), .B(KEYINPUT4), .ZN(n532) );
  OR2_X1 U587 ( .A1(n529), .A2(n654), .ZN(n530) );
  XNOR2_X2 U588 ( .A(KEYINPUT65), .B(n530), .ZN(n658) );
  NAND2_X1 U589 ( .A1(G76), .A2(n658), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U591 ( .A(KEYINPUT5), .B(n533), .ZN(n534) );
  XNOR2_X1 U592 ( .A(KEYINPUT73), .B(n534), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U594 ( .A(KEYINPUT7), .B(n537), .Z(G168) );
  XOR2_X1 U595 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  XNOR2_X2 U597 ( .A(n539), .B(n538), .ZN(n870) );
  XNOR2_X1 U598 ( .A(n540), .B(KEYINPUT88), .ZN(n542) );
  INV_X1 U599 ( .A(G2105), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n871), .A2(G102), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n874), .A2(G126), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G2105), .A2(G2104), .ZN(n544) );
  XOR2_X1 U604 ( .A(KEYINPUT64), .B(n544), .Z(n559) );
  BUF_X1 U605 ( .A(n559), .Z(n875) );
  NAND2_X1 U606 ( .A1(G114), .A2(n875), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X2 U608 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U609 ( .A1(G91), .A2(n657), .ZN(n550) );
  NAND2_X1 U610 ( .A1(G78), .A2(n658), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G53), .A2(n662), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G65), .A2(n663), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT68), .B(n555), .Z(G299) );
  NAND2_X1 U617 ( .A1(n870), .A2(G137), .ZN(n558) );
  NAND2_X1 U618 ( .A1(G101), .A2(n871), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT23), .B(n556), .Z(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n874), .A2(G125), .ZN(n561) );
  NAND2_X1 U622 ( .A1(G113), .A2(n559), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X2 U624 ( .A1(n563), .A2(n562), .ZN(G160) );
  XNOR2_X1 U625 ( .A(G2435), .B(G2443), .ZN(n573) );
  XOR2_X1 U626 ( .A(G2454), .B(G2430), .Z(n565) );
  XNOR2_X1 U627 ( .A(G2446), .B(KEYINPUT109), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n565), .B(n564), .ZN(n569) );
  XOR2_X1 U629 ( .A(G2451), .B(G2427), .Z(n567) );
  XNOR2_X1 U630 ( .A(G1348), .B(G1341), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U632 ( .A(n569), .B(n568), .Z(n571) );
  XNOR2_X1 U633 ( .A(KEYINPUT108), .B(G2438), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n573), .B(n572), .ZN(n574) );
  AND2_X1 U636 ( .A1(n574), .A2(G14), .ZN(G401) );
  NAND2_X1 U637 ( .A1(G52), .A2(n662), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G64), .A2(n663), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G90), .A2(n657), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G77), .A2(n658), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n579), .Z(n580) );
  NOR2_X1 U644 ( .A1(n581), .A2(n580), .ZN(G171) );
  INV_X1 U645 ( .A(G57), .ZN(G237) );
  INV_X1 U646 ( .A(G82), .ZN(G220) );
  NAND2_X1 U647 ( .A1(G94), .A2(G452), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U649 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(KEYINPUT10), .ZN(n584) );
  XNOR2_X1 U651 ( .A(KEYINPUT70), .B(n584), .ZN(G223) );
  INV_X1 U652 ( .A(G223), .ZN(n845) );
  NAND2_X1 U653 ( .A1(n845), .A2(G567), .ZN(n585) );
  XOR2_X1 U654 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U655 ( .A1(n657), .A2(G81), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G68), .A2(n658), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G43), .A2(n662), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n522), .A2(n590), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n663), .A2(G56), .ZN(n591) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(n591), .Z(n592) );
  NOR2_X2 U663 ( .A1(n593), .A2(n592), .ZN(n977) );
  NAND2_X1 U664 ( .A1(n977), .A2(G860), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G66), .A2(n663), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G92), .A2(n657), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G54), .A2(n662), .ZN(n597) );
  NAND2_X1 U670 ( .A1(G79), .A2(n658), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U672 ( .A(KEYINPUT71), .B(n598), .Z(n599) );
  NOR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT15), .B(n601), .ZN(n716) );
  INV_X1 U675 ( .A(G868), .ZN(n613) );
  NAND2_X1 U676 ( .A1(n716), .A2(n613), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT72), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(G284) );
  NOR2_X1 U680 ( .A1(G286), .A2(n613), .ZN(n606) );
  NOR2_X1 U681 ( .A1(G299), .A2(G868), .ZN(n605) );
  NOR2_X1 U682 ( .A1(n606), .A2(n605), .ZN(G297) );
  INV_X1 U683 ( .A(G860), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G559), .A2(n607), .ZN(n608) );
  XNOR2_X1 U685 ( .A(KEYINPUT74), .B(n608), .ZN(n609) );
  INV_X1 U686 ( .A(n716), .ZN(n632) );
  NAND2_X1 U687 ( .A1(n609), .A2(n632), .ZN(n610) );
  XNOR2_X1 U688 ( .A(KEYINPUT16), .B(n610), .ZN(G148) );
  NOR2_X1 U689 ( .A1(n716), .A2(n613), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n611), .B(KEYINPUT75), .ZN(n612) );
  NOR2_X1 U691 ( .A1(G559), .A2(n612), .ZN(n615) );
  AND2_X1 U692 ( .A1(n613), .A2(n977), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U694 ( .A1(G123), .A2(n874), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT18), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n617), .B(KEYINPUT76), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G99), .A2(n871), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G135), .A2(n870), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G111), .A2(n875), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n935) );
  XOR2_X1 U703 ( .A(G2096), .B(n935), .Z(n624) );
  NOR2_X1 U704 ( .A1(G2100), .A2(n624), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT77), .B(n625), .ZN(G156) );
  NAND2_X1 U706 ( .A1(G93), .A2(n657), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G80), .A2(n658), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G55), .A2(n662), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G67), .A2(n663), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n680) );
  NAND2_X1 U713 ( .A1(n632), .A2(G559), .ZN(n669) );
  XOR2_X1 U714 ( .A(n977), .B(n669), .Z(n633) );
  NOR2_X1 U715 ( .A1(G860), .A2(n633), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n680), .B(n634), .ZN(G145) );
  NAND2_X1 U717 ( .A1(G47), .A2(n662), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G60), .A2(n663), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U720 ( .A(KEYINPUT66), .B(n637), .Z(n641) );
  NAND2_X1 U721 ( .A1(G85), .A2(n657), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G72), .A2(n658), .ZN(n638) );
  AND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U725 ( .A1(G86), .A2(n657), .ZN(n642) );
  XOR2_X1 U726 ( .A(KEYINPUT78), .B(n642), .Z(n645) );
  NAND2_X1 U727 ( .A1(n658), .A2(G73), .ZN(n643) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n663), .A2(G61), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U732 ( .A(n648), .B(KEYINPUT79), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G48), .A2(n662), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(G305) );
  NAND2_X1 U735 ( .A1(G49), .A2(n662), .ZN(n652) );
  NAND2_X1 U736 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U738 ( .A1(n663), .A2(n653), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n654), .A2(G87), .ZN(n655) );
  NAND2_X1 U740 ( .A1(n656), .A2(n655), .ZN(G288) );
  NAND2_X1 U741 ( .A1(G88), .A2(n657), .ZN(n660) );
  NAND2_X1 U742 ( .A1(G75), .A2(n658), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U744 ( .A(KEYINPUT81), .B(n661), .ZN(n668) );
  NAND2_X1 U745 ( .A1(G50), .A2(n662), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G62), .A2(n663), .ZN(n664) );
  NAND2_X1 U747 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U748 ( .A(KEYINPUT80), .B(n666), .Z(n667) );
  NAND2_X1 U749 ( .A1(n668), .A2(n667), .ZN(G303) );
  INV_X1 U750 ( .A(G303), .ZN(G166) );
  XOR2_X1 U751 ( .A(KEYINPUT84), .B(n669), .Z(n678) );
  XNOR2_X1 U752 ( .A(G299), .B(G290), .ZN(n670) );
  XNOR2_X1 U753 ( .A(n670), .B(G305), .ZN(n674) );
  XNOR2_X1 U754 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n672) );
  XNOR2_X1 U755 ( .A(G288), .B(KEYINPUT82), .ZN(n671) );
  XNOR2_X1 U756 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U757 ( .A(n674), .B(n673), .Z(n676) );
  XNOR2_X1 U758 ( .A(G166), .B(n680), .ZN(n675) );
  XNOR2_X1 U759 ( .A(n676), .B(n675), .ZN(n677) );
  XOR2_X1 U760 ( .A(n977), .B(n677), .Z(n894) );
  XNOR2_X1 U761 ( .A(n678), .B(n894), .ZN(n679) );
  NAND2_X1 U762 ( .A1(n679), .A2(G868), .ZN(n682) );
  OR2_X1 U763 ( .A1(G868), .A2(n680), .ZN(n681) );
  NAND2_X1 U764 ( .A1(n682), .A2(n681), .ZN(G295) );
  NAND2_X1 U765 ( .A1(G2078), .A2(G2084), .ZN(n683) );
  XOR2_X1 U766 ( .A(KEYINPUT20), .B(n683), .Z(n684) );
  NAND2_X1 U767 ( .A1(G2090), .A2(n684), .ZN(n685) );
  XNOR2_X1 U768 ( .A(KEYINPUT21), .B(n685), .ZN(n686) );
  NAND2_X1 U769 ( .A1(n686), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U770 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U771 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n687) );
  XOR2_X1 U773 ( .A(KEYINPUT22), .B(n687), .Z(n688) );
  NOR2_X1 U774 ( .A1(G218), .A2(n688), .ZN(n689) );
  XOR2_X1 U775 ( .A(KEYINPUT85), .B(n689), .Z(n690) );
  NAND2_X1 U776 ( .A1(G96), .A2(n690), .ZN(n851) );
  NAND2_X1 U777 ( .A1(n851), .A2(G2106), .ZN(n696) );
  NAND2_X1 U778 ( .A1(G120), .A2(G69), .ZN(n691) );
  NOR2_X1 U779 ( .A1(G237), .A2(n691), .ZN(n692) );
  XNOR2_X1 U780 ( .A(KEYINPUT86), .B(n692), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n693), .A2(G108), .ZN(n850) );
  NAND2_X1 U782 ( .A1(G567), .A2(n850), .ZN(n694) );
  XOR2_X1 U783 ( .A(KEYINPUT87), .B(n694), .Z(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n852) );
  NAND2_X1 U785 ( .A1(G483), .A2(G661), .ZN(n697) );
  NOR2_X1 U786 ( .A1(n852), .A2(n697), .ZN(n849) );
  NAND2_X1 U787 ( .A1(n849), .A2(G36), .ZN(G176) );
  NAND2_X1 U788 ( .A1(G40), .A2(G160), .ZN(n781) );
  XNOR2_X1 U789 ( .A(n781), .B(KEYINPUT89), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n782), .A2(n698), .ZN(n742) );
  NAND2_X1 U791 ( .A1(G8), .A2(n699), .ZN(n819) );
  INV_X1 U792 ( .A(KEYINPUT104), .ZN(n774) );
  NOR2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n773) );
  NAND2_X1 U794 ( .A1(n774), .A2(n773), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n773), .A2(KEYINPUT33), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n700), .A2(KEYINPUT104), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n819), .A2(n703), .ZN(n780) );
  XOR2_X1 U799 ( .A(G1996), .B(KEYINPUT96), .Z(n959) );
  NOR2_X1 U800 ( .A1(n959), .A2(n742), .ZN(n704) );
  XNOR2_X1 U801 ( .A(n704), .B(KEYINPUT26), .ZN(n707) );
  NAND2_X1 U802 ( .A1(G1341), .A2(n742), .ZN(n705) );
  XNOR2_X1 U803 ( .A(n705), .B(KEYINPUT97), .ZN(n706) );
  NAND2_X1 U804 ( .A1(n708), .A2(n977), .ZN(n715) );
  INV_X1 U805 ( .A(KEYINPUT98), .ZN(n709) );
  XNOR2_X1 U806 ( .A(n710), .B(n709), .ZN(n714) );
  NAND2_X1 U807 ( .A1(G1348), .A2(n699), .ZN(n712) );
  NAND2_X1 U808 ( .A1(G2067), .A2(n735), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n727) );
  INV_X1 U813 ( .A(n735), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n719), .A2(G1956), .ZN(n723) );
  NAND2_X1 U815 ( .A1(n735), .A2(G2072), .ZN(n721) );
  INV_X1 U816 ( .A(KEYINPUT27), .ZN(n720) );
  XNOR2_X1 U817 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U818 ( .A1(n723), .A2(n722), .ZN(n725) );
  INV_X1 U819 ( .A(KEYINPUT95), .ZN(n724) );
  XNOR2_X1 U820 ( .A(n725), .B(n724), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U822 ( .A(KEYINPUT99), .B(n728), .ZN(n732) );
  NAND2_X1 U823 ( .A1(G299), .A2(n729), .ZN(n730) );
  XOR2_X1 U824 ( .A(n730), .B(KEYINPUT28), .Z(n731) );
  XNOR2_X1 U825 ( .A(KEYINPUT29), .B(KEYINPUT100), .ZN(n733) );
  XNOR2_X1 U826 ( .A(n734), .B(n733), .ZN(n740) );
  XNOR2_X1 U827 ( .A(G2078), .B(KEYINPUT25), .ZN(n950) );
  NAND2_X1 U828 ( .A1(n735), .A2(n950), .ZN(n736) );
  XNOR2_X1 U829 ( .A(n736), .B(KEYINPUT94), .ZN(n738) );
  INV_X1 U830 ( .A(G1961), .ZN(n1016) );
  NAND2_X1 U831 ( .A1(n1016), .A2(n699), .ZN(n737) );
  NAND2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U833 ( .A1(G171), .A2(n741), .ZN(n739) );
  NAND2_X1 U834 ( .A1(n740), .A2(n739), .ZN(n752) );
  NOR2_X1 U835 ( .A1(G171), .A2(n741), .ZN(n748) );
  NOR2_X1 U836 ( .A1(G1966), .A2(n819), .ZN(n767) );
  NOR2_X1 U837 ( .A1(G2084), .A2(n742), .ZN(n743) );
  XOR2_X1 U838 ( .A(KEYINPUT92), .B(n743), .Z(n763) );
  NAND2_X1 U839 ( .A1(G8), .A2(n763), .ZN(n744) );
  NOR2_X1 U840 ( .A1(n767), .A2(n744), .ZN(n745) );
  XOR2_X1 U841 ( .A(KEYINPUT30), .B(n745), .Z(n746) );
  NOR2_X1 U842 ( .A1(G168), .A2(n746), .ZN(n747) );
  NOR2_X1 U843 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U844 ( .A(n749), .B(KEYINPUT31), .ZN(n750) );
  XNOR2_X1 U845 ( .A(n750), .B(KEYINPUT101), .ZN(n751) );
  NAND2_X1 U846 ( .A1(n752), .A2(n751), .ZN(n765) );
  NAND2_X1 U847 ( .A1(n765), .A2(G286), .ZN(n758) );
  NOR2_X1 U848 ( .A1(G1971), .A2(n819), .ZN(n753) );
  XNOR2_X1 U849 ( .A(n753), .B(KEYINPUT102), .ZN(n755) );
  NOR2_X1 U850 ( .A1(n699), .A2(G2090), .ZN(n754) );
  NOR2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U852 ( .A1(n756), .A2(G303), .ZN(n757) );
  NAND2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U854 ( .A(n760), .B(n759), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n761), .A2(G8), .ZN(n762) );
  XNOR2_X1 U856 ( .A(n762), .B(KEYINPUT32), .ZN(n771) );
  INV_X1 U857 ( .A(n763), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n764), .A2(G8), .ZN(n769) );
  INV_X1 U859 ( .A(n765), .ZN(n766) );
  NOR2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n817) );
  NOR2_X1 U863 ( .A1(G1971), .A2(G303), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n983) );
  NAND2_X1 U865 ( .A1(n817), .A2(n983), .ZN(n777) );
  OR2_X1 U866 ( .A1(n819), .A2(n774), .ZN(n775) );
  NOR2_X1 U867 ( .A1(KEYINPUT33), .A2(n778), .ZN(n779) );
  NOR2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n811) );
  XOR2_X1 U869 ( .A(G1981), .B(G305), .Z(n974) );
  XOR2_X1 U870 ( .A(n781), .B(KEYINPUT89), .Z(n783) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n839) );
  XNOR2_X1 U872 ( .A(G2067), .B(KEYINPUT37), .ZN(n837) );
  NAND2_X1 U873 ( .A1(G140), .A2(n870), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G104), .A2(n871), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n786), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n874), .A2(G128), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G116), .A2(n875), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U880 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U882 ( .A(KEYINPUT36), .B(n792), .ZN(n889) );
  NOR2_X1 U883 ( .A1(n837), .A2(n889), .ZN(n944) );
  NAND2_X1 U884 ( .A1(n839), .A2(n944), .ZN(n835) );
  XOR2_X1 U885 ( .A(KEYINPUT90), .B(G1991), .Z(n949) );
  NAND2_X1 U886 ( .A1(G131), .A2(n870), .ZN(n794) );
  NAND2_X1 U887 ( .A1(G95), .A2(n871), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n874), .A2(G119), .ZN(n796) );
  NAND2_X1 U890 ( .A1(G107), .A2(n875), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n868) );
  NOR2_X1 U893 ( .A1(n949), .A2(n868), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G141), .A2(n870), .ZN(n800) );
  NAND2_X1 U895 ( .A1(G129), .A2(n874), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n871), .A2(G105), .ZN(n801) );
  XOR2_X1 U898 ( .A(KEYINPUT38), .B(n801), .Z(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U900 ( .A1(G117), .A2(n875), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n869) );
  AND2_X1 U902 ( .A1(G1996), .A2(n869), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n938) );
  XNOR2_X1 U904 ( .A(KEYINPUT91), .B(n839), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n938), .A2(n808), .ZN(n831) );
  INV_X1 U906 ( .A(n831), .ZN(n809) );
  AND2_X1 U907 ( .A1(n835), .A2(n809), .ZN(n812) );
  AND2_X1 U908 ( .A1(n974), .A2(n812), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n826) );
  INV_X1 U910 ( .A(n812), .ZN(n824) );
  NOR2_X1 U911 ( .A1(G1981), .A2(G305), .ZN(n813) );
  XOR2_X1 U912 ( .A(n813), .B(KEYINPUT24), .Z(n814) );
  OR2_X1 U913 ( .A1(n819), .A2(n814), .ZN(n822) );
  NOR2_X1 U914 ( .A1(G2090), .A2(G303), .ZN(n815) );
  XOR2_X1 U915 ( .A(KEYINPUT105), .B(n815), .Z(n816) );
  NAND2_X1 U916 ( .A1(G8), .A2(n816), .ZN(n818) );
  NAND2_X1 U917 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n828) );
  XNOR2_X1 U921 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U922 ( .A1(n981), .A2(n839), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n842) );
  NOR2_X1 U924 ( .A1(G1996), .A2(n869), .ZN(n930) );
  AND2_X1 U925 ( .A1(n949), .A2(n868), .ZN(n936) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n829) );
  XNOR2_X1 U927 ( .A(KEYINPUT106), .B(n829), .ZN(n830) );
  NOR2_X1 U928 ( .A1(n936), .A2(n830), .ZN(n832) );
  NOR2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U930 ( .A1(n930), .A2(n833), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT39), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n837), .A2(n889), .ZN(n927) );
  NAND2_X1 U934 ( .A1(n838), .A2(n927), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(n844) );
  XOR2_X1 U937 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n843) );
  XNOR2_X1 U938 ( .A(n844), .B(n843), .ZN(G329) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n845), .ZN(G217) );
  NAND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n846) );
  XOR2_X1 U941 ( .A(KEYINPUT110), .B(n846), .Z(n847) );
  NAND2_X1 U942 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U944 ( .A1(n849), .A2(n848), .ZN(G188) );
  XNOR2_X1 U945 ( .A(G96), .B(KEYINPUT111), .ZN(G221) );
  INV_X1 U947 ( .A(G120), .ZN(G236) );
  INV_X1 U948 ( .A(G108), .ZN(G238) );
  INV_X1 U949 ( .A(G69), .ZN(G235) );
  NOR2_X1 U950 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U951 ( .A(G325), .ZN(G261) );
  INV_X1 U952 ( .A(n852), .ZN(G319) );
  NAND2_X1 U953 ( .A1(G124), .A2(n874), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G136), .A2(n870), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n854), .B(KEYINPUT114), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G100), .A2(n871), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G112), .A2(n875), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U961 ( .A1(n860), .A2(n859), .ZN(G162) );
  NAND2_X1 U962 ( .A1(n874), .A2(G130), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G118), .A2(n875), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G142), .A2(n870), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G106), .A2(n871), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(KEYINPUT45), .B(n865), .Z(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n883) );
  XOR2_X1 U970 ( .A(n869), .B(n868), .Z(n881) );
  NAND2_X1 U971 ( .A1(G139), .A2(n870), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G103), .A2(n871), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n880) );
  NAND2_X1 U974 ( .A1(n874), .A2(G127), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G115), .A2(n875), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n923) );
  XNOR2_X1 U979 ( .A(n881), .B(n923), .ZN(n882) );
  XOR2_X1 U980 ( .A(n883), .B(n882), .Z(n885) );
  XNOR2_X1 U981 ( .A(G164), .B(G160), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n891) );
  XOR2_X1 U983 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n887) );
  XNOR2_X1 U984 ( .A(G162), .B(n935), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U988 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U989 ( .A(G171), .B(G286), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n893), .B(KEYINPUT115), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n716), .B(n894), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U993 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U994 ( .A(G2100), .B(G2096), .Z(n899) );
  XNOR2_X1 U995 ( .A(KEYINPUT42), .B(G2678), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U997 ( .A(KEYINPUT43), .B(G2090), .Z(n901) );
  XNOR2_X1 U998 ( .A(G2067), .B(G2072), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G2078), .B(G2084), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(G227) );
  XOR2_X1 U1003 ( .A(KEYINPUT113), .B(G1976), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G1986), .B(G1956), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1006 ( .A(n908), .B(KEYINPUT41), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G1996), .B(G1991), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1009 ( .A(G1981), .B(G1971), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G1966), .B(G1961), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1012 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1013 ( .A(KEYINPUT112), .B(G2474), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(G229) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n917), .B(KEYINPUT116), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n918), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n919), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT49), .B(n920), .Z(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(KEYINPUT55), .ZN(n970) );
  XNOR2_X1 U1024 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n946) );
  XOR2_X1 U1025 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(n926), .B(KEYINPUT50), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(G2090), .B(G162), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(n929), .B(KEYINPUT117), .ZN(n931) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(KEYINPUT51), .B(n932), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n940) );
  XOR2_X1 U1037 ( .A(G160), .B(G2084), .Z(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n946), .B(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n970), .A2(n947), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n948), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n964) );
  XNOR2_X1 U1045 ( .A(n949), .B(G25), .ZN(n958) );
  XNOR2_X1 U1046 ( .A(G27), .B(n950), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(G28), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(G2072), .B(G33), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n954), .B(KEYINPUT119), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1054 ( .A(n959), .B(G32), .Z(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n965), .B(KEYINPUT120), .ZN(n968) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n966), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(n970), .B(n969), .ZN(n972) );
  INV_X1 U1063 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n973), .ZN(n1029) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT57), .B(n976), .ZN(n996) );
  XNOR2_X1 U1070 ( .A(n977), .B(G1341), .ZN(n993) );
  XOR2_X1 U1071 ( .A(G1348), .B(n716), .Z(n988) );
  INV_X1 U1072 ( .A(G299), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(G1956), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(G1971), .A2(G303), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n523), .A2(n981), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n986), .B(KEYINPUT122), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1081 ( .A(G1961), .B(G301), .Z(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT121), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(KEYINPUT123), .B(n994), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1027) );
  INV_X1 U1088 ( .A(G16), .ZN(n1025) );
  XOR2_X1 U1089 ( .A(G1976), .B(G23), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(G1986), .B(KEYINPUT127), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(n999), .B(G24), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(G22), .B(G1971), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1095 ( .A(KEYINPUT58), .B(n1004), .Z(n1022) );
  XOR2_X1 U1096 ( .A(G1966), .B(G21), .Z(n1015) );
  XOR2_X1 U1097 ( .A(G4), .B(KEYINPUT125), .Z(n1006) );
  XNOR2_X1 U1098 ( .A(G1348), .B(KEYINPUT59), .ZN(n1005) );
  XNOR2_X1 U1099 ( .A(n1006), .B(n1005), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(G1981), .B(G6), .ZN(n1007) );
  NOR2_X1 U1102 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1103 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1104 ( .A(G20), .B(G1956), .ZN(n1011) );
  NOR2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1106 ( .A(KEYINPUT60), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(KEYINPUT124), .B(n1016), .Z(n1017) );
  XNOR2_X1 U1109 ( .A(G5), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1111 ( .A(KEYINPUT126), .B(n1020), .Z(n1021) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

