//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G221), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n187), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G125), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n193), .A2(KEYINPUT77), .A3(G140), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n194), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n197), .B1(new_n202), .B2(new_n196), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n205), .B(new_n197), .C1(new_n202), .C2(new_n196), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G110), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT76), .B1(new_n209), .B2(G128), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n210), .A2(KEYINPUT23), .B1(new_n209), .B2(G128), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n212));
  OAI211_X1 g026(.A(KEYINPUT76), .B(new_n212), .C1(new_n209), .C2(G128), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n208), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(KEYINPUT24), .A2(G110), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT74), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT24), .A2(G110), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT24), .A2(G110), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT74), .B1(new_n220), .B2(new_n215), .ZN(new_n221));
  XNOR2_X1  g035(.A(G119), .B(G128), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT75), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT75), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n219), .A2(new_n221), .A3(new_n225), .A4(new_n222), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n214), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n207), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT64), .B(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n193), .A2(G140), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n195), .A3(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n211), .A2(new_n208), .A3(new_n213), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n222), .B1(new_n219), .B2(new_n221), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n204), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n228), .A2(KEYINPUT78), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT78), .B1(new_n228), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n192), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n234), .A3(new_n191), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n237), .A2(KEYINPUT25), .A3(new_n238), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(G217), .B1(new_n189), .B2(G902), .ZN(new_n245));
  XOR2_X1   g059(.A(new_n245), .B(KEYINPUT73), .Z(new_n246));
  AOI21_X1  g060(.A(KEYINPUT79), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n248));
  INV_X1    g062(.A(new_n246), .ZN(new_n249));
  AOI211_X1 g063(.A(new_n248), .B(new_n249), .C1(new_n242), .C2(new_n243), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n237), .A2(new_n239), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n238), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT80), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT32), .ZN(new_n257));
  NOR2_X1   g071(.A1(G472), .A2(G902), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  INV_X1    g075(.A(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT64), .A2(G146), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT64), .A2(G146), .ZN(new_n268));
  OAI21_X1  g082(.A(G143), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n205), .A2(G143), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AND4_X1   g085(.A1(new_n266), .A2(new_n269), .A3(G128), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n269), .B2(KEYINPUT1), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n205), .A2(G143), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n267), .A2(new_n268), .ZN(new_n277));
  INV_X1    g091(.A(G143), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT69), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n281));
  OR2_X1    g095(.A1(KEYINPUT64), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT64), .A2(G146), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n275), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n266), .B1(new_n229), .B2(G143), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n281), .B(new_n285), .C1(new_n286), .C2(new_n273), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n272), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G137), .ZN(new_n289));
  OR3_X1    g103(.A1(new_n289), .A2(KEYINPUT68), .A3(G134), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(G134), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT68), .B1(new_n289), .B2(G134), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT11), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n289), .A3(G134), .ZN(new_n296));
  INV_X1    g110(.A(G134), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n294), .A2(new_n296), .B1(new_n297), .B2(G137), .ZN(new_n298));
  INV_X1    g112(.A(G131), .ZN(new_n299));
  MUX2_X1   g113(.A(new_n293), .B(new_n298), .S(new_n299), .Z(new_n300));
  OR2_X1    g114(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT2), .B(G113), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(G116), .B(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n209), .A2(G116), .ZN(new_n306));
  INV_X1    g120(.A(G116), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n302), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(KEYINPUT70), .A3(new_n310), .ZN(new_n311));
  OR3_X1    g125(.A1(new_n303), .A2(KEYINPUT70), .A3(new_n304), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n298), .B(new_n299), .ZN(new_n315));
  AND2_X1   g129(.A1(KEYINPUT0), .A2(G128), .ZN(new_n316));
  NOR2_X1   g130(.A1(KEYINPUT0), .A2(G128), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n284), .B2(new_n275), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n269), .A2(new_n271), .A3(new_n316), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n269), .A2(KEYINPUT65), .A3(new_n271), .A4(new_n316), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n319), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n315), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n301), .A2(new_n314), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT28), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n315), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  AOI211_X1 g143(.A(KEYINPUT66), .B(new_n319), .C1(new_n322), .C2(new_n323), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT67), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n319), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n270), .B1(new_n229), .B2(G143), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT65), .B1(new_n333), .B2(new_n316), .ZN(new_n334));
  INV_X1    g148(.A(new_n323), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT66), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n324), .A2(new_n328), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n337), .A2(new_n338), .A3(new_n315), .A4(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n340), .A3(new_n301), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n313), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n265), .B1(new_n327), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n301), .A2(KEYINPUT30), .A3(new_n325), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n313), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT31), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n265), .A4(new_n326), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n265), .A3(new_n326), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT31), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n343), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n350), .A3(KEYINPUT31), .ZN(new_n355));
  AOI211_X1 g169(.A(new_n257), .B(new_n259), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n353), .ZN(new_n357));
  INV_X1    g171(.A(new_n343), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT32), .B1(new_n359), .B2(new_n258), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n301), .A2(new_n325), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n313), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n327), .A2(KEYINPUT29), .A3(new_n265), .A4(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n365), .B2(new_n364), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n347), .A2(new_n326), .ZN(new_n368));
  INV_X1    g182(.A(new_n265), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n327), .A2(new_n342), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n265), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G472), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n256), .B1(new_n361), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n322), .A2(new_n323), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n193), .B1(new_n376), .B2(new_n332), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n193), .B2(new_n288), .ZN(new_n378));
  INV_X1    g192(.A(G953), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G224), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n378), .A2(KEYINPUT90), .A3(KEYINPUT7), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n280), .A2(new_n287), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n333), .A2(new_n266), .A3(G128), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n193), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n336), .A2(G125), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT7), .A4(new_n380), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT3), .B1(new_n390), .B2(G107), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  INV_X1    g206(.A(G107), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G104), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n390), .A2(KEYINPUT81), .A3(G107), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT81), .B1(new_n390), .B2(G107), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n391), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT82), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n393), .B2(G104), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n390), .A2(KEYINPUT81), .A3(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n391), .A4(new_n394), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(G101), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n402), .A2(new_n262), .A3(new_n391), .A4(new_n394), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n406), .A2(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n398), .A2(new_n409), .A3(G101), .A4(new_n404), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n313), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n393), .A2(G104), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n390), .A2(G107), .ZN(new_n413));
  OAI21_X1  g227(.A(G101), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n406), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n306), .A2(KEYINPUT5), .ZN(new_n417));
  INV_X1    g231(.A(G113), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n304), .A2(KEYINPUT5), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n419), .A2(new_n420), .B1(new_n304), .B2(new_n303), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G110), .B(G122), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n411), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT86), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n411), .A2(new_n426), .A3(new_n422), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n380), .ZN(new_n429));
  AOI211_X1 g243(.A(G125), .B(new_n272), .C1(new_n280), .C2(new_n287), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(new_n377), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT7), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n430), .B2(new_n377), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n421), .B(new_n434), .C1(new_n415), .C2(KEYINPUT88), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT87), .B(KEYINPUT8), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n423), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT89), .B1(new_n416), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n421), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n434), .B2(new_n415), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n435), .B(new_n437), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n431), .A2(new_n433), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n389), .A2(new_n428), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n238), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(KEYINPUT91), .A3(new_n238), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n423), .B1(new_n411), .B2(new_n422), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n449), .A2(KEYINPUT6), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n425), .B2(new_n427), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n378), .A2(new_n380), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n431), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n447), .A2(new_n448), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n445), .A2(new_n446), .B1(new_n453), .B2(new_n455), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n458), .A3(new_n448), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(KEYINPUT92), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G214), .B1(G237), .B2(G902), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n458), .B1(new_n461), .B2(new_n448), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n275), .A2(KEYINPUT1), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G128), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n278), .B1(new_n282), .B2(new_n283), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n270), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n272), .B1(new_n472), .B2(KEYINPUT83), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(KEYINPUT83), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n415), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n476), .A2(KEYINPUT10), .ZN(new_n477));
  INV_X1    g291(.A(new_n315), .ZN(new_n478));
  INV_X1    g292(.A(new_n288), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT10), .A3(new_n416), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n408), .A2(new_n324), .A3(new_n410), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(new_n478), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G110), .B(G140), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n379), .A2(G227), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n477), .A2(new_n480), .A3(new_n481), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n315), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n482), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n382), .A2(new_n383), .A3(new_n415), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n269), .A2(new_n271), .B1(new_n469), .B2(G128), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n383), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n416), .B1(new_n495), .B2(new_n474), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT12), .A3(new_n315), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n382), .A2(new_n383), .A3(new_n415), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n476), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n492), .A2(new_n496), .A3(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n315), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT12), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n499), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n478), .B1(new_n497), .B2(new_n500), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT12), .B1(new_n509), .B2(new_n503), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT85), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n491), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(G469), .B(new_n490), .C1(new_n512), .C2(new_n485), .ZN(new_n513));
  INV_X1    g327(.A(G469), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n486), .B1(new_n508), .B2(new_n511), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n485), .B1(new_n489), .B2(new_n482), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(new_n238), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n514), .A2(new_n238), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  XOR2_X1   g334(.A(KEYINPUT9), .B(G234), .Z(new_n521));
  AOI21_X1  g335(.A(new_n188), .B1(new_n521), .B2(new_n238), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n278), .A2(G128), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT95), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n273), .A2(G143), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n297), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(G134), .A3(new_n527), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n531), .A3(G134), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n526), .A2(new_n531), .A3(G134), .A4(new_n527), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n307), .A2(G122), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n307), .A2(G122), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G107), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n536), .A3(new_n393), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n533), .A2(new_n534), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n535), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n544));
  OAI21_X1  g358(.A(G107), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n539), .B(KEYINPUT96), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n529), .A3(new_n530), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n521), .A2(G217), .A3(new_n379), .ZN(new_n551));
  OR3_X1    g365(.A1(new_n541), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n541), .B2(new_n550), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(KEYINPUT98), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(new_n551), .C1(new_n541), .C2(new_n550), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n238), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G478), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n557), .B(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G475), .A2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G113), .B(G122), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(new_n390), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n565));
  AOI21_X1  g379(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT18), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(new_n299), .ZN(new_n569));
  OAI211_X1 g383(.A(KEYINPUT18), .B(G131), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n231), .B1(new_n202), .B2(new_n205), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT93), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT93), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n569), .A2(new_n574), .A3(new_n571), .A4(new_n570), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n577));
  OAI21_X1  g391(.A(G131), .B1(new_n565), .B2(new_n566), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n204), .B(new_n206), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n567), .A2(new_n299), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n578), .ZN(new_n581));
  OAI22_X1  g395(.A1(new_n579), .A2(KEYINPUT94), .B1(KEYINPUT17), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n564), .B(new_n576), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT19), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n195), .A2(new_n230), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n202), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n581), .B(new_n204), .C1(new_n277), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n576), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n564), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n562), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT20), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n576), .B1(new_n582), .B2(new_n583), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n590), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n596), .A2(new_n584), .ZN(new_n597));
  OAI21_X1  g411(.A(G475), .B1(new_n597), .B2(G902), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n379), .A2(G952), .ZN(new_n600));
  INV_X1    g414(.A(G237), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n600), .B1(new_n189), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n238), .B(new_n379), .C1(G234), .C2(G237), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT21), .B(G898), .Z(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n560), .A2(new_n599), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n468), .A2(new_n524), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n375), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  NAND2_X1  g426(.A1(new_n244), .A2(new_n246), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n248), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n244), .A2(KEYINPUT79), .A3(new_n246), .ZN(new_n615));
  AND4_X1   g429(.A1(new_n614), .A2(new_n615), .A3(new_n255), .A4(new_n523), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n520), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n359), .A2(new_n258), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n354), .B2(new_n355), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n607), .ZN(new_n622));
  AND4_X1   g436(.A1(new_n458), .A2(new_n447), .A3(new_n448), .A4(new_n456), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n464), .B(new_n622), .C1(new_n623), .C2(new_n465), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n557), .A2(new_n558), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n553), .A2(KEYINPUT99), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n553), .A2(KEYINPUT99), .ZN(new_n627));
  OAI211_X1 g441(.A(KEYINPUT33), .B(new_n552), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n554), .A2(new_n629), .A3(new_n556), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n238), .A2(G478), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n625), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n599), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT100), .B1(new_n624), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n464), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n460), .B2(new_n462), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n638));
  INV_X1    g452(.A(new_n634), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n637), .A2(new_n638), .A3(new_n622), .A4(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n617), .B(new_n621), .C1(new_n635), .C2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT101), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT34), .B(G104), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NOR3_X1   g458(.A1(new_n621), .A2(new_n607), .A3(new_n617), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n598), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g461(.A(KEYINPUT102), .B(G475), .C1(new_n597), .C2(G902), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n647), .A2(new_n594), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n645), .A2(new_n560), .A3(new_n637), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT103), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT35), .B(G107), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n524), .A2(new_n609), .ZN(new_n654));
  INV_X1    g468(.A(new_n468), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n259), .B1(new_n354), .B2(new_n355), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n359), .A2(new_n238), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(G472), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n235), .A2(new_n236), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n659), .B(new_n660), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n254), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n614), .A2(new_n615), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n251), .A2(KEYINPUT104), .A3(new_n662), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n654), .A2(new_n655), .A3(new_n658), .A4(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  NAND4_X1  g484(.A1(new_n560), .A2(new_n647), .A3(new_n594), .A4(new_n648), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n604), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n602), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n663), .A2(new_n664), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT104), .B1(new_n251), .B2(new_n662), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n676), .B(new_n637), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n618), .A2(new_n257), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n656), .A2(KEYINPUT32), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n374), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n498), .B1(new_n510), .B2(KEYINPUT85), .ZN(new_n684));
  AOI211_X1 g498(.A(new_n507), .B(KEYINPUT12), .C1(new_n509), .C2(new_n503), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n487), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n516), .ZN(new_n687));
  AOI21_X1  g501(.A(G902), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n518), .B1(new_n688), .B2(new_n514), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n522), .B1(new_n689), .B2(new_n513), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n680), .A2(new_n683), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  NAND2_X1  g506(.A1(new_n463), .A2(new_n467), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT38), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n674), .B(KEYINPUT39), .Z(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  INV_X1    g513(.A(new_n560), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n594), .A2(new_n598), .ZN(new_n701));
  NOR4_X1   g515(.A1(new_n663), .A2(new_n700), .A3(new_n636), .A4(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n695), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n368), .A2(new_n369), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n326), .A2(new_n369), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(G902), .B1(new_n707), .B2(new_n363), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(G472), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n681), .A2(new_n682), .A3(new_n710), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n704), .B(new_n711), .C1(KEYINPUT40), .C2(new_n698), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  OAI21_X1  g527(.A(new_n464), .B1(new_n623), .B2(new_n465), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n666), .B2(new_n665), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n634), .A2(new_n675), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n683), .A2(new_n715), .A3(new_n690), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  OR2_X1    g532(.A1(new_n688), .A2(new_n514), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n523), .A3(new_n517), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n635), .B2(new_n640), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n375), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NOR4_X1   g538(.A1(new_n720), .A2(new_n714), .A3(new_n607), .A4(new_n671), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n375), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT105), .B(G116), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G18));
  INV_X1    g542(.A(new_n720), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n683), .A2(new_n715), .A3(new_n608), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  NOR3_X1   g545(.A1(new_n624), .A2(new_n701), .A3(new_n700), .ZN(new_n732));
  INV_X1    g546(.A(new_n256), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n327), .A2(new_n363), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n353), .B(new_n349), .C1(new_n265), .C2(new_n734), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n657), .A2(G472), .B1(new_n258), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n732), .A2(new_n733), .A3(new_n729), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n720), .A2(new_n714), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n663), .A3(new_n736), .A4(new_n716), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT106), .B(G125), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G27));
  AND3_X1   g556(.A1(new_n693), .A2(new_n690), .A3(new_n464), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n733), .A3(new_n683), .A4(new_n716), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n375), .A2(KEYINPUT42), .A3(new_n716), .A4(new_n743), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  AND4_X1   g563(.A1(new_n733), .A2(new_n743), .A3(new_n683), .A4(new_n676), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n297), .ZN(G36));
  OAI21_X1  g565(.A(new_n482), .B1(new_n684), .B2(new_n685), .ZN(new_n752));
  INV_X1    g566(.A(new_n485), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n752), .A2(new_n753), .B1(new_n489), .B2(new_n487), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(G469), .A3(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(KEYINPUT107), .Z(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n518), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n759), .A2(KEYINPUT46), .B1(new_n514), .B2(new_n688), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n522), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n621), .A2(KEYINPUT108), .A3(new_n663), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n701), .A2(new_n633), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT43), .Z(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT108), .B1(new_n621), .B2(new_n663), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n764), .A2(new_n697), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n771), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n464), .A3(new_n693), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n289), .ZN(G39));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(KEYINPUT109), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(KEYINPUT109), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n764), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n762), .A2(new_n763), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n523), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n779), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n693), .A2(new_n464), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n716), .A2(new_n256), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n683), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT110), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  AND2_X1   g606(.A1(new_n719), .A2(new_n517), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT49), .ZN(new_n794));
  INV_X1    g608(.A(new_n711), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n256), .A2(new_n766), .A3(new_n636), .A4(new_n522), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n694), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n787), .A2(new_n602), .A3(new_n720), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n795), .A3(new_n733), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n600), .B1(new_n799), .B2(new_n634), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n767), .ZN(new_n801));
  INV_X1    g615(.A(new_n375), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT48), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n767), .A2(new_n603), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n736), .A2(new_n733), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n800), .B(new_n804), .C1(new_n739), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n807), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n783), .A2(new_n786), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n793), .A2(new_n522), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n787), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n799), .A2(new_n599), .A3(new_n633), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n807), .A2(new_n636), .A3(new_n694), .A4(new_n729), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT50), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n736), .A2(new_n663), .ZN(new_n816));
  INV_X1    g630(.A(new_n801), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n813), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT51), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n808), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n809), .A2(new_n787), .ZN(new_n821));
  INV_X1    g635(.A(new_n810), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n811), .B(KEYINPUT115), .Z(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT51), .B1(new_n824), .B2(new_n818), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n750), .B1(new_n746), .B2(new_n747), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT111), .B1(new_n633), .B2(new_n599), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n634), .B1(new_n700), .B2(new_n599), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n828), .B2(KEYINPUT111), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n468), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n375), .A2(new_n725), .B1(new_n645), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n375), .B1(new_n721), .B2(new_n610), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n560), .A2(new_n675), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n649), .B(new_n834), .C1(new_n677), .C2(new_n678), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n361), .B2(new_n374), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n736), .A2(new_n663), .A3(new_n716), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n743), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n730), .A2(new_n737), .A3(new_n668), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n826), .A2(new_n833), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n614), .A2(new_n615), .A3(new_n662), .A4(new_n674), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT112), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n700), .A2(new_n701), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n251), .A2(new_n845), .A3(new_n662), .A4(new_n674), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n637), .A2(new_n843), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n711), .A3(new_n690), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n691), .A2(new_n717), .A3(new_n848), .A4(new_n740), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n637), .B(new_n716), .C1(new_n677), .C2(new_n678), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n683), .B(new_n690), .C1(new_n680), .C2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n740), .A4(new_n848), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n840), .A2(new_n841), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n750), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n748), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n839), .A2(new_n838), .A3(new_n832), .A4(new_n831), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n850), .A2(new_n862), .A3(new_n855), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n850), .B2(new_n855), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n841), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n857), .B1(new_n866), .B2(KEYINPUT114), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n865), .A2(new_n869), .A3(new_n841), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n841), .B1(new_n840), .B2(new_n856), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n865), .B2(new_n841), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n820), .A2(new_n825), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT116), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n797), .B1(new_n876), .B2(new_n878), .ZN(G75));
  NOR2_X1   g693(.A1(new_n379), .A2(G952), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n856), .A2(KEYINPUT113), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n850), .A2(new_n862), .A3(new_n855), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n840), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT114), .B1(new_n884), .B2(KEYINPUT53), .ZN(new_n885));
  INV_X1    g699(.A(new_n857), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n870), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(G210), .A3(G902), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n453), .B(new_n455), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  AOI22_X1  g705(.A1(new_n888), .A2(new_n889), .B1(KEYINPUT117), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(KEYINPUT117), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n881), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n892), .B2(new_n893), .ZN(G51));
  NAND2_X1  g709(.A1(new_n887), .A2(KEYINPUT54), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n871), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n518), .B(KEYINPUT57), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n516), .B2(new_n515), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n887), .A2(G902), .A3(new_n758), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n880), .B1(new_n900), .B2(new_n901), .ZN(G54));
  AND4_X1   g716(.A1(KEYINPUT58), .A2(new_n887), .A3(G475), .A4(G902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n584), .A2(new_n591), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n881), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n904), .B2(new_n903), .ZN(G60));
  XNOR2_X1  g720(.A(new_n631), .B(KEYINPUT118), .ZN(new_n907));
  NAND2_X1  g721(.A1(G478), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT59), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT119), .B1(new_n897), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n913), .B(new_n910), .C1(new_n896), .C2(new_n871), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n907), .B1(new_n875), .B2(new_n909), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n912), .A2(new_n914), .A3(new_n915), .A4(new_n880), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT60), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n252), .B1(new_n887), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT121), .B1(new_n920), .B2(new_n880), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n867), .B2(new_n870), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n922), .B(new_n881), .C1(new_n923), .C2(new_n252), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n661), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n920), .A2(new_n880), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(KEYINPUT61), .A3(new_n925), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(G66));
  AOI21_X1  g745(.A(new_n379), .B1(new_n605), .B2(G224), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n833), .A2(new_n839), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n379), .ZN(new_n934));
  OAI221_X1 g748(.A(new_n450), .B1(G898), .B2(new_n379), .C1(new_n451), .C2(new_n452), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(G69));
  NAND2_X1  g750(.A1(new_n345), .A2(new_n346), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(new_n587), .Z(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT122), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n853), .A2(new_n740), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n712), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n712), .A2(KEYINPUT62), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n791), .A2(new_n946), .ZN(new_n947));
  OR4_X1    g761(.A1(new_n802), .A2(new_n698), .A3(new_n787), .A4(new_n829), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n773), .B2(new_n775), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT123), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n951), .B(new_n948), .C1(new_n773), .C2(new_n775), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n939), .B1(new_n953), .B2(G953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n764), .A2(new_n697), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n375), .A2(new_n637), .A3(new_n844), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n941), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n776), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n958), .A2(new_n379), .A3(new_n791), .A4(new_n826), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n938), .B1(G900), .B2(G953), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n379), .B1(G227), .B2(G900), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n959), .A2(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n961), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n954), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n954), .B2(new_n963), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(G72));
  INV_X1    g782(.A(new_n705), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n620), .A2(new_n238), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n873), .A2(new_n370), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n972), .ZN(new_n974));
  INV_X1    g788(.A(new_n933), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n953), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n973), .B1(new_n976), .B2(new_n969), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n958), .A2(new_n791), .A3(new_n826), .A4(new_n975), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(new_n972), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n370), .B(KEYINPUT126), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  OAI211_X1 g795(.A(KEYINPUT127), .B(new_n881), .C1(new_n979), .C2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n978), .B2(new_n972), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n880), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n977), .B1(new_n982), .B2(new_n985), .ZN(G57));
endmodule


