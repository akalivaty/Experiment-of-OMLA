

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X2 U556 ( .A1(G2104), .A2(n551), .ZN(n903) );
  XOR2_X1 U557 ( .A(KEYINPUT70), .B(n581), .Z(n524) );
  NOR2_X1 U558 ( .A1(n753), .A2(n754), .ZN(n525) );
  XOR2_X1 U559 ( .A(n748), .B(KEYINPUT97), .Z(n526) );
  INV_X1 U560 ( .A(KEYINPUT31), .ZN(n696) );
  INV_X1 U561 ( .A(KEYINPUT95), .ZN(n740) );
  NOR2_X1 U562 ( .A1(G1966), .A2(n805), .ZN(n729) );
  INV_X1 U563 ( .A(KEYINPUT99), .ZN(n758) );
  NOR2_X1 U564 ( .A1(G543), .A2(n533), .ZN(n534) );
  XNOR2_X1 U565 ( .A(KEYINPUT15), .B(n585), .ZN(n984) );
  NOR2_X1 U566 ( .A1(G651), .A2(n649), .ZN(n642) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n632) );
  NAND2_X1 U568 ( .A1(n632), .A2(G89), .ZN(n527) );
  XNOR2_X1 U569 ( .A(n527), .B(KEYINPUT4), .ZN(n529) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n649) );
  INV_X1 U571 ( .A(G651), .ZN(n533) );
  NOR2_X1 U572 ( .A1(n649), .A2(n533), .ZN(n635) );
  NAND2_X1 U573 ( .A1(G76), .A2(n635), .ZN(n528) );
  NAND2_X1 U574 ( .A1(n529), .A2(n528), .ZN(n532) );
  XOR2_X1 U575 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n530) );
  XNOR2_X1 U576 ( .A(KEYINPUT5), .B(n530), .ZN(n531) );
  XNOR2_X1 U577 ( .A(n532), .B(n531), .ZN(n539) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n534), .Z(n647) );
  NAND2_X1 U579 ( .A1(G63), .A2(n647), .ZN(n536) );
  NAND2_X1 U580 ( .A1(G51), .A2(n642), .ZN(n535) );
  NAND2_X1 U581 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U582 ( .A(KEYINPUT6), .B(n537), .Z(n538) );
  NAND2_X1 U583 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U584 ( .A(KEYINPUT7), .B(n540), .ZN(G168) );
  XNOR2_X1 U585 ( .A(G168), .B(KEYINPUT8), .ZN(n541) );
  XNOR2_X1 U586 ( .A(n541), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U587 ( .A1(G72), .A2(n635), .ZN(n543) );
  NAND2_X1 U588 ( .A1(G85), .A2(n632), .ZN(n542) );
  NAND2_X1 U589 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U590 ( .A1(G60), .A2(n647), .ZN(n545) );
  NAND2_X1 U591 ( .A1(G47), .A2(n642), .ZN(n544) );
  NAND2_X1 U592 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U593 ( .A1(n547), .A2(n546), .ZN(G290) );
  AND2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n904) );
  NAND2_X1 U595 ( .A1(G114), .A2(n904), .ZN(n556) );
  NOR2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n548) );
  XOR2_X2 U597 ( .A(n548), .B(KEYINPUT17), .Z(n907) );
  NAND2_X1 U598 ( .A1(G138), .A2(n907), .ZN(n550) );
  INV_X1 U599 ( .A(G2105), .ZN(n551) );
  AND2_X1 U600 ( .A1(n551), .A2(G2104), .ZN(n909) );
  NAND2_X1 U601 ( .A1(G102), .A2(n909), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U603 ( .A1(n903), .A2(G126), .ZN(n552) );
  XOR2_X1 U604 ( .A(KEYINPUT84), .B(n552), .Z(n553) );
  NAND2_X1 U605 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U606 ( .A(n557), .B(KEYINPUT85), .ZN(G164) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(G7), .A2(G661), .ZN(n558) );
  XOR2_X1 U612 ( .A(n558), .B(KEYINPUT10), .Z(n829) );
  NAND2_X1 U613 ( .A1(n829), .A2(G567), .ZN(n559) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  XOR2_X1 U615 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n561) );
  NAND2_X1 U616 ( .A1(G56), .A2(n647), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n561), .B(n560), .ZN(n568) );
  NAND2_X1 U618 ( .A1(n635), .A2(G68), .ZN(n562) );
  XNOR2_X1 U619 ( .A(KEYINPUT69), .B(n562), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n632), .A2(G81), .ZN(n563) );
  XOR2_X1 U621 ( .A(KEYINPUT12), .B(n563), .Z(n564) );
  NOR2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U623 ( .A(n566), .B(KEYINPUT13), .ZN(n567) );
  NOR2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n642), .A2(G43), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n978) );
  INV_X1 U627 ( .A(G860), .ZN(n599) );
  OR2_X1 U628 ( .A1(n978), .A2(n599), .ZN(G153) );
  NAND2_X1 U629 ( .A1(G52), .A2(n642), .ZN(n571) );
  XOR2_X1 U630 ( .A(KEYINPUT64), .B(n571), .Z(n578) );
  NAND2_X1 U631 ( .A1(G77), .A2(n635), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G90), .A2(n632), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U634 ( .A(n574), .B(KEYINPUT9), .ZN(n576) );
  NAND2_X1 U635 ( .A1(G64), .A2(n647), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U637 ( .A1(n578), .A2(n577), .ZN(G171) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U640 ( .A1(n642), .A2(G54), .ZN(n584) );
  NAND2_X1 U641 ( .A1(G79), .A2(n635), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G92), .A2(n632), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n647), .A2(G66), .ZN(n581) );
  NOR2_X1 U645 ( .A1(n582), .A2(n524), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U647 ( .A(n984), .ZN(n708) );
  INV_X1 U648 ( .A(G868), .ZN(n663) );
  NAND2_X1 U649 ( .A1(n708), .A2(n663), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U651 ( .A1(n642), .A2(G53), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT66), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G65), .A2(n647), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(KEYINPUT67), .B(n591), .ZN(n596) );
  NAND2_X1 U656 ( .A1(G78), .A2(n635), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G91), .A2(n632), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U659 ( .A(KEYINPUT65), .B(n594), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(G299) );
  NOR2_X1 U661 ( .A1(G286), .A2(n663), .ZN(n598) );
  NOR2_X1 U662 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U663 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U664 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n600), .A2(n984), .ZN(n601) );
  XNOR2_X1 U666 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U667 ( .A1(n984), .A2(G868), .ZN(n602) );
  NOR2_X1 U668 ( .A1(G559), .A2(n602), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n603), .B(KEYINPUT74), .ZN(n605) );
  NOR2_X1 U670 ( .A1(n978), .A2(G868), .ZN(n604) );
  NOR2_X1 U671 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G123), .A2(n903), .ZN(n606) );
  XNOR2_X1 U673 ( .A(n606), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U674 ( .A1(G111), .A2(n904), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G99), .A2(n909), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U677 ( .A(KEYINPUT76), .B(n609), .Z(n610) );
  NAND2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U679 ( .A1(G135), .A2(n907), .ZN(n612) );
  XNOR2_X1 U680 ( .A(KEYINPUT75), .B(n612), .ZN(n613) );
  NOR2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n953) );
  XNOR2_X1 U682 ( .A(G2096), .B(n953), .ZN(n615) );
  INV_X1 U683 ( .A(G2100), .ZN(n865) );
  NAND2_X1 U684 ( .A1(n615), .A2(n865), .ZN(G156) );
  NAND2_X1 U685 ( .A1(G67), .A2(n647), .ZN(n617) );
  NAND2_X1 U686 ( .A1(G93), .A2(n632), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U688 ( .A1(G80), .A2(n635), .ZN(n618) );
  XNOR2_X1 U689 ( .A(KEYINPUT77), .B(n618), .ZN(n619) );
  NOR2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n642), .A2(G55), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n662) );
  NAND2_X1 U693 ( .A1(n984), .A2(G559), .ZN(n660) );
  XNOR2_X1 U694 ( .A(n978), .B(n660), .ZN(n623) );
  NOR2_X1 U695 ( .A1(G860), .A2(n623), .ZN(n624) );
  XOR2_X1 U696 ( .A(n662), .B(n624), .Z(G145) );
  NAND2_X1 U697 ( .A1(G88), .A2(n632), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G50), .A2(n642), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G62), .A2(n647), .ZN(n628) );
  NAND2_X1 U701 ( .A1(G75), .A2(n635), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U704 ( .A(n631), .B(KEYINPUT81), .Z(G166) );
  INV_X1 U705 ( .A(G166), .ZN(G303) );
  NAND2_X1 U706 ( .A1(G61), .A2(n647), .ZN(n634) );
  NAND2_X1 U707 ( .A1(G86), .A2(n632), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U710 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n642), .A2(G48), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U714 ( .A1(G651), .A2(G74), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(KEYINPUT78), .ZN(n644) );
  NAND2_X1 U716 ( .A1(G49), .A2(n642), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U718 ( .A(KEYINPUT79), .B(n645), .Z(n646) );
  NOR2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n648), .B(KEYINPUT80), .ZN(n651) );
  NAND2_X1 U721 ( .A1(G87), .A2(n649), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(G288) );
  XNOR2_X1 U723 ( .A(KEYINPUT19), .B(KEYINPUT83), .ZN(n653) );
  XNOR2_X1 U724 ( .A(G290), .B(KEYINPUT82), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n654), .B(G305), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n655), .B(n662), .ZN(n656) );
  XOR2_X1 U728 ( .A(G303), .B(n656), .Z(n659) );
  XOR2_X1 U729 ( .A(G299), .B(n978), .Z(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(G288), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n659), .B(n658), .ZN(n872) );
  XNOR2_X1 U732 ( .A(n660), .B(n872), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n661), .A2(G868), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U742 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U743 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U744 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U745 ( .A1(G96), .A2(n672), .ZN(n833) );
  NAND2_X1 U746 ( .A1(n833), .A2(G2106), .ZN(n676) );
  NAND2_X1 U747 ( .A1(G69), .A2(G120), .ZN(n673) );
  NOR2_X1 U748 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U749 ( .A1(G108), .A2(n674), .ZN(n834) );
  NAND2_X1 U750 ( .A1(n834), .A2(G567), .ZN(n675) );
  NAND2_X1 U751 ( .A1(n676), .A2(n675), .ZN(n846) );
  NAND2_X1 U752 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U753 ( .A1(n846), .A2(n677), .ZN(n832) );
  NAND2_X1 U754 ( .A1(n832), .A2(G36), .ZN(G176) );
  NAND2_X1 U755 ( .A1(n904), .A2(G113), .ZN(n680) );
  NAND2_X1 U756 ( .A1(G101), .A2(n909), .ZN(n678) );
  XOR2_X1 U757 ( .A(KEYINPUT23), .B(n678), .Z(n679) );
  NAND2_X1 U758 ( .A1(n680), .A2(n679), .ZN(n684) );
  NAND2_X1 U759 ( .A1(G125), .A2(n903), .ZN(n682) );
  NAND2_X1 U760 ( .A1(G137), .A2(n907), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U762 ( .A1(n684), .A2(n683), .ZN(G160) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n776) );
  INV_X1 U764 ( .A(n776), .ZN(n686) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n777) );
  NOR2_X2 U766 ( .A1(n686), .A2(n777), .ZN(n712) );
  INV_X1 U767 ( .A(n712), .ZN(n734) );
  NOR2_X1 U768 ( .A1(G2084), .A2(n734), .ZN(n690) );
  NAND2_X1 U769 ( .A1(G8), .A2(n690), .ZN(n731) );
  NAND2_X1 U770 ( .A1(G8), .A2(n734), .ZN(n805) );
  NAND2_X1 U771 ( .A1(G1961), .A2(n734), .ZN(n688) );
  XOR2_X1 U772 ( .A(KEYINPUT25), .B(G2078), .Z(n925) );
  NAND2_X1 U773 ( .A1(n712), .A2(n925), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n698) );
  NAND2_X1 U775 ( .A1(G301), .A2(n698), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n689), .B(KEYINPUT93), .ZN(n695) );
  NOR2_X1 U777 ( .A1(n729), .A2(n690), .ZN(n691) );
  NAND2_X1 U778 ( .A1(G8), .A2(n691), .ZN(n692) );
  XNOR2_X1 U779 ( .A(n692), .B(KEYINPUT30), .ZN(n693) );
  NOR2_X1 U780 ( .A1(n693), .A2(G168), .ZN(n694) );
  NOR2_X1 U781 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U782 ( .A(n697), .B(n696), .ZN(n727) );
  OR2_X1 U783 ( .A1(G301), .A2(n698), .ZN(n725) );
  AND2_X1 U784 ( .A1(n712), .A2(G1996), .ZN(n699) );
  XOR2_X1 U785 ( .A(n699), .B(KEYINPUT26), .Z(n701) );
  NAND2_X1 U786 ( .A1(n734), .A2(G1341), .ZN(n700) );
  NAND2_X1 U787 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U788 ( .A1(n978), .A2(n702), .ZN(n706) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n734), .ZN(n704) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n712), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n704), .A2(n703), .ZN(n707) );
  NOR2_X1 U792 ( .A1(n708), .A2(n707), .ZN(n705) );
  OR2_X1 U793 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U794 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U795 ( .A1(n710), .A2(n709), .ZN(n716) );
  INV_X1 U796 ( .A(G299), .ZN(n979) );
  NAND2_X1 U797 ( .A1(n712), .A2(G2072), .ZN(n711) );
  XNOR2_X1 U798 ( .A(n711), .B(KEYINPUT27), .ZN(n714) );
  INV_X1 U799 ( .A(G1956), .ZN(n849) );
  NOR2_X1 U800 ( .A1(n849), .A2(n712), .ZN(n713) );
  NOR2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U802 ( .A1(n979), .A2(n717), .ZN(n715) );
  NAND2_X1 U803 ( .A1(n716), .A2(n715), .ZN(n721) );
  NOR2_X1 U804 ( .A1(n979), .A2(n717), .ZN(n719) );
  XNOR2_X1 U805 ( .A(KEYINPUT28), .B(KEYINPUT91), .ZN(n718) );
  XNOR2_X1 U806 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U807 ( .A1(n721), .A2(n720), .ZN(n723) );
  XOR2_X1 U808 ( .A(KEYINPUT92), .B(KEYINPUT29), .Z(n722) );
  XNOR2_X1 U809 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U811 ( .A1(n727), .A2(n726), .ZN(n732) );
  INV_X1 U812 ( .A(n732), .ZN(n728) );
  NOR2_X1 U813 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U814 ( .A1(n731), .A2(n730), .ZN(n745) );
  NAND2_X1 U815 ( .A1(n732), .A2(G286), .ZN(n739) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n805), .ZN(n733) );
  XNOR2_X1 U817 ( .A(n733), .B(KEYINPUT94), .ZN(n736) );
  NOR2_X1 U818 ( .A1(n734), .A2(G2090), .ZN(n735) );
  NOR2_X1 U819 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U820 ( .A1(n737), .A2(G303), .ZN(n738) );
  NAND2_X1 U821 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U822 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U823 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U824 ( .A(n743), .B(KEYINPUT32), .ZN(n744) );
  NAND2_X1 U825 ( .A1(n745), .A2(n744), .ZN(n799) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n746) );
  NOR2_X1 U828 ( .A1(n750), .A2(n746), .ZN(n998) );
  XNOR2_X1 U829 ( .A(KEYINPUT96), .B(n998), .ZN(n747) );
  NAND2_X1 U830 ( .A1(n799), .A2(n747), .ZN(n748) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U832 ( .A(n987), .ZN(n749) );
  OR2_X1 U833 ( .A1(n805), .A2(n749), .ZN(n753) );
  NAND2_X1 U834 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  NOR2_X1 U835 ( .A1(n805), .A2(n751), .ZN(n752) );
  XNOR2_X1 U836 ( .A(n752), .B(KEYINPUT98), .ZN(n754) );
  NAND2_X1 U837 ( .A1(n526), .A2(n525), .ZN(n757) );
  INV_X1 U838 ( .A(n754), .ZN(n755) );
  NAND2_X1 U839 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  NAND2_X1 U840 ( .A1(n757), .A2(n756), .ZN(n759) );
  XNOR2_X1 U841 ( .A(n759), .B(n758), .ZN(n796) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n993) );
  NAND2_X1 U843 ( .A1(G129), .A2(n903), .ZN(n761) );
  NAND2_X1 U844 ( .A1(G117), .A2(n904), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U846 ( .A1(n909), .A2(G105), .ZN(n762) );
  XOR2_X1 U847 ( .A(KEYINPUT38), .B(n762), .Z(n763) );
  NOR2_X1 U848 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U849 ( .A(n765), .B(KEYINPUT90), .ZN(n767) );
  NAND2_X1 U850 ( .A1(G141), .A2(n907), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n767), .A2(n766), .ZN(n900) );
  AND2_X1 U852 ( .A1(n900), .A2(G1996), .ZN(n775) );
  INV_X1 U853 ( .A(G1991), .ZN(n933) );
  NAND2_X1 U854 ( .A1(G119), .A2(n903), .ZN(n769) );
  NAND2_X1 U855 ( .A1(G107), .A2(n904), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G95), .A2(n909), .ZN(n771) );
  NAND2_X1 U858 ( .A1(G131), .A2(n907), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n885) );
  NOR2_X1 U861 ( .A1(n933), .A2(n885), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n960) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U864 ( .A(n778), .B(KEYINPUT87), .Z(n791) );
  INV_X1 U865 ( .A(n791), .ZN(n821) );
  NOR2_X1 U866 ( .A1(n960), .A2(n821), .ZN(n814) );
  XNOR2_X1 U867 ( .A(KEYINPUT86), .B(G1986), .ZN(n779) );
  XNOR2_X1 U868 ( .A(n779), .B(G290), .ZN(n990) );
  NAND2_X1 U869 ( .A1(n990), .A2(n791), .ZN(n780) );
  XNOR2_X1 U870 ( .A(n780), .B(KEYINPUT88), .ZN(n793) );
  XOR2_X1 U871 ( .A(G2067), .B(KEYINPUT37), .Z(n810) );
  NAND2_X1 U872 ( .A1(G128), .A2(n903), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G116), .A2(n904), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U875 ( .A(n783), .B(KEYINPUT35), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n909), .A2(G104), .ZN(n784) );
  XOR2_X1 U877 ( .A(KEYINPUT89), .B(n784), .Z(n786) );
  NAND2_X1 U878 ( .A1(n907), .A2(G140), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U880 ( .A(KEYINPUT34), .B(n787), .Z(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U882 ( .A(n790), .B(KEYINPUT36), .ZN(n889) );
  NAND2_X1 U883 ( .A1(n810), .A2(n889), .ZN(n817) );
  INV_X1 U884 ( .A(n817), .ZN(n958) );
  NAND2_X1 U885 ( .A1(n958), .A2(n791), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U887 ( .A1(n814), .A2(n794), .ZN(n807) );
  AND2_X1 U888 ( .A1(n993), .A2(n807), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n827) );
  NOR2_X1 U890 ( .A1(G2090), .A2(G303), .ZN(n797) );
  NAND2_X1 U891 ( .A1(G8), .A2(n797), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U893 ( .A(n800), .B(KEYINPUT100), .ZN(n802) );
  AND2_X1 U894 ( .A1(n805), .A2(n807), .ZN(n801) );
  AND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n809) );
  NOR2_X1 U896 ( .A1(G1981), .A2(G305), .ZN(n803) );
  XOR2_X1 U897 ( .A(n803), .B(KEYINPUT24), .Z(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n806) );
  AND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n825) );
  NOR2_X1 U901 ( .A1(n810), .A2(n889), .ZN(n968) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n900), .ZN(n963) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n811) );
  AND2_X1 U904 ( .A1(n933), .A2(n885), .ZN(n954) );
  NOR2_X1 U905 ( .A1(n811), .A2(n954), .ZN(n812) );
  XOR2_X1 U906 ( .A(KEYINPUT101), .B(n812), .Z(n813) );
  NOR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U908 ( .A1(n963), .A2(n815), .ZN(n816) );
  XNOR2_X1 U909 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U911 ( .A(KEYINPUT102), .B(n819), .Z(n820) );
  NOR2_X1 U912 ( .A1(n968), .A2(n820), .ZN(n822) );
  NOR2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U914 ( .A(n823), .B(KEYINPUT103), .ZN(n824) );
  AND2_X1 U915 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U916 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U917 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n829), .ZN(G217) );
  INV_X1 U919 ( .A(n829), .ZN(G223) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U921 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U930 ( .A(KEYINPUT104), .B(G2454), .ZN(n843) );
  XNOR2_X1 U931 ( .A(G2430), .B(G2435), .ZN(n841) );
  XOR2_X1 U932 ( .A(G2451), .B(G2427), .Z(n836) );
  XNOR2_X1 U933 ( .A(G2438), .B(G2446), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n837), .B(G2443), .Z(n839) );
  XNOR2_X1 U936 ( .A(G1341), .B(G1348), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n844), .A2(G14), .ZN(n845) );
  XNOR2_X1 U941 ( .A(KEYINPUT105), .B(n845), .ZN(G401) );
  INV_X1 U942 ( .A(n846), .ZN(G319) );
  XOR2_X1 U943 ( .A(G1961), .B(G1966), .Z(n848) );
  XOR2_X1 U944 ( .A(n933), .B(G1996), .Z(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n859) );
  XOR2_X1 U946 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n851) );
  XOR2_X1 U947 ( .A(n849), .B(KEYINPUT108), .Z(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U949 ( .A(G1976), .B(G1981), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1971), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(G2474), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U955 ( .A(n859), .B(n858), .Z(G229) );
  XOR2_X1 U956 ( .A(G2096), .B(G2678), .Z(n861) );
  XNOR2_X1 U957 ( .A(G2067), .B(KEYINPUT43), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U959 ( .A(n862), .B(KEYINPUT42), .Z(n864) );
  XNOR2_X1 U960 ( .A(G2072), .B(G2090), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(n869) );
  XNOR2_X1 U962 ( .A(KEYINPUT106), .B(n865), .ZN(n867) );
  XNOR2_X1 U963 ( .A(G2078), .B(G2084), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(G227) );
  XOR2_X1 U966 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n871) );
  XOR2_X1 U967 ( .A(G301), .B(G286), .Z(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(n874) );
  XOR2_X1 U969 ( .A(n984), .B(n872), .Z(n873) );
  XNOR2_X1 U970 ( .A(n874), .B(n873), .ZN(n875) );
  NOR2_X1 U971 ( .A1(G37), .A2(n875), .ZN(n876) );
  XOR2_X1 U972 ( .A(KEYINPUT115), .B(n876), .Z(G397) );
  NAND2_X1 U973 ( .A1(n907), .A2(G136), .ZN(n883) );
  NAND2_X1 U974 ( .A1(G112), .A2(n904), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G100), .A2(n909), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n903), .A2(G124), .ZN(n879) );
  XOR2_X1 U978 ( .A(KEYINPUT44), .B(n879), .Z(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  NAND2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U981 ( .A(KEYINPUT110), .B(n884), .Z(G162) );
  XOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n887) );
  XNOR2_X1 U983 ( .A(n885), .B(n953), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(G162), .B(n888), .ZN(n891) );
  XNOR2_X1 U986 ( .A(G164), .B(n889), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n899) );
  NAND2_X1 U988 ( .A1(G103), .A2(n909), .ZN(n893) );
  NAND2_X1 U989 ( .A1(G139), .A2(n907), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n898) );
  NAND2_X1 U991 ( .A1(G127), .A2(n903), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G115), .A2(n904), .ZN(n894) );
  NAND2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U995 ( .A1(n898), .A2(n897), .ZN(n948) );
  XOR2_X1 U996 ( .A(n899), .B(n948), .Z(n902) );
  XOR2_X1 U997 ( .A(n900), .B(G160), .Z(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n916) );
  NAND2_X1 U999 ( .A1(G130), .A2(n903), .ZN(n906) );
  NAND2_X1 U1000 ( .A1(G118), .A2(n904), .ZN(n905) );
  NAND2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n914) );
  NAND2_X1 U1002 ( .A1(n907), .A2(G142), .ZN(n908) );
  XOR2_X1 U1003 ( .A(KEYINPUT111), .B(n908), .Z(n911) );
  NAND2_X1 U1004 ( .A1(n909), .A2(G106), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1006 ( .A(n912), .B(KEYINPUT45), .Z(n913) );
  NOR2_X1 U1007 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1008 ( .A(n916), .B(n915), .Z(n917) );
  NOR2_X1 U1009 ( .A1(n917), .A2(G37), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(n918), .B(KEYINPUT112), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n919) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n919), .Z(n920) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n920), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1015 ( .A(KEYINPUT116), .B(n922), .ZN(n924) );
  NOR2_X1 U1016 ( .A1(G397), .A2(G395), .ZN(n923) );
  NAND2_X1 U1017 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1020 ( .A(G32), .B(G1996), .Z(n929) );
  XNOR2_X1 U1021 ( .A(G2067), .B(G26), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(G27), .B(n925), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(G33), .B(G2072), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1027 ( .A(KEYINPUT120), .B(n932), .Z(n935) );
  XOR2_X1 U1028 ( .A(n933), .B(G25), .Z(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(G28), .A2(n936), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(KEYINPUT53), .B(n937), .ZN(n939) );
  XOR2_X1 U1032 ( .A(G2090), .B(G35), .Z(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(KEYINPUT121), .B(n940), .ZN(n944) );
  XOR2_X1 U1035 ( .A(KEYINPUT122), .B(G34), .Z(n942) );
  XNOR2_X1 U1036 ( .A(G2084), .B(KEYINPUT54), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(n942), .B(n941), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1039 ( .A(KEYINPUT55), .B(n945), .Z(n946) );
  INV_X1 U1040 ( .A(G29), .ZN(n974) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n974), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(G11), .A2(n947), .ZN(n977) );
  XNOR2_X1 U1043 ( .A(G2072), .B(n948), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(n949), .B(KEYINPUT119), .ZN(n951) );
  XOR2_X1 U1045 ( .A(G2078), .B(G164), .Z(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1047 ( .A(KEYINPUT50), .B(n952), .Z(n971) );
  XNOR2_X1 U1048 ( .A(G160), .B(G2084), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(KEYINPUT117), .B(n961), .ZN(n966) );
  XOR2_X1 U1054 ( .A(G2090), .B(G162), .Z(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1056 ( .A(KEYINPUT51), .B(n964), .Z(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1059 ( .A(KEYINPUT118), .B(n969), .Z(n970) );
  NOR2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1061 ( .A(KEYINPUT52), .B(n972), .Z(n973) );
  NOR2_X1 U1062 ( .A1(KEYINPUT55), .A2(n973), .ZN(n975) );
  NOR2_X1 U1063 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1064 ( .A1(n977), .A2(n976), .ZN(n1029) );
  XNOR2_X1 U1065 ( .A(n978), .B(G1341), .ZN(n981) );
  XOR2_X1 U1066 ( .A(n979), .B(G1956), .Z(n980) );
  NOR2_X1 U1067 ( .A1(n981), .A2(n980), .ZN(n992) );
  XOR2_X1 U1068 ( .A(G301), .B(G1961), .Z(n983) );
  NAND2_X1 U1069 ( .A1(G1971), .A2(G303), .ZN(n982) );
  NAND2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1071 ( .A(G1348), .B(n984), .Z(n985) );
  NOR2_X1 U1072 ( .A1(n986), .A2(n985), .ZN(n988) );
  NAND2_X1 U1073 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1074 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1075 ( .A1(n992), .A2(n991), .ZN(n1000) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n994) );
  NAND2_X1 U1077 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1078 ( .A(n995), .B(KEYINPUT57), .ZN(n996) );
  XOR2_X1 U1079 ( .A(KEYINPUT123), .B(n996), .Z(n997) );
  NAND2_X1 U1080 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1081 ( .A1(n1000), .A2(n999), .ZN(n1030) );
  INV_X1 U1082 ( .A(n1030), .ZN(n1001) );
  NAND2_X1 U1083 ( .A1(n1001), .A2(KEYINPUT56), .ZN(n1026) );
  XOR2_X1 U1084 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n1024) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G21), .ZN(n1003) );
  XNOR2_X1 U1086 ( .A(G5), .B(G1961), .ZN(n1002) );
  NOR2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1022) );
  XOR2_X1 U1088 ( .A(G1971), .B(KEYINPUT126), .Z(n1004) );
  XNOR2_X1 U1089 ( .A(G22), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G23), .B(G1976), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(n1009), .B(KEYINPUT58), .ZN(n1020) );
  XNOR2_X1 U1095 ( .A(KEYINPUT59), .B(G1348), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(n1010), .B(G4), .ZN(n1016) );
  XOR2_X1 U1097 ( .A(G1341), .B(G19), .Z(n1012) );
  XOR2_X1 U1098 ( .A(G1956), .B(G20), .Z(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G6), .B(G1981), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(n1017), .B(KEYINPUT60), .Z(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT125), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(n1024), .B(n1023), .ZN(n1031) );
  OR2_X1 U1108 ( .A1(n1031), .A2(KEYINPUT124), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(G16), .ZN(n1028) );
  NAND2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1037) );
  NOR2_X1 U1112 ( .A1(KEYINPUT56), .A2(n1030), .ZN(n1034) );
  INV_X1 U1113 ( .A(KEYINPUT124), .ZN(n1032) );
  NOR2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1115 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1116 ( .A1(G16), .A2(n1035), .ZN(n1036) );
  NOR2_X1 U1117 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1118 ( .A(n1038), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

