//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n202), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n212), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n219), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  OAI21_X1  g0046(.A(KEYINPUT72), .B1(new_n246), .B2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT72), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n246), .A2(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n247), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n207), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(KEYINPUT73), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT73), .B1(new_n253), .B2(new_n254), .ZN(new_n258));
  OAI21_X1  g0058(.A(G68), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G58), .ZN(new_n260));
  INV_X1    g0060(.A(G68), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n262), .B2(new_n201), .ZN(new_n263));
  INV_X1    g0063(.A(G159), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  XOR2_X1   g0067(.A(new_n267), .B(KEYINPUT74), .Z(new_n268));
  NAND3_X1  g0068(.A1(new_n259), .A2(new_n268), .A3(KEYINPUT16), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n267), .B(KEYINPUT74), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n207), .B1(KEYINPUT76), .B2(KEYINPUT7), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n251), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT76), .ZN(new_n279));
  AOI21_X1  g0079(.A(G20), .B1(new_n279), .B2(new_n254), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(new_n272), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n276), .A2(new_n281), .A3(G68), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n270), .B1(new_n271), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n213), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n269), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n285), .B1(new_n206), .B2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(new_n293), .B2(new_n288), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G226), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(G1698), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n299), .A2(new_n247), .A3(new_n250), .A4(new_n251), .ZN(new_n300));
  INV_X1    g0100(.A(G87), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n249), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT77), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(KEYINPUT77), .C1(new_n249), .C2(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT78), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G41), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(G1), .A3(G13), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G232), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G41), .ZN(new_n314));
  INV_X1    g0114(.A(G45), .ZN(new_n315));
  AOI21_X1  g0115(.A(G1), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G274), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT79), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n302), .A2(new_n303), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT78), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(new_n306), .A4(new_n305), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n308), .A2(new_n309), .A3(new_n320), .A4(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n318), .B1(new_n304), .B2(new_n307), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n296), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT18), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT18), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n296), .A2(new_n332), .A3(new_n329), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n308), .A2(new_n334), .A3(new_n320), .A4(new_n323), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n286), .A2(new_n338), .A3(new_n295), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT17), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n286), .A2(new_n338), .A3(KEYINPUT17), .A4(new_n295), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n331), .A2(new_n333), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n265), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n207), .A2(G33), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n287), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n285), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n289), .A2(new_n202), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n292), .B2(new_n202), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(KEYINPUT9), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g0150(.A(new_n350), .B(KEYINPUT69), .Z(new_n351));
  INV_X1    g0151(.A(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n274), .A2(G222), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n274), .A2(G1698), .ZN(new_n355));
  OAI221_X1 g0155(.A(new_n353), .B1(new_n354), .B2(new_n274), .C1(new_n355), .C2(new_n298), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n306), .ZN(new_n357));
  INV_X1    g0157(.A(new_n317), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n306), .A2(new_n316), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(G226), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT9), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n347), .A2(new_n349), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n362), .A2(G190), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(G200), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n351), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT10), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT10), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n351), .A2(new_n365), .A3(new_n369), .A4(new_n366), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n311), .A2(G238), .A3(new_n312), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n317), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n277), .A2(new_n251), .A3(G226), .A4(new_n352), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n277), .A2(new_n251), .A3(G232), .A4(G1698), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G97), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI211_X1 g0177(.A(KEYINPUT13), .B(new_n373), .C1(new_n306), .C2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n306), .ZN(new_n380));
  INV_X1    g0180(.A(new_n373), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(G169), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT70), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n373), .B1(new_n377), .B2(new_n306), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n379), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT70), .B1(new_n387), .B2(new_n379), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n386), .A2(G179), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT14), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(G169), .C1(new_n378), .C2(new_n382), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n384), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n266), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n345), .A2(new_n354), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n285), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT11), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n396), .A2(new_n397), .B1(G68), .B2(new_n292), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n206), .A2(G13), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n400), .A2(new_n207), .A3(G68), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT12), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT71), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(KEYINPUT71), .A3(new_n402), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n402), .B2(new_n401), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n398), .B(new_n399), .C1(new_n403), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n393), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n387), .B(new_n379), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n408), .B2(G200), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n386), .A2(G190), .A3(new_n388), .A4(new_n389), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n288), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT68), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n413), .A2(new_n414), .B1(new_n345), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n413), .A2(new_n414), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n285), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n289), .A2(new_n354), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n292), .B2(new_n354), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n274), .A2(G232), .A3(new_n352), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  INV_X1    g0224(.A(G238), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n423), .B1(new_n424), .B2(new_n274), .C1(new_n355), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n306), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n358), .B1(new_n359), .B2(G244), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(G200), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n429), .A2(G190), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n422), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n362), .A2(new_n326), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n361), .A2(new_n309), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n364), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(G169), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n429), .A2(new_n309), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n421), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n433), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  NOR4_X1   g0241(.A1(new_n343), .A2(new_n371), .A3(new_n412), .A4(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT5), .B(G41), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n315), .A2(G1), .ZN(new_n444));
  INV_X1    g0244(.A(new_n213), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n443), .A2(new_n444), .B1(new_n445), .B2(new_n310), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT86), .B1(new_n446), .B2(G264), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n206), .A2(G45), .ZN(new_n448));
  OR2_X1    g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NAND2_X1  g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT86), .ZN(new_n452));
  INV_X1    g0252(.A(G264), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n451), .A2(new_n306), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G257), .A2(G1698), .ZN(new_n456));
  INV_X1    g0256(.A(G250), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G1698), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(new_n247), .A3(new_n250), .A4(new_n251), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G294), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n306), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n451), .A2(G274), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n455), .A2(new_n334), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n444), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n311), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n452), .B1(new_n468), .B2(new_n453), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n446), .A2(KEYINPUT86), .A3(G264), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n462), .A2(new_n469), .A3(new_n470), .A4(new_n463), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n336), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n285), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n424), .A2(KEYINPUT23), .A3(G20), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT23), .B1(new_n424), .B2(G20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G116), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n475), .A2(new_n476), .B1(G20), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT22), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(new_n207), .A3(G87), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT85), .B1(new_n278), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n480), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT85), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n274), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n247), .A2(new_n250), .A3(new_n207), .A4(new_n251), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT22), .B1(new_n486), .B2(new_n301), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n478), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n474), .B1(new_n488), .B2(KEYINPUT24), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT24), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(KEYINPUT72), .B2(new_n277), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n207), .A3(G87), .A4(new_n250), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n493), .A2(KEYINPUT22), .B1(new_n484), .B2(new_n481), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n490), .B1(new_n494), .B2(new_n478), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n400), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G20), .A3(new_n424), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT25), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n206), .A2(G33), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n289), .A2(new_n500), .A3(new_n213), .A4(new_n284), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n499), .B1(G107), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n473), .A2(new_n496), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n311), .B1(new_n459), .B2(new_n460), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n447), .A2(new_n454), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G179), .A3(new_n463), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n471), .A2(G169), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n496), .A2(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT87), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n496), .A2(new_n503), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT87), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n473), .A2(new_n496), .A3(new_n503), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  AND2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n424), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(G20), .B1(G77), .B2(new_n265), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n276), .A2(new_n281), .A3(G107), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n285), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n289), .A2(G97), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n502), .B2(G97), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n518), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n474), .B1(new_n525), .B2(new_n526), .ZN(new_n532));
  INV_X1    g0332(.A(new_n530), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n532), .A2(KEYINPUT81), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G257), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n463), .B1(new_n468), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n277), .A2(new_n251), .A3(G250), .A4(G1698), .ZN(new_n538));
  AND2_X1   g0338(.A1(KEYINPUT4), .A2(G244), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n277), .A2(new_n251), .A3(new_n539), .A4(new_n352), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G283), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n247), .A2(new_n250), .A3(G244), .A4(new_n251), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(G1698), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n537), .B1(new_n546), .B2(new_n306), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n309), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n311), .B1(new_n542), .B2(new_n545), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n326), .B1(new_n549), .B2(new_n537), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT82), .B1(new_n535), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n548), .A2(new_n550), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT82), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n528), .A2(new_n518), .A3(new_n530), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT81), .B1(new_n532), .B2(new_n533), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n547), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT80), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(G200), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT80), .B1(new_n547), .B2(new_n336), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n547), .A2(G190), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n532), .A2(new_n533), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n552), .A2(new_n558), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT21), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n289), .A2(G116), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n502), .B2(G116), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n249), .A2(G97), .ZN(new_n571));
  AOI21_X1  g0371(.A(G20), .B1(new_n571), .B2(new_n541), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n207), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n285), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n570), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G169), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n247), .A2(new_n250), .A3(new_n352), .A4(new_n251), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n581), .A2(new_n536), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n278), .A2(G303), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT84), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n453), .A2(new_n352), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n492), .A2(new_n584), .A3(new_n250), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G264), .A2(G1698), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT84), .B1(new_n252), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n582), .A2(new_n583), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n467), .A2(G270), .A3(new_n311), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n463), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT83), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT83), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n463), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n589), .A2(new_n306), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n568), .B1(new_n580), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n586), .A2(new_n588), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n583), .B1(new_n581), .B2(new_n536), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n306), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n592), .A2(new_n594), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n601), .A2(KEYINPUT21), .A3(G169), .A4(new_n579), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(G179), .A3(new_n579), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n596), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n336), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n595), .A2(new_n334), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n579), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n477), .B1(new_n544), .B2(new_n352), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n581), .A2(new_n425), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n306), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n444), .B2(new_n457), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n311), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n309), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n415), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n289), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n207), .B1(new_n376), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(G97), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n301), .A2(new_n619), .A3(new_n424), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n618), .A2(new_n620), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n261), .B2(new_n486), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n616), .B1(new_n623), .B2(new_n285), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n502), .A2(new_n615), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n610), .A2(new_n613), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n614), .B(new_n626), .C1(new_n627), .C2(G169), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n610), .A2(G190), .A3(new_n613), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n501), .A2(new_n301), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n616), .B(new_n630), .C1(new_n623), .C2(new_n285), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n629), .B(new_n631), .C1(new_n627), .C2(new_n336), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n604), .A2(new_n607), .A3(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n442), .A2(new_n517), .A3(new_n567), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n436), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n331), .A2(new_n333), .ZN(new_n637));
  INV_X1    g0437(.A(new_n439), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n422), .B1(new_n638), .B2(new_n437), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n411), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n407), .ZN(new_n641));
  XOR2_X1   g0441(.A(new_n641), .B(KEYINPUT91), .Z(new_n642));
  NAND2_X1  g0442(.A1(new_n341), .A2(new_n342), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n637), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT92), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT92), .B1(new_n368), .B2(new_n370), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n636), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n613), .B(KEYINPUT88), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n610), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n651), .B2(new_n326), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n614), .A2(new_n626), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(G169), .B1(new_n650), .B2(new_n610), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n649), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n629), .A2(new_n631), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(G200), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n654), .A2(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n659), .B(new_n515), .C1(new_n509), .C2(new_n604), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n563), .A2(new_n566), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n535), .A2(KEYINPUT82), .A3(new_n551), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n554), .B1(new_n553), .B2(new_n557), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n628), .A2(new_n632), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n552), .A2(new_n666), .A3(new_n558), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT26), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n654), .A2(new_n656), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n548), .B2(new_n550), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n548), .A2(new_n670), .A3(new_n550), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n565), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n659), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n668), .A2(new_n669), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n442), .B1(new_n665), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n648), .A2(new_n678), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n497), .A2(new_n207), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT93), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n604), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n511), .A2(new_n686), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n517), .A2(KEYINPUT94), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT94), .B1(new_n517), .B2(new_n690), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n513), .A2(new_n686), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n517), .A2(new_n690), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT94), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n509), .A2(new_n686), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n517), .A2(KEYINPUT94), .A3(new_n690), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n686), .A2(new_n579), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n604), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n604), .B2(new_n607), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n696), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n210), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR4_X1   g0513(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G1), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n218), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n713), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n517), .A2(new_n567), .A3(new_n634), .A4(new_n687), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n599), .A2(new_n600), .A3(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n610), .A2(new_n613), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n462), .A2(new_n469), .A3(new_n470), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT95), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT95), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n506), .A2(new_n724), .A3(new_n610), .A4(new_n613), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n720), .A2(new_n723), .A3(new_n547), .A4(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT96), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AND4_X1   g0529(.A1(G179), .A2(new_n547), .A3(new_n600), .A4(new_n599), .ZN(new_n730));
  INV_X1    g0530(.A(new_n728), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n723), .A3(new_n725), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n651), .B(KEYINPUT97), .Z(new_n734));
  AND4_X1   g0534(.A1(new_n309), .A2(new_n601), .A3(new_n559), .A4(new_n471), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n729), .A2(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n687), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n719), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n664), .A2(KEYINPUT98), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT98), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n567), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n657), .A2(new_n658), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n669), .A2(new_n515), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n604), .A2(new_n509), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n565), .ZN(new_n753));
  INV_X1    g0553(.A(new_n673), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(new_n671), .ZN(new_n755));
  INV_X1    g0555(.A(new_n656), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n614), .B(new_n626), .C1(new_n655), .C2(new_n649), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n748), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT26), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n552), .A2(new_n666), .A3(new_n558), .A4(new_n675), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n759), .A2(new_n669), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n686), .B1(new_n752), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT29), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n687), .B1(new_n677), .B2(new_n665), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT29), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n744), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n718), .B1(new_n767), .B2(G1), .ZN(G364));
  AND2_X1   g0568(.A1(new_n207), .A2(G13), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n206), .B1(new_n769), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n712), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n708), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n706), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G330), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n213), .B1(G20), .B2(new_n326), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n207), .A2(new_n334), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n336), .A2(G179), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G303), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n278), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n309), .A2(G200), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n207), .A2(G190), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G179), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G322), .A2(new_n789), .B1(new_n793), .B2(G329), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n790), .A2(new_n784), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n790), .A2(new_n788), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n794), .B1(new_n795), .B2(new_n796), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n207), .B1(new_n791), .B2(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n787), .B(new_n800), .C1(G294), .C2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT100), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT100), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n805), .A2(G190), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G326), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n805), .A2(new_n334), .A3(new_n806), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI211_X1 g0611(.A(new_n803), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT101), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n789), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n815), .A2(new_n260), .B1(new_n799), .B2(new_n354), .ZN(new_n816));
  INV_X1    g0616(.A(new_n796), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(G107), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n792), .A2(new_n264), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT32), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n274), .B1(new_n785), .B2(new_n301), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G97), .B2(new_n802), .ZN(new_n822));
  INV_X1    g0622(.A(new_n810), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G50), .A2(new_n808), .B1(new_n823), .B2(G68), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n818), .A2(new_n820), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n812), .B2(new_n813), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n782), .B1(new_n814), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n772), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n244), .A2(G45), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT99), .ZN(new_n830));
  INV_X1    g0630(.A(new_n252), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n711), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n830), .B(new_n832), .C1(G45), .C2(new_n716), .ZN(new_n833));
  INV_X1    g0633(.A(G355), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n210), .A2(new_n274), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(G116), .B2(new_n210), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n779), .A2(new_n782), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n828), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n827), .A2(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n774), .A2(new_n776), .B1(new_n781), .B2(new_n839), .ZN(G396));
  INV_X1    g0640(.A(new_n782), .ZN(new_n841));
  INV_X1    g0641(.A(G294), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n815), .A2(new_n842), .B1(new_n792), .B2(new_n797), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n799), .A2(new_n573), .B1(new_n301), .B2(new_n796), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n278), .B1(new_n801), .B2(new_n619), .C1(new_n424), .C2(new_n785), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n795), .B2(new_n810), .C1(new_n786), .C2(new_n807), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT102), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G143), .A2(new_n789), .B1(new_n798), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n850), .B2(new_n807), .C1(new_n851), .C2(new_n810), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n831), .B1(new_n260), .B2(new_n801), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n796), .A2(new_n261), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n785), .A2(new_n202), .B1(new_n792), .B2(new_n857), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n852), .A2(new_n853), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n854), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n841), .B1(new_n848), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n782), .A2(new_n777), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n828), .B(new_n862), .C1(new_n354), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n686), .A2(new_n421), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n639), .B1(new_n433), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n440), .A2(new_n686), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n864), .B1(new_n778), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n868), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n764), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n687), .B(new_n868), .C1(new_n677), .C2(new_n665), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n744), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT103), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n744), .A2(new_n871), .A3(new_n872), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n828), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(KEYINPUT103), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n869), .B1(new_n876), .B2(new_n877), .ZN(G384));
  OAI211_X1 g0678(.A(G116), .B(new_n214), .C1(new_n524), .C2(KEYINPUT35), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(KEYINPUT35), .B2(new_n524), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT36), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n218), .B(G77), .C1(new_n260), .C2(new_n261), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n202), .A2(G68), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n206), .B(G13), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n412), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n686), .A2(new_n406), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n407), .A2(KEYINPUT104), .A3(new_n411), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n888), .ZN(new_n891));
  AOI221_X4 g0691(.A(new_n886), .B1(new_n409), .B2(new_n410), .C1(new_n393), .C2(new_n406), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT104), .B1(new_n407), .B2(new_n411), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n867), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n872), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n253), .A2(new_n254), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT73), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n255), .A3(new_n256), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n271), .B1(new_n901), .B2(G68), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n474), .B1(new_n902), .B2(KEYINPUT16), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n259), .A2(new_n268), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n270), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n294), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n339), .B1(new_n906), .B2(new_n684), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n328), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n684), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n296), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n330), .A2(new_n911), .A3(new_n912), .A4(new_n339), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n906), .A2(new_n684), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n343), .A2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT38), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n914), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n897), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n637), .B2(new_n910), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n407), .A2(new_n686), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT39), .B1(new_n917), .B2(new_n918), .ZN(new_n923));
  INV_X1    g0723(.A(new_n911), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n343), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n330), .A2(new_n911), .A3(new_n339), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n913), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT38), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT38), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n922), .B1(new_n923), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n920), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n763), .A2(new_n442), .A3(new_n766), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n648), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n719), .A2(new_n738), .A3(new_n741), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n890), .A2(new_n894), .A3(new_n868), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n917), .B2(new_n918), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n931), .A2(new_n933), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n943), .A2(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n442), .A2(new_n742), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n707), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n939), .A2(new_n950), .B1(new_n206), .B2(new_n769), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n939), .A2(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n885), .B1(new_n951), .B2(new_n952), .ZN(G367));
  NOR2_X1   g0753(.A1(new_n755), .A2(new_n687), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n745), .A2(new_n747), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n686), .A2(new_n753), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n702), .A3(new_n689), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n957), .A2(new_n513), .B1(new_n662), .B2(new_n663), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n959), .A2(KEYINPUT42), .B1(new_n960), .B2(new_n687), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT42), .B2(new_n959), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n687), .A2(new_n631), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n659), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n669), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(KEYINPUT105), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(KEYINPUT105), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n962), .A2(new_n966), .B1(KEYINPUT107), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(KEYINPUT107), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n709), .A2(new_n957), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n971), .B(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n712), .B(KEYINPUT41), .Z(new_n976));
  INV_X1    g0776(.A(new_n708), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n691), .A2(new_n692), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n977), .B1(new_n978), .B2(new_n700), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n702), .A2(new_n708), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n688), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n977), .A3(new_n700), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(new_n709), .A3(new_n689), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n767), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT110), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n693), .A2(new_n695), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT109), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n989), .A3(new_n957), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n989), .B1(new_n988), .B2(new_n957), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT109), .B1(new_n696), .B2(new_n958), .ZN(new_n994));
  INV_X1    g0794(.A(new_n987), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n990), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n696), .A2(new_n958), .A3(KEYINPUT45), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n988), .B2(new_n957), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n993), .A2(new_n996), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n979), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n993), .A2(new_n996), .A3(new_n709), .A4(new_n1000), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n986), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n976), .B1(new_n1004), .B2(new_n767), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n975), .B1(new_n1005), .B2(new_n771), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n832), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n837), .B1(new_n210), .B2(new_n415), .C1(new_n1007), .C2(new_n236), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n772), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT111), .Z(new_n1010));
  OAI221_X1 g0810(.A(new_n274), .B1(new_n261), .B2(new_n801), .C1(new_n799), .C2(new_n202), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n785), .A2(new_n260), .B1(new_n796), .B2(new_n354), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n815), .A2(new_n851), .B1(new_n792), .B2(new_n850), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n264), .B2(new_n810), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G143), .B2(new_n808), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT112), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n785), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(G116), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT46), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n252), .C1(new_n424), .C2(new_n801), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n815), .A2(new_n786), .B1(new_n799), .B2(new_n795), .ZN(new_n1022));
  INV_X1    g0822(.A(G317), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n796), .A2(new_n619), .B1(new_n792), .B2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G294), .A2(new_n823), .B1(new_n808), .B2(G311), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1017), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(KEYINPUT47), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n782), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(KEYINPUT47), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1010), .B1(new_n780), .B2(new_n965), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1006), .A2(new_n1031), .ZN(G387));
  AOI22_X1  g0832(.A1(G317), .A2(new_n789), .B1(new_n798), .B2(G303), .ZN(new_n1033));
  INV_X1    g0833(.A(G322), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1033), .B1(new_n797), .B2(new_n810), .C1(new_n1034), .C2(new_n807), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT116), .Z(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT48), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(KEYINPUT48), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1018), .A2(G294), .B1(new_n802), .B2(G283), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT49), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n796), .A2(new_n573), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n831), .B(new_n1044), .C1(G326), .C2(new_n793), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n808), .A2(G159), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT115), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n823), .A2(new_n288), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1018), .A2(G77), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n261), .B2(new_n799), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G50), .B2(new_n789), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n796), .A2(new_n619), .B1(new_n792), .B2(new_n851), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n801), .A2(new_n415), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1053), .A2(new_n252), .A3(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n841), .B1(new_n1046), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n287), .A2(G50), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1059));
  XNOR2_X1  g0859(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n714), .B(new_n315), .C1(new_n261), .C2(new_n354), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT113), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n832), .B1(new_n1060), .B2(new_n1062), .C1(new_n233), .C2(new_n315), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(G107), .B2(new_n210), .C1(new_n714), .C2(new_n835), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n828), .B(new_n1057), .C1(new_n837), .C2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT117), .Z(new_n1066));
  NAND3_X1  g0866(.A1(new_n978), .A2(new_n700), .A3(new_n779), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n981), .A2(new_n983), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1066), .A2(new_n1067), .B1(new_n771), .B2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n984), .A2(new_n712), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n767), .B2(new_n1069), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(G393));
  NAND3_X1  g0873(.A1(new_n1002), .A2(new_n771), .A3(new_n1003), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n241), .A2(new_n1007), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n837), .B1(new_n619), .B2(new_n210), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n772), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n808), .A2(G317), .B1(G311), .B2(new_n789), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n810), .A2(new_n786), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G322), .A2(new_n793), .B1(new_n798), .B2(G294), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n795), .B2(new_n785), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n278), .B1(new_n801), .B2(new_n573), .C1(new_n424), .C2(new_n796), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT118), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G87), .A2(new_n817), .B1(new_n793), .B2(G143), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n261), .B2(new_n785), .C1(new_n287), .C2(new_n799), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n801), .A2(new_n354), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1087), .A2(new_n252), .A3(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n264), .A2(new_n815), .B1(new_n807), .B2(new_n851), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(new_n202), .C2(new_n810), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1084), .A2(KEYINPUT118), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1085), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1077), .B1(new_n1094), .B2(new_n782), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n958), .B2(new_n780), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1074), .A2(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1004), .A2(new_n712), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n984), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1097), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  OAI211_X1 g0902(.A(new_n923), .B(new_n934), .C1(new_n921), .C2(new_n897), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n866), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n867), .B1(new_n762), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n945), .B(new_n922), .C1(new_n1105), .C2(new_n895), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n895), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1107), .A2(G330), .A3(new_n742), .A4(new_n868), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1103), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n948), .A2(G330), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n648), .A2(new_n1112), .A3(new_n937), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT119), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n743), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n742), .A2(KEYINPUT119), .A3(G330), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n870), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1114), .B1(new_n1118), .B2(new_n1107), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n895), .B1(new_n743), .B2(new_n870), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1108), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n872), .A2(new_n896), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1113), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n712), .B1(new_n1111), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1108), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT120), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1103), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1128), .A2(new_n1124), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT120), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1125), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n923), .A2(new_n934), .A3(new_n777), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n793), .A2(G125), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1136), .B1(new_n799), .B2(new_n1137), .C1(new_n857), .C2(new_n815), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n785), .A2(new_n851), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT53), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n264), .B2(new_n801), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n274), .B1(new_n202), .B2(new_n796), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1138), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n807), .C1(new_n850), .C2(new_n810), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n815), .A2(new_n573), .B1(new_n796), .B2(new_n261), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n799), .A2(new_n619), .B1(new_n792), .B2(new_n842), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n278), .B1(new_n785), .B2(new_n301), .ZN(new_n1149));
  NOR4_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1088), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n424), .B2(new_n810), .C1(new_n795), .C2(new_n807), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n841), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n828), .B(new_n1152), .C1(new_n287), .C2(new_n863), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1135), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1111), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n770), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1134), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(G378));
  OR2_X1    g0958(.A1(new_n920), .A2(new_n935), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT38), .B1(new_n925), .B2(new_n928), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n942), .B(KEYINPUT40), .C1(new_n917), .C2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n742), .A2(new_n868), .A3(new_n894), .A4(new_n890), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n914), .A2(new_n916), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n930), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n1164), .B2(new_n933), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1161), .B(G330), .C1(new_n1165), .C2(KEYINPUT40), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  NAND2_X1  g0967(.A1(new_n910), .A2(new_n364), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n647), .A2(new_n436), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n647), .B2(new_n436), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1167), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1166), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n947), .B2(G330), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1159), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT123), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1166), .A2(new_n1177), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n947), .A2(G330), .A3(new_n1176), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n936), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n936), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT123), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n771), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n828), .B1(new_n202), .B2(new_n863), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n815), .A2(new_n424), .B1(new_n792), .B2(new_n795), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1050), .B1(new_n260), .B2(new_n796), .C1(new_n261), .C2(new_n801), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n615), .C2(new_n798), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G97), .A2(new_n823), .B1(new_n808), .B2(G116), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n314), .A3(new_n252), .A4(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G50), .B1(new_n249), .B2(new_n314), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n831), .B2(G41), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n810), .A2(new_n857), .B1(new_n799), .B2(new_n850), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT121), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1137), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1018), .A2(new_n1203), .B1(new_n789), .B2(G128), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT122), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n808), .A2(G125), .B1(G150), .B2(new_n802), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT59), .Z(new_n1208));
  OAI211_X1 g1008(.A(new_n249), .B(new_n314), .C1(new_n796), .C2(new_n264), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G124), .B2(new_n793), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1196), .B(new_n1200), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1189), .B1(new_n841), .B2(new_n1211), .C1(new_n1176), .C2(new_n778), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1188), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT124), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1188), .A2(KEYINPUT124), .A3(new_n1212), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1113), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1129), .B1(new_n1111), .B2(new_n1124), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1131), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1221), .A2(KEYINPUT123), .A3(new_n1159), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1186), .A2(KEYINPUT123), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1184), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1113), .B1(new_n1133), .B2(new_n1131), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1184), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1186), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n712), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1215), .B(new_n1216), .C1(new_n1225), .C2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n895), .A2(new_n777), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n815), .A2(new_n795), .B1(new_n792), .B2(new_n786), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n799), .A2(new_n424), .B1(new_n619), .B2(new_n785), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n278), .B1(new_n796), .B2(new_n354), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1054), .A4(new_n1235), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n573), .B2(new_n810), .C1(new_n842), .C2(new_n807), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n815), .A2(new_n850), .B1(new_n796), .B2(new_n260), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n252), .B(new_n1238), .C1(G50), .C2(new_n802), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n785), .A2(new_n264), .B1(new_n792), .B2(new_n1145), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G150), .B2(new_n798), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G132), .A2(new_n808), .B1(new_n823), .B2(new_n1203), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n841), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n828), .B(new_n1244), .C1(new_n261), .C2(new_n863), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1231), .A2(new_n771), .B1(new_n1232), .B2(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1124), .A2(new_n976), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1231), .A2(new_n1217), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1247), .B2(new_n1248), .ZN(G381));
  OR2_X1    g1049(.A1(G375), .A2(G378), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1101), .A2(new_n1006), .A3(new_n1031), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  INV_X1    g1052(.A(G384), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OR4_X1    g1054(.A1(G381), .A2(new_n1250), .A3(new_n1251), .A4(new_n1254), .ZN(G407));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  INV_X1    g1056(.A(G396), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1252), .A2(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1101), .A2(new_n1006), .A3(new_n1031), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1101), .B1(new_n1006), .B2(new_n1031), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1259), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G387), .A2(G390), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1251), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT126), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1266), .B(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1226), .A2(new_n1269), .A3(new_n976), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n771), .B1(new_n1227), .B2(new_n1186), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1212), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1157), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(G375), .B2(new_n1157), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n685), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1248), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT60), .B1(new_n1231), .B2(new_n1217), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1124), .A2(new_n713), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G384), .B(new_n1246), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1246), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1253), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1276), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT57), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1226), .B2(new_n1269), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1292), .B(new_n712), .C1(new_n1226), .C2(new_n1228), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1293), .A2(G378), .A3(new_n1216), .A4(new_n1215), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1290), .B1(new_n1294), .B2(new_n1273), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1276), .A2(KEYINPUT125), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1282), .A2(new_n1285), .A3(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1290), .A2(G2897), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1297), .B(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1288), .B(new_n1289), .C1(new_n1295), .C2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1275), .B1(new_n1295), .B2(new_n1287), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1268), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1287), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1299), .B1(new_n1276), .B2(new_n1274), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1262), .A2(new_n1265), .A3(new_n1289), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1274), .A2(new_n1276), .A3(new_n1287), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1308), .B2(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1302), .A2(new_n1310), .ZN(G405));
  NAND2_X1  g1111(.A1(G375), .A2(G378), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT127), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1286), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1250), .A2(new_n1312), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1266), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1286), .A2(new_n1313), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1266), .A2(new_n1250), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1318), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(G402));
endmodule


