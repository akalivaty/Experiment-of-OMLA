//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(G137), .A3(new_n463), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  AOI21_X1  g051(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI211_X1 g060(.A(G138), .B(new_n463), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n468), .A2(new_n488), .A3(G138), .A4(new_n463), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n463), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT68), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n477), .A2(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n490), .A2(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n512), .A2(G50), .A3(G543), .A4(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n512), .A2(new_n518), .A3(G88), .A4(new_n514), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n509), .A2(new_n515), .A3(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  AND3_X1   g096(.A1(new_n512), .A2(G543), .A3(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n513), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n514), .B1(new_n504), .B2(new_n505), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n518), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n523), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n522), .A2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n506), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n528), .A2(G90), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT70), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n537), .A2(new_n545), .A3(new_n542), .A4(new_n541), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n506), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n513), .B1(new_n550), .B2(KEYINPUT71), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n551), .B1(KEYINPUT71), .B2(new_n550), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT72), .B(G43), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n522), .A2(new_n553), .B1(new_n528), .B2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G860), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND3_X1  g137(.A1(new_n512), .A2(new_n514), .A3(new_n518), .ZN(new_n563));
  INV_X1    g138(.A(G91), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT74), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n528), .A2(new_n566), .A3(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n506), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n565), .A2(new_n567), .B1(G651), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n512), .A2(G53), .A3(G543), .A4(new_n514), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND2_X1  g150(.A1(new_n522), .A2(G49), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n522), .A2(new_n578), .A3(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n528), .A2(G87), .ZN(new_n581));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n513), .B1(new_n506), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(G288));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n516), .B2(new_n517), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n512), .A2(new_n518), .A3(G86), .A4(new_n514), .ZN(new_n590));
  AND2_X1   g165(.A1(G48), .A2(G543), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n512), .A2(new_n514), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n522), .A2(G47), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n528), .A2(G85), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n594), .B(new_n595), .C1(new_n513), .C2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(new_n528), .A2(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n506), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n522), .A2(G54), .B1(G651), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G868), .B2(G171), .ZN(G321));
  XOR2_X1   g182(.A(G321), .B(KEYINPUT76), .Z(G284));
  AOI21_X1  g183(.A(G868), .B1(G299), .B2(KEYINPUT78), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(KEYINPUT78), .B2(G299), .ZN(new_n610));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT77), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n612), .ZN(G297));
  NAND2_X1  g188(.A1(new_n610), .A2(new_n612), .ZN(G280));
  INV_X1    g189(.A(new_n605), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n555), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n605), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n468), .A2(new_n473), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT79), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n482), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n477), .A2(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n463), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  OAI211_X1 g209(.A(new_n628), .B(new_n634), .C1(new_n626), .C2(new_n625), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT83), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2427), .B(G2430), .Z(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n638), .A2(new_n639), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  OR2_X1    g226(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(new_n626), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT18), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n657), .A2(new_n658), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2096), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n662), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n670), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n670), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT85), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT86), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  NAND2_X1  g263(.A1(new_n482), .A2(G139), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT25), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n468), .A2(G127), .ZN(new_n692));
  NAND2_X1  g267(.A1(G115), .A2(G2104), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n689), .B(new_n691), .C1(new_n694), .C2(new_n463), .ZN(new_n695));
  MUX2_X1   g270(.A(G33), .B(new_n695), .S(G29), .Z(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(G2072), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT93), .Z(new_n698));
  XOR2_X1   g273(.A(KEYINPUT89), .B(G16), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G19), .ZN(new_n701));
  INV_X1    g276(.A(new_n555), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1341), .Z(new_n704));
  NOR2_X1   g279(.A1(G29), .A2(G35), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G162), .B2(G29), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n698), .B(new_n704), .C1(G2090), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n615), .A2(G16), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G4), .B2(G16), .ZN(new_n711));
  INV_X1    g286(.A(G1348), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G27), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G164), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2078), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n711), .A2(new_n712), .ZN(new_n718));
  NOR4_X1   g293(.A1(new_n709), .A2(new_n713), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n708), .A2(G2090), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT99), .ZN(new_n721));
  NOR2_X1   g296(.A1(G5), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G171), .B2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1961), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n699), .A2(G20), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT23), .Z(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G299), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G1956), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G21), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(G16), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G286), .B2(G16), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT95), .B(G1966), .Z(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n477), .A2(G129), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT94), .Z(new_n737));
  AND2_X1   g312(.A1(new_n473), .A2(G105), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT26), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n738), .B(new_n740), .C1(G141), .C2(new_n482), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n714), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n714), .B2(G32), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n735), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n714), .A2(G26), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT28), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n482), .A2(G140), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n477), .A2(G128), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n463), .A2(G116), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT92), .Z(new_n756));
  AOI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n696), .A2(G2072), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n633), .A2(new_n714), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n714), .B1(new_n763), .B2(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n763), .B2(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G160), .B2(G29), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n760), .B(new_n762), .C1(G2084), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n733), .A2(new_n734), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(G2084), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G28), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT97), .Z(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(new_n714), .C1(new_n771), .C2(G28), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n748), .A2(new_n759), .A3(new_n767), .A4(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n719), .A2(new_n721), .A3(new_n730), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n482), .A2(G131), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n477), .A2(G119), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n463), .A2(G107), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT87), .Z(new_n783));
  MUX2_X1   g358(.A(G25), .B(new_n783), .S(G29), .Z(new_n784));
  XOR2_X1   g359(.A(KEYINPUT35), .B(G1991), .Z(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n786), .A2(KEYINPUT88), .A3(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n700), .A2(G24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G290), .B2(new_n699), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT90), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1986), .Z(new_n792));
  AOI21_X1  g367(.A(KEYINPUT88), .B1(new_n786), .B2(new_n787), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n788), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT91), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT32), .B(G1981), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G23), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(G16), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G288), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n700), .A2(G22), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n700), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1971), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n796), .B2(new_n797), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n798), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT34), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n794), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT36), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n794), .A2(new_n810), .A3(new_n814), .A4(new_n811), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n777), .B1(new_n813), .B2(new_n815), .ZN(G311));
  XNOR2_X1  g391(.A(G311), .B(KEYINPUT100), .ZN(G150));
  AOI22_X1  g392(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(new_n513), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n512), .A2(G55), .A3(G543), .A4(new_n514), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n563), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n528), .A2(G93), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT101), .B1(new_n825), .B2(new_n820), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n819), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(KEYINPUT102), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(new_n819), .C1(new_n824), .C2(new_n826), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n831), .A2(new_n702), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n702), .B1(new_n831), .B2(new_n833), .ZN(new_n835));
  OR3_X1    g410(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT38), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n605), .A2(new_n616), .ZN(new_n837));
  OAI21_X1  g412(.A(KEYINPUT38), .B1(new_n834), .B2(new_n835), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n830), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n556), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n839), .A2(new_n840), .A3(new_n830), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n829), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT103), .ZN(G145));
  XOR2_X1   g420(.A(new_n624), .B(new_n782), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n482), .A2(G142), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT105), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n477), .A2(G130), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n463), .A2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n846), .B(new_n852), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n756), .B(new_n742), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(G164), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(G164), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n695), .B(KEYINPUT104), .Z(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n855), .B2(new_n856), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n853), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G160), .B(new_n633), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n859), .A2(new_n861), .A3(KEYINPUT106), .A4(new_n853), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n859), .A2(new_n853), .A3(new_n861), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  INV_X1    g446(.A(new_n867), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n864), .B1(new_n872), .B2(new_n862), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  OAI22_X1  g450(.A1(new_n834), .A2(new_n835), .B1(G559), .B2(new_n605), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n831), .A2(new_n833), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n555), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n831), .A2(new_n702), .A3(new_n833), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n620), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n600), .A2(new_n573), .A3(new_n571), .A4(new_n604), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n600), .A2(new_n604), .B1(new_n571), .B2(new_n573), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n876), .A2(new_n880), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n883), .A2(new_n884), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n876), .B2(new_n880), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n889), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G288), .B(G305), .ZN(new_n898));
  XNOR2_X1  g473(.A(G290), .B(G166), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n898), .B(new_n899), .Z(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n898), .B(new_n899), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n618), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n827), .A2(new_n618), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n904), .A2(KEYINPUT107), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT107), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(G295));
  OR2_X1    g483(.A1(new_n904), .A2(new_n905), .ZN(G331));
  AOI21_X1  g484(.A(G286), .B1(new_n544), .B2(new_n546), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n544), .A2(G286), .A3(new_n546), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n834), .B2(new_n835), .ZN(new_n914));
  INV_X1    g489(.A(new_n912), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n878), .A2(new_n916), .A3(new_n879), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n888), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n917), .A3(new_n891), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n900), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n871), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n914), .A2(new_n917), .A3(new_n891), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n888), .B1(new_n914), .B2(new_n917), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n902), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n922), .A2(new_n871), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n920), .A2(new_n921), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT108), .B1(new_n930), .B2(new_n902), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  AOI211_X1 g507(.A(new_n932), .B(new_n900), .C1(new_n920), .C2(new_n921), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n928), .B1(new_n934), .B2(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n926), .A2(new_n922), .A3(new_n938), .A4(new_n871), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT44), .ZN(new_n940));
  AOI211_X1 g515(.A(KEYINPUT109), .B(new_n940), .C1(KEYINPUT43), .C2(new_n934), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(new_n940), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n937), .B1(new_n941), .B2(new_n945), .ZN(G397));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n490), .B2(new_n501), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT110), .B(G40), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n471), .A2(new_n475), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT111), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n756), .B(new_n758), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n743), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT126), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n952), .A2(G1996), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT46), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT47), .Z(new_n962));
  INV_X1    g537(.A(G1996), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n955), .B1(new_n963), .B2(new_n743), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n964), .A2(new_n953), .B1(new_n743), .B2(new_n959), .ZN(new_n965));
  INV_X1    g540(.A(new_n785), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n782), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n953), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n952), .A2(G1986), .A3(G290), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT48), .Z(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n756), .A2(G2067), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n783), .A2(new_n966), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n954), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n962), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n487), .A2(new_n489), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n493), .A2(new_n498), .B1(new_n477), .B2(G126), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n951), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI211_X1 g557(.A(KEYINPUT50), .B(G1384), .C1(new_n978), .C2(new_n979), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n728), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n948), .A2(new_n949), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT56), .B(G2072), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n985), .A2(new_n951), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(G299), .A2(KEYINPUT57), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n571), .A2(new_n990), .A3(new_n573), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n984), .A2(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n984), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n993), .A2(new_n615), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n712), .B1(new_n982), .B2(new_n983), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n951), .A2(new_n980), .A3(new_n758), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n995), .A2(KEYINPUT121), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT121), .B1(new_n995), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n992), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT60), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT60), .B1(new_n997), .B2(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n615), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT60), .B(new_n605), .C1(new_n997), .C2(new_n998), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n985), .A2(new_n963), .A3(new_n951), .A4(new_n986), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n951), .A2(new_n980), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT58), .B(G1341), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n702), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT59), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1013), .A3(new_n702), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT61), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n984), .A2(new_n988), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n989), .A2(new_n991), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1012), .A2(new_n1014), .B1(new_n1018), .B2(new_n993), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n993), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT61), .B1(new_n992), .B2(KEYINPUT122), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1000), .B1(new_n1005), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n985), .A2(new_n951), .A3(new_n986), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n734), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n948), .A2(KEYINPUT50), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n980), .A2(new_n981), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n951), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(G2084), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(G8), .A3(G286), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT123), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(G8), .C1(new_n1032), .C2(G286), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT124), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(KEYINPUT51), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n982), .A2(new_n983), .ZN(new_n1039));
  INV_X1    g614(.A(G2084), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1039), .A2(new_n1040), .B1(new_n1027), .B2(new_n734), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1041), .B2(G168), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT124), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT124), .B1(new_n1042), .B2(new_n1034), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1033), .B(new_n1037), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G305), .A2(G1981), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT116), .B(G1981), .Z(new_n1050));
  NAND4_X1  g625(.A1(new_n589), .A2(new_n590), .A3(new_n592), .A4(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1051), .A2(KEYINPUT117), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(KEYINPUT117), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1048), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n590), .A2(new_n1050), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n592), .A4(new_n589), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1051), .A2(KEYINPUT117), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1059), .A2(new_n1060), .B1(G1981), .B2(G305), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1054), .A2(KEYINPUT118), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1056), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT49), .B1(new_n1054), .B2(KEYINPUT118), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1048), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1038), .B1(new_n951), .B2(new_n980), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  INV_X1    g646(.A(G288), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT115), .B(G1976), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1069), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT112), .B(G1971), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1027), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(G2090), .B2(new_n1031), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(G303), .B2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(G303), .A2(G8), .A3(new_n1084), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1087), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1089), .A2(new_n1085), .A3(KEYINPUT114), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1082), .A2(G8), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G2090), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1039), .A2(new_n1093), .B1(new_n1027), .B2(new_n1080), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1094), .A2(new_n1038), .B1(new_n1089), .B2(new_n1085), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1070), .A2(new_n1079), .A3(new_n1092), .A4(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(G171), .B(KEYINPUT54), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1039), .A2(G1961), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1027), .B2(G2078), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(G2078), .ZN(new_n1101));
  AND3_X1   g676(.A1(G160), .A2(G40), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n985), .A2(new_n1102), .A3(new_n986), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .A4(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n985), .A2(new_n951), .A3(new_n986), .A4(new_n1101), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1098), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1104), .B1(new_n1106), .B2(new_n1097), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1096), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1026), .A2(new_n1047), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1094), .A2(new_n1038), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1070), .A2(new_n1079), .A3(new_n1110), .A4(new_n1091), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1112));
  NOR2_X1   g687(.A1(G288), .A2(G1976), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1070), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1069), .B(KEYINPUT120), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1111), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1041), .A2(new_n1038), .A3(G286), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1096), .B2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1070), .A2(new_n1079), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1095), .A2(new_n1092), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT63), .A4(new_n1118), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1116), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1109), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1109), .B2(new_n1124), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1047), .A2(KEYINPUT62), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(new_n1044), .A3(new_n1043), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n1033), .A4(new_n1037), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1096), .A2(G301), .A3(new_n1106), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1128), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1126), .A2(new_n1127), .A3(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(G290), .B(G1986), .Z(new_n1136));
  OAI21_X1  g711(.A(new_n969), .B1(new_n952), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n977), .B1(new_n1135), .B2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g713(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1140));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n1141));
  AND2_X1   g715(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1143));
  NOR3_X1   g717(.A1(G229), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g718(.A1(new_n935), .A2(new_n874), .A3(new_n1144), .ZN(G225));
  INV_X1    g719(.A(G225), .ZN(G308));
endmodule


