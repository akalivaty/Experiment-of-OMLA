//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT10), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G107), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n191), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n194), .B2(new_n192), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT82), .B(KEYINPUT3), .C1(new_n193), .C2(G107), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n197), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(G101), .B1(new_n194), .B2(new_n191), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G146), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT65), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n206), .B(G143), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n205), .A2(new_n211), .A3(new_n212), .A4(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n202), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT84), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI211_X1 g037(.A(KEYINPUT84), .B(new_n202), .C1(new_n220), .C2(new_n217), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n189), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT83), .A3(G101), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT4), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n200), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n205), .A2(new_n230), .A3(new_n211), .A4(new_n212), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n207), .A2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n214), .B1(new_n234), .B2(G143), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n229), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n204), .B1(new_n232), .B2(new_n233), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n243));
  OAI21_X1  g057(.A(G128), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n235), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n220), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n202), .A2(KEYINPUT85), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n200), .A2(new_n248), .A3(new_n201), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n247), .A2(KEYINPUT86), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT86), .B1(new_n247), .B2(new_n249), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT10), .B(new_n246), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n256), .A2(new_n253), .A3(KEYINPUT11), .A4(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n253), .A2(G134), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n253), .A2(G134), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n258), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n258), .B2(new_n262), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n225), .A2(new_n241), .A3(new_n252), .A4(new_n266), .ZN(new_n267));
  XOR2_X1   g081(.A(G110), .B(G140), .Z(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT81), .ZN(new_n269));
  INV_X1    g083(.A(G227), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n247), .A2(new_n249), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n245), .A3(new_n220), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n223), .B2(new_n224), .ZN(new_n275));
  INV_X1    g089(.A(new_n266), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n275), .A2(KEYINPUT12), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT12), .B1(new_n275), .B2(new_n276), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n267), .B(new_n272), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n225), .A2(new_n241), .A3(new_n252), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n276), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n272), .B1(new_n282), .B2(new_n267), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n187), .B(new_n188), .C1(new_n280), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(G469), .A2(G902), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n267), .B1(new_n277), .B2(new_n278), .ZN(new_n286));
  INV_X1    g100(.A(new_n272), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n282), .A2(new_n267), .A3(new_n272), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n284), .B(new_n285), .C1(new_n187), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G221), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT9), .B(G234), .Z(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n188), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G110), .B(G122), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT89), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G116), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G119), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT2), .B(G113), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n303), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G113), .B1(new_n308), .B2(new_n300), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n251), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n247), .A2(KEYINPUT86), .A3(new_n249), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(new_n303), .B(new_n304), .Z(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(new_n228), .B2(new_n200), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n298), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n316), .ZN(new_n318));
  INV_X1    g132(.A(new_n311), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n250), .B2(new_n251), .ZN(new_n320));
  INV_X1    g134(.A(new_n298), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n317), .A2(new_n322), .A3(KEYINPUT6), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT6), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n324), .B(new_n298), .C1(new_n314), .C2(new_n316), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n239), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n245), .A2(new_n220), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G224), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G953), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n323), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT7), .B1(new_n330), .B2(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n335), .B(KEYINPUT90), .Z(new_n336));
  XOR2_X1   g150(.A(new_n298), .B(KEYINPUT8), .Z(new_n337));
  AOI21_X1  g151(.A(new_n310), .B1(KEYINPUT5), .B2(new_n307), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n273), .A2(new_n305), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n311), .A2(new_n202), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n329), .A2(new_n334), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n336), .A2(new_n341), .A3(new_n322), .A4(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n333), .A2(new_n188), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G210), .B1(G237), .B2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n333), .A2(new_n188), .A3(new_n343), .A4(new_n345), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G214), .B1(G237), .B2(G902), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n350), .B(KEYINPUT87), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G116), .B(G122), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n190), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n301), .A2(KEYINPUT14), .A3(G122), .ZN(new_n356));
  INV_X1    g170(.A(new_n354), .ZN(new_n357));
  OAI211_X1 g171(.A(G107), .B(new_n356), .C1(new_n357), .C2(KEYINPUT14), .ZN(new_n358));
  XOR2_X1   g172(.A(G128), .B(G143), .Z(new_n359));
  INV_X1    g173(.A(KEYINPUT94), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G134), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n361), .A2(new_n362), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n355), .B(new_n358), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n362), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT93), .B(KEYINPUT13), .Z(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(G128), .A3(new_n204), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n368), .B(G134), .C1(new_n367), .C2(new_n359), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n354), .B(new_n190), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G953), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n293), .A2(G217), .A3(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n374), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n188), .ZN(new_n378));
  INV_X1    g192(.A(G478), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(KEYINPUT15), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n378), .B(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G475), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n193), .ZN(new_n385));
  XNOR2_X1  g199(.A(G125), .B(G140), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT19), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n386), .B1(KEYINPUT91), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT91), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT19), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n389), .A3(KEYINPUT19), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n203), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(KEYINPUT92), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n386), .B2(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G146), .ZN(new_n397));
  INV_X1    g211(.A(G237), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n373), .A3(G214), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(G143), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n263), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n393), .A2(KEYINPUT92), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n394), .A2(new_n397), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n400), .A2(new_n263), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT18), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n400), .B1(new_n406), .B2(new_n263), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n234), .A2(new_n386), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n209), .B2(new_n386), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n385), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n396), .B(new_n209), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n404), .A2(KEYINPUT17), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n412), .B(new_n413), .C1(new_n401), .C2(KEYINPUT17), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n414), .A2(new_n385), .A3(new_n410), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n383), .B(new_n188), .C1(new_n411), .C2(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n416), .A2(KEYINPUT20), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(KEYINPUT20), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n385), .B1(new_n414), .B2(new_n410), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n188), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n417), .A2(new_n418), .B1(G475), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n373), .A2(G952), .ZN(new_n422));
  NAND2_X1  g236(.A1(G234), .A2(G237), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT21), .B(G898), .Z(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(G902), .A3(G953), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n382), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n296), .A2(new_n353), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n299), .A2(G128), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT74), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(G119), .B2(new_n218), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT24), .B(G110), .Z(new_n433));
  OR3_X1    g247(.A1(new_n432), .A2(KEYINPUT77), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT77), .B1(new_n432), .B2(new_n433), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(KEYINPUT23), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT76), .B1(new_n218), .B2(G119), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n434), .B(new_n435), .C1(G110), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n408), .A3(new_n397), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n432), .A2(new_n433), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT75), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n412), .B1(G110), .B2(new_n438), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(G137), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n373), .A2(G221), .A3(G234), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n450), .B(KEYINPUT79), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n440), .B2(new_n445), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n188), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT25), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n450), .B(KEYINPUT79), .Z(new_n457));
  NAND2_X1  g271(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n446), .B2(new_n451), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT25), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n188), .ZN(new_n461));
  INV_X1    g275(.A(G217), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(G234), .B2(new_n188), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n456), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(G902), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n465), .B(KEYINPUT80), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(G101), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n398), .A2(new_n373), .A3(G210), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n315), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n266), .A2(new_n239), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n258), .A2(new_n262), .A3(new_n263), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n362), .A2(G137), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n259), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n245), .B2(new_n220), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n476), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n478), .A2(new_n480), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n246), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n231), .B(new_n238), .C1(new_n264), .C2(new_n265), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n315), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n475), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT28), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n473), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n485), .A2(new_n493), .A3(new_n486), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n485), .B2(new_n486), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n476), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n473), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n487), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT29), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n485), .A2(new_n315), .A3(new_n486), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n315), .B1(new_n485), .B2(new_n486), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n490), .B1(new_n502), .B2(new_n489), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n473), .A2(KEYINPUT29), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n188), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G472), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT72), .B(G472), .C1(new_n499), .C2(new_n505), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT32), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n497), .B1(new_n488), .B2(new_n491), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n487), .A2(new_n473), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n496), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT30), .B1(new_n477), .B2(new_n482), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n485), .A2(new_n493), .A3(new_n486), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n315), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT31), .B1(new_n520), .B2(new_n512), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT68), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n496), .B2(new_n513), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT68), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n517), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G472), .A2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n510), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n520), .A2(new_n512), .A3(new_n514), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n474), .B1(new_n500), .B2(new_n501), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n473), .B1(new_n532), .B2(new_n490), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n524), .A2(new_n525), .ZN(new_n535));
  AOI211_X1 g349(.A(KEYINPUT68), .B(new_n523), .C1(new_n496), .C2(new_n513), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT32), .A3(new_n528), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT71), .B(new_n510), .C1(new_n527), .C2(new_n529), .ZN(new_n541));
  AOI221_X4 g355(.A(KEYINPUT73), .B1(new_n508), .B2(new_n509), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n541), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n508), .A2(new_n509), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n429), .B(new_n469), .C1(new_n542), .C2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(G101), .ZN(G3));
  NAND2_X1  g362(.A1(new_n420), .A2(G475), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n416), .A2(KEYINPUT20), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n416), .A2(KEYINPUT20), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n376), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n372), .A2(new_n374), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT33), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n375), .A2(new_n556), .A3(new_n376), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n557), .A3(G478), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n377), .A2(new_n379), .A3(new_n188), .ZN(new_n559));
  NAND2_X1  g373(.A1(G478), .A2(G902), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n552), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT95), .Z(new_n563));
  AOI21_X1  g377(.A(new_n351), .B1(new_n347), .B2(new_n348), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n427), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n468), .A2(new_n294), .ZN(new_n567));
  INV_X1    g381(.A(G472), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n537), .B2(new_n188), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n528), .B2(new_n537), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n567), .A2(new_n291), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(new_n193), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n572), .B(new_n574), .ZN(G6));
  NAND2_X1  g389(.A1(new_n417), .A2(new_n418), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n549), .B(KEYINPUT97), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n565), .A2(new_n382), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n571), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G107), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT98), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n580), .B(new_n582), .ZN(G9));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n457), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n446), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n440), .A2(new_n457), .A3(new_n584), .A4(new_n445), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n466), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n464), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n429), .A2(new_n570), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n592), .B(KEYINPUT37), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G110), .ZN(G12));
  NAND2_X1  g408(.A1(new_n544), .A2(new_n545), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT73), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n544), .A2(new_n543), .A3(new_n545), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n296), .A2(new_n353), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n426), .A2(G900), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n424), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n382), .A2(new_n578), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n598), .A2(new_n599), .A3(new_n591), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G128), .ZN(G30));
  XNOR2_X1  g419(.A(new_n601), .B(KEYINPUT39), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n291), .A2(new_n295), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n349), .B(KEYINPUT38), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n552), .A2(new_n381), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n496), .A2(new_n487), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n473), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n502), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n188), .B1(new_n617), .B2(new_n473), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n544), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n591), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n609), .A2(new_n613), .A3(new_n622), .A4(new_n352), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT100), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G143), .ZN(G45));
  NOR2_X1   g439(.A1(new_n562), .A2(new_n602), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n598), .A2(new_n599), .A3(new_n591), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G146), .ZN(G48));
  AOI21_X1  g442(.A(new_n468), .B1(new_n596), .B2(new_n597), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n282), .A2(new_n267), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n287), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n279), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n188), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G469), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(KEYINPUT101), .A3(new_n284), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n633), .A2(new_n636), .A3(G469), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n294), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n629), .A2(new_n566), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT41), .B(G113), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G15));
  NAND4_X1  g455(.A1(new_n598), .A2(new_n469), .A3(new_n579), .A4(new_n638), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G116), .ZN(G18));
  AND2_X1   g457(.A1(new_n464), .A2(new_n590), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n596), .B2(new_n597), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n635), .A2(new_n637), .ZN(new_n646));
  INV_X1    g460(.A(new_n428), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n564), .A2(new_n646), .A3(new_n295), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G119), .ZN(G21));
  AOI21_X1  g464(.A(new_n524), .B1(new_n497), .B2(new_n503), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n529), .B1(new_n651), .B2(new_n516), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n569), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n646), .A2(new_n469), .A3(new_n295), .A4(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n611), .A2(KEYINPUT102), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n611), .A2(KEYINPUT102), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n564), .A3(new_n427), .A4(new_n656), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G122), .ZN(G24));
  NAND2_X1  g473(.A1(new_n653), .A2(new_n591), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n562), .B2(new_n602), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n552), .A2(new_n561), .A3(KEYINPUT104), .A4(new_n601), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n662), .A2(new_n564), .A3(new_n638), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G125), .ZN(G27));
  NAND3_X1  g482(.A1(new_n347), .A2(new_n352), .A3(new_n348), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n296), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n545), .A2(new_n530), .A3(new_n538), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n469), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AND4_X1   g487(.A1(KEYINPUT42), .A2(new_n670), .A3(new_n673), .A4(new_n666), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n598), .A2(new_n469), .A3(new_n666), .A4(new_n670), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n676));
  AOI21_X1  g490(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n263), .ZN(G33));
  NAND3_X1  g492(.A1(new_n629), .A2(new_n603), .A3(new_n670), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G134), .ZN(G36));
  INV_X1    g494(.A(new_n284), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n682), .B1(new_n290), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n187), .B1(new_n290), .B2(new_n683), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT106), .A4(KEYINPUT45), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n285), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n681), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(KEYINPUT46), .A3(new_n285), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n294), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n421), .A2(new_n561), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n421), .A2(new_n561), .A3(KEYINPUT43), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n570), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n591), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n669), .B1(new_n699), .B2(new_n700), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n692), .A2(new_n701), .A3(new_n606), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G137), .ZN(G39));
  AND3_X1   g518(.A1(new_n687), .A2(KEYINPUT46), .A3(new_n285), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT46), .B1(new_n687), .B2(new_n285), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n705), .A2(new_n706), .A3(new_n681), .ZN(new_n707));
  NOR2_X1   g521(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n708));
  NAND2_X1  g522(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  OAI22_X1  g524(.A1(new_n707), .A2(new_n294), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n692), .A2(new_n709), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n598), .A2(new_n469), .A3(new_n669), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n712), .A3(new_n713), .A4(new_n626), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G140), .ZN(G42));
  NAND2_X1  g529(.A1(new_n646), .A2(new_n295), .ZN(new_n716));
  INV_X1    g530(.A(new_n424), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n697), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n716), .A2(new_n669), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n673), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT48), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n718), .A2(new_n468), .A3(new_n569), .A4(new_n652), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n564), .A3(new_n638), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n721), .A2(new_n422), .A3(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n716), .A2(new_n468), .A3(new_n669), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n717), .A3(new_n621), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n552), .A3(new_n561), .ZN(new_n727));
  OR4_X1    g541(.A1(new_n352), .A2(new_n654), .A3(new_n610), .A4(new_n718), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n729));
  AOI21_X1  g543(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n669), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n711), .A2(new_n712), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n295), .B1(new_n635), .B2(new_n637), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n731), .B(new_n722), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n719), .A2(new_n662), .ZN(new_n735));
  OR3_X1    g549(.A1(new_n728), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n730), .A2(new_n734), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT51), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT51), .B1(new_n737), .B2(new_n738), .ZN(new_n740));
  OAI221_X1 g554(.A(new_n724), .B1(new_n563), .B2(new_n726), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n644), .A2(new_n291), .A3(new_n295), .A4(new_n601), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(KEYINPUT111), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n655), .A2(new_n564), .A3(new_n656), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(KEYINPUT111), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n620), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n604), .A2(new_n627), .A3(new_n667), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n645), .B(new_n599), .C1(new_n603), .C2(new_n626), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(KEYINPUT52), .A3(new_n667), .A4(new_n747), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n639), .A2(new_n649), .A3(new_n642), .A4(new_n658), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n562), .B1(new_n382), .B2(new_n552), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n571), .A2(new_n564), .A3(new_n427), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n547), .A2(new_n756), .A3(new_n592), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n754), .A2(new_n677), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n381), .A2(new_n602), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n591), .B(new_n760), .C1(new_n542), .C2(new_n546), .ZN(new_n761));
  INV_X1    g575(.A(new_n670), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n761), .A2(new_n578), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n660), .A2(new_n661), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT103), .B1(new_n653), .B2(new_n591), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n670), .B(new_n666), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n469), .B(new_n670), .C1(new_n542), .C2(new_n546), .ZN(new_n767));
  INV_X1    g581(.A(new_n603), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n759), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n578), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n645), .A2(new_n771), .A3(new_n670), .A4(new_n760), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n679), .A3(KEYINPUT110), .A4(new_n766), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n753), .A2(new_n758), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n753), .A2(new_n758), .A3(new_n774), .A4(KEYINPUT53), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n777), .A2(KEYINPUT54), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT54), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n742), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n782));
  INV_X1    g596(.A(new_n666), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n676), .B1(new_n767), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n674), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n469), .B(new_n638), .C1(new_n542), .C2(new_n546), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n788), .A2(new_n579), .B1(new_n645), .B2(new_n648), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n654), .A2(new_n657), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n788), .B2(new_n566), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n547), .A2(new_n592), .A3(new_n756), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n770), .B2(new_n773), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT53), .B1(new_n794), .B2(new_n753), .ZN(new_n795));
  INV_X1    g609(.A(new_n778), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n782), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n777), .A2(KEYINPUT54), .A3(new_n778), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(KEYINPUT112), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n741), .B1(new_n781), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(G952), .A2(G953), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT115), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n567), .A2(new_n352), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT108), .ZN(new_n804));
  INV_X1    g618(.A(new_n693), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n646), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n610), .B1(new_n807), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n646), .A2(new_n806), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n621), .A3(new_n811), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n800), .A2(new_n802), .B1(new_n809), .B2(new_n812), .ZN(G75));
  AOI21_X1  g627(.A(new_n188), .B1(new_n777), .B2(new_n778), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT56), .B1(new_n814), .B2(G210), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n323), .A2(new_n325), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(new_n332), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT55), .Z(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n815), .A2(new_n819), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n373), .A2(G952), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(G51));
  XOR2_X1   g637(.A(new_n285), .B(KEYINPUT57), .Z(new_n824));
  NAND3_X1  g638(.A1(new_n797), .A2(new_n798), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n632), .ZN(new_n826));
  INV_X1    g640(.A(new_n687), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n814), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n822), .B1(new_n826), .B2(new_n828), .ZN(G54));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n383), .ZN(new_n832));
  NAND3_X1  g646(.A1(KEYINPUT116), .A2(KEYINPUT58), .A3(G475), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n814), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n411), .A2(new_n415), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n834), .A2(new_n836), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n837), .A2(new_n838), .A3(new_n822), .ZN(G60));
  NAND2_X1  g653(.A1(new_n555), .A2(new_n557), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT117), .Z(new_n841));
  XOR2_X1   g655(.A(new_n560), .B(KEYINPUT59), .Z(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n797), .A2(new_n798), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n797), .A2(KEYINPUT118), .A3(new_n798), .A4(new_n843), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n822), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n842), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n781), .A2(new_n799), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n841), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n848), .A2(new_n851), .ZN(G63));
  INV_X1    g666(.A(new_n822), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n777), .A2(new_n778), .ZN(new_n854));
  NAND2_X1  g668(.A1(G217), .A2(G902), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT60), .Z(new_n856));
  NAND2_X1  g670(.A1(new_n586), .A2(new_n587), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT119), .Z(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n854), .A2(new_n856), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n853), .B(new_n859), .C1(new_n860), .C2(new_n459), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(G66));
  INV_X1    g677(.A(new_n425), .ZN(new_n864));
  OAI21_X1  g678(.A(G953), .B1(new_n864), .B2(new_n330), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n754), .A2(new_n757), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n816), .B1(G898), .B2(new_n373), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(G69));
  NAND2_X1  g683(.A1(new_n518), .A2(new_n519), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n391), .A2(new_n392), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n870), .B(new_n871), .Z(new_n872));
  NAND3_X1  g686(.A1(new_n751), .A2(new_n623), .A3(new_n667), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n755), .A2(new_n606), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT120), .B1(new_n767), .B2(new_n876), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n767), .A2(KEYINPUT120), .A3(new_n876), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n703), .A2(new_n714), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n872), .B1(new_n880), .B2(G953), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n692), .A2(new_n606), .A3(new_n745), .A4(new_n673), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n786), .A2(new_n714), .A3(new_n679), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n703), .A2(new_n751), .A3(new_n667), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT121), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n703), .A2(new_n751), .A3(new_n886), .A4(new_n667), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT122), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n883), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n890), .A2(new_n373), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n872), .ZN(new_n894));
  INV_X1    g708(.A(G900), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n373), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n881), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n373), .B1(G227), .B2(G900), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT123), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n897), .B(new_n899), .Z(G72));
  NAND3_X1  g714(.A1(new_n875), .A2(new_n866), .A3(new_n879), .ZN(new_n901));
  XOR2_X1   g715(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n902));
  NOR2_X1   g716(.A1(new_n568), .A2(new_n188), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n902), .B(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT125), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n901), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n616), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT126), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n907), .A2(new_n912), .A3(new_n616), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n890), .A2(new_n866), .A3(new_n892), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(new_n905), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n915), .B(new_n853), .C1(new_n917), .C2(new_n498), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n854), .A2(new_n498), .A3(new_n615), .A4(new_n905), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n498), .B1(new_n916), .B2(new_n905), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT127), .B1(new_n920), .B2(new_n822), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n914), .A2(new_n918), .A3(new_n919), .A4(new_n921), .ZN(G57));
endmodule


