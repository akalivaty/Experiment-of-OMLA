

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X2 U323 ( .A(G218GAT), .B(G162GAT), .Z(n429) );
  XNOR2_X1 U324 ( .A(n375), .B(n374), .ZN(n554) );
  XNOR2_X1 U325 ( .A(n398), .B(KEYINPUT64), .ZN(n399) );
  XNOR2_X1 U326 ( .A(n400), .B(n399), .ZN(n415) );
  XNOR2_X1 U327 ( .A(n373), .B(n412), .ZN(n374) );
  XNOR2_X1 U328 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U329 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n296) );
  XOR2_X1 U331 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n292) );
  XNOR2_X1 U332 ( .A(G43GAT), .B(G99GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n294) );
  XNOR2_X1 U334 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n293), .B(KEYINPUT80), .ZN(n313) );
  XNOR2_X1 U336 ( .A(n294), .B(n313), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U338 ( .A(G190GAT), .B(G134GAT), .Z(n364) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n405) );
  XOR2_X1 U340 ( .A(n364), .B(n405), .Z(n298) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U343 ( .A(n300), .B(n299), .Z(n306) );
  XOR2_X1 U344 ( .A(G113GAT), .B(G15GAT), .Z(n351) );
  XNOR2_X1 U345 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n301), .B(KEYINPUT19), .ZN(n302) );
  XOR2_X1 U347 ( .A(n302), .B(KEYINPUT18), .Z(n304) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G176GAT), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n340) );
  XNOR2_X1 U350 ( .A(n351), .B(n340), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n504) );
  XOR2_X1 U352 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n308) );
  XNOR2_X1 U353 ( .A(KEYINPUT89), .B(G57GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U355 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n310) );
  XNOR2_X1 U356 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U358 ( .A(n312), .B(n311), .Z(n318) );
  XOR2_X1 U359 ( .A(G85GAT), .B(n313), .Z(n315) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U362 ( .A(G29GAT), .B(n316), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U364 ( .A(G162GAT), .B(G120GAT), .Z(n320) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G134GAT), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U367 ( .A(n322), .B(n321), .Z(n330) );
  XOR2_X1 U368 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n324) );
  XNOR2_X1 U369 ( .A(KEYINPUT87), .B(G155GAT), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U371 ( .A(KEYINPUT2), .B(n325), .Z(n440) );
  XOR2_X1 U372 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n327) );
  XNOR2_X1 U373 ( .A(G141GAT), .B(G148GAT), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U375 ( .A(n440), .B(n328), .ZN(n329) );
  XNOR2_X1 U376 ( .A(n330), .B(n329), .ZN(n513) );
  XOR2_X1 U377 ( .A(G64GAT), .B(G190GAT), .Z(n332) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(G8GAT), .ZN(n331) );
  XNOR2_X1 U379 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U380 ( .A(G92GAT), .B(KEYINPUT93), .Z(n334) );
  XNOR2_X1 U381 ( .A(G218GAT), .B(KEYINPUT92), .ZN(n333) );
  XNOR2_X1 U382 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U383 ( .A(n336), .B(n335), .Z(n338) );
  NAND2_X1 U384 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U385 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U386 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U387 ( .A(KEYINPUT85), .B(G211GAT), .Z(n342) );
  XNOR2_X1 U388 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n341) );
  XNOR2_X1 U389 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U390 ( .A(G197GAT), .B(n343), .ZN(n441) );
  XNOR2_X1 U391 ( .A(n344), .B(n441), .ZN(n502) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n345) );
  XNOR2_X1 U393 ( .A(n345), .B(G29GAT), .ZN(n346) );
  XOR2_X1 U394 ( .A(n346), .B(KEYINPUT7), .Z(n348) );
  XNOR2_X1 U395 ( .A(G43GAT), .B(G50GAT), .ZN(n347) );
  XNOR2_X1 U396 ( .A(n348), .B(n347), .ZN(n373) );
  XOR2_X1 U397 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n350) );
  XNOR2_X1 U398 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n349) );
  XNOR2_X1 U399 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U400 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U401 ( .A(G141GAT), .B(G22GAT), .Z(n436) );
  XOR2_X1 U402 ( .A(n436), .B(KEYINPUT69), .Z(n354) );
  NAND2_X1 U403 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U405 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U406 ( .A(G1GAT), .B(G8GAT), .Z(n384) );
  XOR2_X1 U407 ( .A(n357), .B(n384), .Z(n359) );
  XNOR2_X1 U408 ( .A(G169GAT), .B(G197GAT), .ZN(n358) );
  XNOR2_X1 U409 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n373), .B(n360), .ZN(n569) );
  XNOR2_X1 U411 ( .A(KEYINPUT70), .B(n569), .ZN(n557) );
  INV_X1 U412 ( .A(KEYINPUT77), .ZN(n376) );
  XOR2_X1 U413 ( .A(KEYINPUT75), .B(KEYINPUT65), .Z(n362) );
  XNOR2_X1 U414 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U416 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n363) );
  XNOR2_X1 U417 ( .A(n429), .B(n363), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U419 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U420 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U422 ( .A(KEYINPUT72), .B(G92GAT), .Z(n371) );
  XNOR2_X1 U423 ( .A(G99GAT), .B(G85GAT), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U425 ( .A(G106GAT), .B(n372), .Z(n412) );
  XNOR2_X1 U426 ( .A(n376), .B(n554), .ZN(n450) );
  NAND2_X1 U427 ( .A1(n450), .A2(KEYINPUT102), .ZN(n378) );
  OR2_X1 U428 ( .A1(n450), .A2(KEYINPUT102), .ZN(n377) );
  NAND2_X1 U429 ( .A1(n378), .A2(n377), .ZN(n379) );
  XNOR2_X1 U430 ( .A(n379), .B(KEYINPUT36), .ZN(n580) );
  XOR2_X1 U431 ( .A(G78GAT), .B(G155GAT), .Z(n381) );
  XNOR2_X1 U432 ( .A(G15GAT), .B(G71GAT), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n381), .B(n380), .ZN(n397) );
  XOR2_X1 U434 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n383) );
  XNOR2_X1 U435 ( .A(G57GAT), .B(G64GAT), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n383), .B(n382), .ZN(n404) );
  XOR2_X1 U437 ( .A(n404), .B(G127GAT), .Z(n386) );
  XNOR2_X1 U438 ( .A(n384), .B(G183GAT), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U440 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n388) );
  NAND2_X1 U441 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U443 ( .A(n390), .B(n389), .Z(n395) );
  XOR2_X1 U444 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n392) );
  XNOR2_X1 U445 ( .A(G22GAT), .B(G211GAT), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n393), .B(KEYINPUT15), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n578) );
  NAND2_X1 U450 ( .A1(n580), .A2(n578), .ZN(n400) );
  XOR2_X1 U451 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n398) );
  XOR2_X1 U452 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n402) );
  XNOR2_X1 U453 ( .A(G176GAT), .B(G204GAT), .ZN(n401) );
  XNOR2_X1 U454 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U455 ( .A(n404), .B(n403), .Z(n407) );
  XOR2_X1 U456 ( .A(G148GAT), .B(G78GAT), .Z(n428) );
  XNOR2_X1 U457 ( .A(n405), .B(n428), .ZN(n406) );
  XNOR2_X1 U458 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U459 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n409) );
  NAND2_X1 U460 ( .A1(G230GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U462 ( .A(n411), .B(n410), .Z(n414) );
  XNOR2_X1 U463 ( .A(n412), .B(KEYINPUT73), .ZN(n413) );
  XNOR2_X1 U464 ( .A(n414), .B(n413), .ZN(n572) );
  NAND2_X1 U465 ( .A1(n415), .A2(n572), .ZN(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT113), .B(n416), .Z(n417) );
  NOR2_X1 U467 ( .A1(n557), .A2(n417), .ZN(n423) );
  XNOR2_X1 U468 ( .A(n572), .B(KEYINPUT41), .ZN(n547) );
  NAND2_X1 U469 ( .A1(n569), .A2(n547), .ZN(n418) );
  XNOR2_X1 U470 ( .A(KEYINPUT46), .B(n418), .ZN(n419) );
  INV_X1 U471 ( .A(n578), .ZN(n451) );
  NAND2_X1 U472 ( .A1(n419), .A2(n451), .ZN(n420) );
  NOR2_X1 U473 ( .A1(n554), .A2(n420), .ZN(n421) );
  XOR2_X1 U474 ( .A(KEYINPUT47), .B(n421), .Z(n422) );
  NOR2_X1 U475 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U476 ( .A(KEYINPUT48), .B(n424), .ZN(n541) );
  NOR2_X1 U477 ( .A1(n502), .A2(n541), .ZN(n426) );
  INV_X1 U478 ( .A(KEYINPUT54), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n426), .B(n425), .ZN(n427) );
  NOR2_X1 U480 ( .A1(n513), .A2(n427), .ZN(n568) );
  XOR2_X1 U481 ( .A(G106GAT), .B(n428), .Z(n431) );
  XNOR2_X1 U482 ( .A(G50GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U484 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n433) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U487 ( .A(n435), .B(n434), .Z(n438) );
  XNOR2_X1 U488 ( .A(n436), .B(KEYINPUT24), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U491 ( .A(n442), .B(n441), .ZN(n460) );
  NAND2_X1 U492 ( .A1(n568), .A2(n460), .ZN(n444) );
  XNOR2_X1 U493 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X2 U495 ( .A1(n504), .A2(n445), .ZN(n562) );
  NAND2_X1 U496 ( .A1(n562), .A2(n547), .ZN(n449) );
  XOR2_X1 U497 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n447) );
  XNOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n557), .A2(n572), .ZN(n484) );
  BUF_X1 U500 ( .A(n450), .Z(n561) );
  NOR2_X1 U501 ( .A1(n561), .A2(n451), .ZN(n452) );
  XNOR2_X1 U502 ( .A(n452), .B(KEYINPUT16), .ZN(n468) );
  XNOR2_X1 U503 ( .A(KEYINPUT84), .B(n504), .ZN(n455) );
  XOR2_X1 U504 ( .A(KEYINPUT27), .B(n502), .Z(n462) );
  NAND2_X1 U505 ( .A1(n462), .A2(n513), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(KEYINPUT94), .ZN(n544) );
  XOR2_X1 U507 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n454) );
  XNOR2_X1 U508 ( .A(n460), .B(n454), .ZN(n521) );
  NOR2_X1 U509 ( .A1(n544), .A2(n521), .ZN(n527) );
  NAND2_X1 U510 ( .A1(n455), .A2(n527), .ZN(n467) );
  INV_X1 U511 ( .A(n513), .ZN(n498) );
  INV_X1 U512 ( .A(n504), .ZN(n526) );
  INV_X1 U513 ( .A(n502), .ZN(n515) );
  NAND2_X1 U514 ( .A1(n526), .A2(n515), .ZN(n456) );
  NAND2_X1 U515 ( .A1(n456), .A2(n460), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT96), .ZN(n458) );
  XNOR2_X1 U517 ( .A(KEYINPUT25), .B(n458), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT95), .ZN(n464) );
  NOR2_X1 U519 ( .A1(n526), .A2(n460), .ZN(n461) );
  XNOR2_X1 U520 ( .A(KEYINPUT26), .B(n461), .ZN(n567) );
  NAND2_X1 U521 ( .A1(n462), .A2(n567), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n498), .A2(n465), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n481) );
  NAND2_X1 U525 ( .A1(n468), .A2(n481), .ZN(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT97), .B(n469), .Z(n496) );
  NOR2_X1 U527 ( .A1(n484), .A2(n496), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT98), .ZN(n478) );
  NAND2_X1 U529 ( .A1(n513), .A2(n478), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  NAND2_X1 U533 ( .A1(n478), .A2(n515), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT100), .ZN(n475) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(n475), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U537 ( .A1(n478), .A2(n526), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  XOR2_X1 U539 ( .A(G22GAT), .B(KEYINPUT101), .Z(n480) );
  NAND2_X1 U540 ( .A1(n521), .A2(n478), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1327GAT) );
  XOR2_X1 U542 ( .A(G29GAT), .B(KEYINPUT39), .Z(n487) );
  NAND2_X1 U543 ( .A1(n580), .A2(n481), .ZN(n482) );
  NOR2_X1 U544 ( .A1(n482), .A2(n578), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n483), .B(KEYINPUT37), .ZN(n511) );
  NOR2_X1 U546 ( .A1(n511), .A2(n484), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n485), .B(KEYINPUT38), .ZN(n492) );
  NAND2_X1 U548 ( .A1(n513), .A2(n492), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  XOR2_X1 U550 ( .A(G36GAT), .B(KEYINPUT103), .Z(n489) );
  NAND2_X1 U551 ( .A1(n515), .A2(n492), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n492), .A2(n526), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  NAND2_X1 U556 ( .A1(n492), .A2(n521), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U558 ( .A(n547), .ZN(n494) );
  NOR2_X1 U559 ( .A1(n569), .A2(n494), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n495), .B(KEYINPUT105), .ZN(n510) );
  NOR2_X1 U561 ( .A1(n496), .A2(n510), .ZN(n497) );
  XOR2_X1 U562 ( .A(KEYINPUT106), .B(n497), .Z(n507) );
  NOR2_X1 U563 ( .A1(n507), .A2(n498), .ZN(n500) );
  XNOR2_X1 U564 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n501), .Z(G1332GAT) );
  NOR2_X1 U567 ( .A1(n507), .A2(n502), .ZN(n503) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n504), .A2(n507), .ZN(n505) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  INV_X1 U571 ( .A(n521), .ZN(n506) );
  NOR2_X1 U572 ( .A1(n507), .A2(n506), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NOR2_X1 U575 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U576 ( .A(KEYINPUT107), .B(n512), .Z(n522) );
  NAND2_X1 U577 ( .A1(n513), .A2(n522), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n522), .A2(n515), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(KEYINPUT108), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n519) );
  NAND2_X1 U583 ( .A1(n522), .A2(n526), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n520), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n524) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n541), .A2(n528), .ZN(n529) );
  XNOR2_X1 U592 ( .A(KEYINPUT114), .B(n529), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n557), .A2(n536), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U596 ( .A1(n536), .A2(n547), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U598 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n578), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U603 ( .A1(n561), .A2(n536), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n540) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT116), .Z(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n546) );
  INV_X1 U608 ( .A(n541), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n542), .A2(n567), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n555), .A2(n569), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U614 ( .A1(n555), .A2(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .Z(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n578), .A2(n555), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT120), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n562), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(G183GAT), .B(KEYINPUT123), .Z(n560) );
  NAND2_X1 U626 ( .A1(n562), .A2(n578), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT58), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT124), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(n566), .Z(n571) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n573) );
  INV_X1 U635 ( .A(n573), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n581), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n581), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n583) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

