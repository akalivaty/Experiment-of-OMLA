

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582;

  XNOR2_X1 U324 ( .A(n444), .B(KEYINPUT55), .ZN(n445) );
  AND2_X1 U325 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U326 ( .A(n362), .B(n292), .ZN(n342) );
  INV_X1 U327 ( .A(KEYINPUT121), .ZN(n444) );
  XNOR2_X1 U328 ( .A(n343), .B(n342), .ZN(n345) );
  XNOR2_X1 U329 ( .A(n393), .B(KEYINPUT48), .ZN(n394) );
  XNOR2_X1 U330 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U331 ( .A(n395), .B(n394), .ZN(n538) );
  XOR2_X1 U332 ( .A(n312), .B(n311), .Z(n492) );
  XNOR2_X1 U333 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U334 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n294) );
  XNOR2_X1 U336 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n312) );
  XOR2_X1 U338 ( .A(G176GAT), .B(G99GAT), .Z(n296) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(G43GAT), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U341 ( .A(G127GAT), .B(G71GAT), .Z(n298) );
  XNOR2_X1 U342 ( .A(G15GAT), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(n300), .B(n299), .Z(n310) );
  XOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT87), .Z(n302) );
  XNOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U348 ( .A(G120GAT), .B(n303), .Z(n425) );
  XOR2_X1 U349 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n305) );
  XNOR2_X1 U350 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n403) );
  XOR2_X1 U352 ( .A(n403), .B(KEYINPUT20), .Z(n307) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n425), .B(n308), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U357 ( .A(G22GAT), .B(G15GAT), .Z(n354) );
  XOR2_X1 U358 ( .A(G141GAT), .B(KEYINPUT30), .Z(n314) );
  XNOR2_X1 U359 ( .A(G197GAT), .B(G1GAT), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U361 ( .A(n354), .B(n315), .Z(n317) );
  NAND2_X1 U362 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U363 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U364 ( .A(n318), .B(KEYINPUT68), .Z(n321) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G36GAT), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n319), .B(G8GAT), .ZN(n396) );
  XNOR2_X1 U367 ( .A(n396), .B(KEYINPUT29), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n331) );
  XOR2_X1 U369 ( .A(G50GAT), .B(G29GAT), .Z(n323) );
  XNOR2_X1 U370 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U372 ( .A(n324), .B(KEYINPUT70), .Z(n326) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n383) );
  XOR2_X1 U375 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n328) );
  XNOR2_X1 U376 ( .A(G113GAT), .B(KEYINPUT73), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U378 ( .A(n383), .B(n329), .Z(n330) );
  XOR2_X1 U379 ( .A(n331), .B(n330), .Z(n565) );
  XOR2_X1 U380 ( .A(G92GAT), .B(G64GAT), .Z(n333) );
  XNOR2_X1 U381 ( .A(G176GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U383 ( .A(KEYINPUT78), .B(n334), .ZN(n406) );
  XOR2_X1 U384 ( .A(G106GAT), .B(G78GAT), .Z(n336) );
  XNOR2_X1 U385 ( .A(G148GAT), .B(KEYINPUT76), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U387 ( .A(KEYINPUT77), .B(n337), .Z(n438) );
  XOR2_X1 U388 ( .A(n406), .B(n438), .Z(n347) );
  XOR2_X1 U389 ( .A(G99GAT), .B(G85GAT), .Z(n377) );
  XOR2_X1 U390 ( .A(KEYINPUT33), .B(KEYINPUT79), .Z(n339) );
  XNOR2_X1 U391 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U393 ( .A(n377), .B(n340), .Z(n343) );
  XNOR2_X1 U394 ( .A(G71GAT), .B(KEYINPUT75), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n341), .B(KEYINPUT13), .ZN(n362) );
  XNOR2_X1 U396 ( .A(G120GAT), .B(G57GAT), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n570) );
  XNOR2_X1 U399 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n570), .B(n348), .ZN(n543) );
  NOR2_X1 U401 ( .A1(n565), .A2(n543), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n349), .B(KEYINPUT46), .ZN(n367) );
  XOR2_X1 U403 ( .A(KEYINPUT14), .B(G78GAT), .Z(n351) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(G64GAT), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n366) );
  XOR2_X1 U406 ( .A(G155GAT), .B(G57GAT), .Z(n353) );
  XNOR2_X1 U407 ( .A(G1GAT), .B(G127GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n415) );
  XOR2_X1 U409 ( .A(n415), .B(n354), .Z(n356) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT84), .B(KEYINPUT12), .Z(n358) );
  XNOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT85), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U415 ( .A(n360), .B(n359), .Z(n364) );
  XNOR2_X1 U416 ( .A(G183GAT), .B(KEYINPUT83), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n361), .B(G211GAT), .ZN(n402) );
  XNOR2_X1 U418 ( .A(n362), .B(n402), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n575) );
  XNOR2_X1 U421 ( .A(KEYINPUT110), .B(n575), .ZN(n557) );
  NOR2_X1 U422 ( .A1(n367), .A2(n557), .ZN(n386) );
  XOR2_X1 U423 ( .A(KEYINPUT82), .B(G218GAT), .Z(n369) );
  XNOR2_X1 U424 ( .A(G36GAT), .B(G134GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U426 ( .A(KEYINPUT80), .B(KEYINPUT10), .Z(n371) );
  XNOR2_X1 U427 ( .A(G162GAT), .B(KEYINPUT66), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U429 ( .A(n373), .B(n372), .Z(n379) );
  XOR2_X1 U430 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n375) );
  NAND2_X1 U431 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n385) );
  XOR2_X1 U435 ( .A(KEYINPUT81), .B(G106GAT), .Z(n381) );
  XNOR2_X1 U436 ( .A(G190GAT), .B(G92GAT), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U438 ( .A(n383), .B(n382), .Z(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n551) );
  NAND2_X1 U440 ( .A1(n386), .A2(n551), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n387), .B(KEYINPUT47), .ZN(n392) );
  XNOR2_X1 U442 ( .A(KEYINPUT36), .B(n551), .ZN(n580) );
  INV_X1 U443 ( .A(n575), .ZN(n547) );
  NOR2_X1 U444 ( .A1(n580), .A2(n547), .ZN(n388) );
  XNOR2_X1 U445 ( .A(KEYINPUT45), .B(n388), .ZN(n389) );
  NAND2_X1 U446 ( .A1(n389), .A2(n570), .ZN(n390) );
  XOR2_X1 U447 ( .A(KEYINPUT74), .B(n565), .Z(n554) );
  NOR2_X1 U448 ( .A1(n390), .A2(n554), .ZN(n391) );
  NOR2_X1 U449 ( .A1(n392), .A2(n391), .ZN(n395) );
  XOR2_X1 U450 ( .A(KEYINPUT64), .B(KEYINPUT111), .Z(n393) );
  XOR2_X1 U451 ( .A(KEYINPUT98), .B(n396), .Z(n398) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n401) );
  XOR2_X1 U454 ( .A(KEYINPUT21), .B(KEYINPUT92), .Z(n400) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n433) );
  XOR2_X1 U457 ( .A(n401), .B(n433), .Z(n405) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n407) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n512) );
  XOR2_X1 U461 ( .A(KEYINPUT120), .B(n512), .Z(n408) );
  NOR2_X1 U462 ( .A1(n538), .A2(n408), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n409), .B(KEYINPUT54), .ZN(n428) );
  XOR2_X1 U464 ( .A(KEYINPUT6), .B(KEYINPUT96), .Z(n411) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U467 ( .A(n412), .B(KEYINPUT4), .Z(n417) );
  XOR2_X1 U468 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n414) );
  XNOR2_X1 U469 ( .A(G141GAT), .B(G162GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n439) );
  XNOR2_X1 U471 ( .A(n415), .B(n439), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U473 ( .A(KEYINPUT5), .B(G148GAT), .Z(n419) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G85GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n421), .B(n420), .Z(n427) );
  XOR2_X1 U477 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n423) );
  XNOR2_X1 U478 ( .A(KEYINPUT93), .B(KEYINPUT95), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n465) );
  XNOR2_X1 U482 ( .A(KEYINPUT97), .B(n465), .ZN(n484) );
  NAND2_X1 U483 ( .A1(n428), .A2(n484), .ZN(n564) );
  XOR2_X1 U484 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n430) );
  XNOR2_X1 U485 ( .A(G22GAT), .B(G155GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n443) );
  XOR2_X1 U487 ( .A(G211GAT), .B(KEYINPUT80), .Z(n432) );
  XNOR2_X1 U488 ( .A(G50GAT), .B(G204GAT), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n437) );
  XOR2_X1 U490 ( .A(n433), .B(KEYINPUT24), .Z(n435) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U493 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U496 ( .A(n443), .B(n442), .Z(n458) );
  NOR2_X1 U497 ( .A1(n564), .A2(n458), .ZN(n446) );
  NOR2_X1 U498 ( .A1(n492), .A2(n447), .ZN(n559) );
  INV_X1 U499 ( .A(n543), .ZN(n527) );
  NAND2_X1 U500 ( .A1(n559), .A2(n527), .ZN(n451) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT57), .Z(n449) );
  XOR2_X1 U502 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n448) );
  NAND2_X1 U503 ( .A1(n554), .A2(n570), .ZN(n482) );
  XOR2_X1 U504 ( .A(KEYINPUT16), .B(KEYINPUT86), .Z(n453) );
  NAND2_X1 U505 ( .A1(n575), .A2(n551), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n469) );
  XOR2_X1 U507 ( .A(n512), .B(KEYINPUT27), .Z(n461) );
  OR2_X1 U508 ( .A1(n484), .A2(n461), .ZN(n537) );
  XOR2_X1 U509 ( .A(n458), .B(KEYINPUT67), .Z(n454) );
  XNOR2_X1 U510 ( .A(KEYINPUT28), .B(n454), .ZN(n517) );
  NOR2_X1 U511 ( .A1(n537), .A2(n517), .ZN(n521) );
  NAND2_X1 U512 ( .A1(n492), .A2(n521), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT99), .ZN(n467) );
  INV_X1 U514 ( .A(n512), .ZN(n488) );
  NOR2_X1 U515 ( .A1(n492), .A2(n488), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n458), .A2(n456), .ZN(n457) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(n457), .Z(n463) );
  NAND2_X1 U518 ( .A1(n458), .A2(n492), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n459), .B(KEYINPUT100), .ZN(n460) );
  XNOR2_X1 U520 ( .A(KEYINPUT26), .B(n460), .ZN(n563) );
  NOR2_X1 U521 ( .A1(n461), .A2(n563), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U525 ( .A(KEYINPUT101), .B(n468), .ZN(n479) );
  NAND2_X1 U526 ( .A1(n469), .A2(n479), .ZN(n498) );
  NOR2_X1 U527 ( .A1(n482), .A2(n498), .ZN(n477) );
  INV_X1 U528 ( .A(n484), .ZN(n510) );
  NAND2_X1 U529 ( .A1(n477), .A2(n510), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U532 ( .A1(n477), .A2(n512), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(KEYINPUT102), .ZN(n473) );
  XNOR2_X1 U534 ( .A(G8GAT), .B(n473), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n475) );
  INV_X1 U536 ( .A(n492), .ZN(n520) );
  NAND2_X1 U537 ( .A1(n477), .A2(n520), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U539 ( .A(G15GAT), .B(n476), .Z(G1326GAT) );
  NAND2_X1 U540 ( .A1(n517), .A2(n477), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n478), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U542 ( .A1(n547), .A2(n479), .ZN(n480) );
  NOR2_X1 U543 ( .A1(n580), .A2(n480), .ZN(n481) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n481), .ZN(n509) );
  NOR2_X1 U545 ( .A1(n509), .A2(n482), .ZN(n483) );
  XOR2_X1 U546 ( .A(KEYINPUT38), .B(n483), .Z(n495) );
  NOR2_X1 U547 ( .A1(n495), .A2(n484), .ZN(n486) );
  XNOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT39), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(n487), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n495), .A2(n488), .ZN(n489) );
  XOR2_X1 U552 ( .A(G36GAT), .B(n489), .Z(G1329GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n491) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(n494) );
  NOR2_X1 U556 ( .A1(n492), .A2(n495), .ZN(n493) );
  XOR2_X1 U557 ( .A(n494), .B(n493), .Z(G1330GAT) );
  INV_X1 U558 ( .A(n517), .ZN(n496) );
  NOR2_X1 U559 ( .A1(n496), .A2(n495), .ZN(n497) );
  XOR2_X1 U560 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n500) );
  NAND2_X1 U562 ( .A1(n565), .A2(n527), .ZN(n508) );
  NOR2_X1 U563 ( .A1(n508), .A2(n498), .ZN(n504) );
  NAND2_X1 U564 ( .A1(n510), .A2(n504), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n512), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n501), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U568 ( .A(G71GAT), .B(KEYINPUT107), .Z(n503) );
  NAND2_X1 U569 ( .A1(n504), .A2(n520), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n517), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n507), .ZN(G1335GAT) );
  NOR2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n510), .A2(n516), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n516), .A2(n512), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U580 ( .A(G99GAT), .B(KEYINPUT109), .Z(n515) );
  NAND2_X1 U581 ( .A1(n516), .A2(n520), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1338GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT44), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U587 ( .A1(n538), .A2(n522), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n533), .A2(n554), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n525) );
  XNOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT112), .B(n526), .Z(n529) );
  NAND2_X1 U594 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n531) );
  NAND2_X1 U597 ( .A1(n533), .A2(n557), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n535) );
  INV_X1 U601 ( .A(n551), .ZN(n560) );
  NAND2_X1 U602 ( .A1(n533), .A2(n560), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n536), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n563), .A2(n537), .ZN(n540) );
  INV_X1 U606 ( .A(n538), .ZN(n539) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n565), .A2(n550), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  NOR2_X1 U611 ( .A1(n543), .A2(n550), .ZN(n545) );
  XNOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n547), .A2(n550), .ZN(n548) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(n548), .Z(n549) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n549), .ZN(G1346GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n559), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(KEYINPUT122), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1351GAT) );
  XNOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT124), .Z(n567) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n576) );
  INV_X1 U632 ( .A(n576), .ZN(n579) );
  OR2_X1 U633 ( .A1(n579), .A2(n565), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n579), .A2(n570), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n572) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT127), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

