//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n209), .B1(new_n213), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(G232), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT2), .B(G226), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n227), .B(new_n230), .Z(G358));
  XOR2_X1   g0031(.A(G87), .B(G97), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G107), .B(G116), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G58), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  INV_X1    g0039(.A(KEYINPUT10), .ZN(new_n240));
  NAND3_X1  g0040(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n241));
  INV_X1    g0041(.A(KEYINPUT67), .ZN(new_n242));
  AND3_X1   g0042(.A1(new_n241), .A2(new_n242), .A3(new_n210), .ZN(new_n243));
  AOI21_X1  g0043(.A(new_n242), .B1(new_n241), .B2(new_n210), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G50), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n211), .B1(new_n201), .B2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n252), .A2(new_n254), .B1(G150), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n246), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n258), .A2(new_n211), .A3(G1), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n257), .B1(new_n247), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n241), .A2(new_n210), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT67), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n241), .A2(new_n242), .A3(new_n210), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n211), .A2(G1), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G50), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n260), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n253), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1698), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G222), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n275), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G223), .A3(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n279), .C1(new_n280), .C2(new_n278), .ZN(new_n281));
  AND2_X1   g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n210), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(G1), .B(G13), .C1(new_n253), .C2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G41), .A2(G45), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G1), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n288), .A3(G274), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT66), .B1(new_n287), .B2(G1), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT66), .ZN(new_n292));
  INV_X1    g0092(.A(G1), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n292), .B(new_n293), .C1(G41), .C2(G45), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n291), .A2(new_n286), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n290), .B1(new_n295), .B2(G226), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n284), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n240), .B1(new_n272), .B2(new_n303), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n300), .A2(KEYINPUT10), .A3(new_n302), .ZN(new_n305));
  INV_X1    g0105(.A(new_n271), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n270), .B1(new_n260), .B2(new_n267), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n306), .A2(KEYINPUT71), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT71), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n269), .B2(new_n271), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n305), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT72), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT71), .B1(new_n306), .B2(new_n307), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n269), .A2(new_n309), .A3(new_n271), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT72), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n305), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n304), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT16), .ZN(new_n319));
  INV_X1    g0119(.A(G68), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n274), .A2(new_n211), .A3(new_n275), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n275), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(G58), .A2(G68), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n328), .B2(new_n201), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n255), .A2(G159), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n319), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  NOR2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(new_n324), .A3(new_n211), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n321), .A2(KEYINPUT7), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(G68), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n246), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n291), .A2(new_n286), .A3(G232), .A4(new_n294), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n342), .A2(new_n289), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G87), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT76), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(G226), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n347));
  INV_X1    g0147(.A(G1698), .ZN(new_n348));
  OAI211_X1 g0148(.A(G223), .B(new_n348), .C1(new_n333), .C2(new_n334), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n283), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G200), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n251), .A2(new_n265), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n264), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n251), .A2(new_n259), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n343), .A2(new_n351), .A3(G190), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n341), .A2(new_n353), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT17), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n343), .A2(new_n351), .A3(G190), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n299), .B1(new_n343), .B2(new_n351), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n357), .B1(new_n332), .B2(new_n340), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(KEYINPUT17), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n341), .A2(new_n358), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n343), .A2(new_n351), .A3(G179), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n342), .A2(new_n289), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n283), .B2(new_n350), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n369), .A2(KEYINPUT77), .A3(KEYINPUT18), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n343), .A2(new_n351), .A3(G179), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n343), .B2(new_n351), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n376), .B1(new_n379), .B2(new_n366), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n369), .A2(KEYINPUT18), .A3(new_n374), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n368), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n264), .A2(G68), .A3(new_n266), .ZN(new_n386));
  XOR2_X1   g0186(.A(new_n386), .B(KEYINPUT73), .Z(new_n387));
  INV_X1    g0187(.A(new_n255), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n247), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n211), .A2(G33), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n390), .A2(new_n280), .B1(new_n211), .B2(G68), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n245), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT11), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n258), .A2(G1), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G20), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT74), .B1(new_n395), .B2(G68), .ZN(new_n396));
  XOR2_X1   g0196(.A(new_n396), .B(KEYINPUT12), .Z(new_n397));
  NAND3_X1  g0197(.A1(new_n387), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT14), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n276), .A2(G226), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n278), .A2(G232), .A3(G1698), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G97), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n283), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n290), .B1(new_n295), .B2(G238), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n404), .B2(new_n405), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n399), .B(G169), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G179), .ZN(new_n411));
  INV_X1    g0211(.A(new_n409), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n407), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n410), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n399), .B1(new_n413), .B2(G169), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n398), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n398), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(G200), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n412), .A2(G190), .A3(new_n407), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n291), .A2(new_n286), .A3(G244), .A4(new_n294), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n289), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT69), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT69), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(new_n424), .A3(new_n289), .ZN(new_n425));
  OAI211_X1 g0225(.A(G232), .B(new_n348), .C1(new_n333), .C2(new_n334), .ZN(new_n426));
  OAI211_X1 g0226(.A(G238), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n427));
  INV_X1    g0227(.A(G107), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n426), .B(new_n427), .C1(new_n428), .C2(new_n278), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n283), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n423), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G200), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G20), .A2(G77), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n433), .B1(new_n251), .B2(new_n388), .C1(new_n390), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n245), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n264), .A2(G77), .A3(new_n266), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n259), .A2(new_n280), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT70), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n423), .A2(G190), .A3(new_n430), .A4(new_n425), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n432), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n431), .A2(new_n373), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n423), .A2(new_n411), .A3(new_n430), .A4(new_n425), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n440), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n385), .A2(new_n416), .A3(new_n420), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n298), .A2(new_n411), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n297), .A2(new_n373), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n268), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n318), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n293), .A2(G33), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n395), .B(new_n455), .C1(new_n243), .C2(new_n244), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n264), .A2(KEYINPUT80), .A3(G116), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n461), .B(new_n211), .C1(G33), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n457), .A2(G20), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n261), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n466), .ZN(new_n468));
  INV_X1    g0268(.A(new_n464), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n467), .A2(new_n468), .B1(new_n394), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n278), .A2(G264), .A3(G1698), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n278), .A2(G257), .A3(new_n348), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n335), .A2(G303), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n283), .ZN(new_n476));
  INV_X1    g0276(.A(G45), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(G270), .A3(new_n286), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(new_n286), .A3(G274), .A4(new_n478), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n482), .A2(new_n484), .A3(KEYINPUT79), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT79), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n476), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT21), .A3(G169), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n476), .B(G179), .C1(new_n485), .C2(new_n486), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n471), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT21), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(G169), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n471), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT81), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n491), .C1(new_n471), .C2(new_n492), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n487), .A2(G200), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n471), .B(new_n498), .C1(new_n301), .C2(new_n487), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT87), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n481), .A2(G264), .A3(new_n286), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT85), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n481), .A2(new_n504), .A3(G264), .A4(new_n286), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(G274), .B1(new_n282), .B2(new_n210), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n481), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n509));
  OAI211_X1 g0309(.A(G250), .B(new_n348), .C1(new_n333), .C2(new_n334), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n512), .B2(new_n283), .ZN(new_n513));
  AOI211_X1 g0313(.A(new_n501), .B(G200), .C1(new_n506), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n506), .A2(new_n513), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT87), .B1(new_n515), .B2(G190), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n299), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT82), .B1(new_n211), .B2(G107), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT23), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  OAI211_X1 g0321(.A(KEYINPUT82), .B(new_n521), .C1(new_n211), .C2(G107), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n520), .A2(new_n522), .B1(G116), .B2(new_n254), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  AOI21_X1  g0324(.A(G20), .B1(new_n274), .B2(new_n275), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G87), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n211), .B(G87), .C1(new_n333), .C2(new_n334), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n523), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n278), .A2(new_n524), .A3(new_n211), .A4(G87), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(KEYINPUT83), .A3(new_n523), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(KEYINPUT24), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT83), .B1(new_n534), .B2(new_n523), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n246), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n428), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT84), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT25), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n395), .B2(G107), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n544), .ZN(new_n546));
  INV_X1    g0346(.A(new_n456), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n545), .A2(new_n546), .B1(G107), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n518), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n515), .A2(G169), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n411), .B2(new_n515), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT86), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT86), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n552), .B(new_n555), .C1(new_n411), .C2(new_n515), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n549), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G250), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(new_n348), .C1(new_n333), .C2(new_n334), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n461), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT4), .B1(new_n276), .B2(G244), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n283), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n481), .A2(G257), .A3(new_n286), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n484), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n373), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n255), .A2(G77), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  AND2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n428), .A2(KEYINPUT6), .A3(G97), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n568), .B1(new_n575), .B2(new_n211), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n428), .B1(new_n325), .B2(new_n326), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n245), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n395), .A2(G97), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n456), .B2(new_n462), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n565), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n560), .A2(new_n561), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n348), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n461), .A4(new_n559), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n587), .B2(new_n283), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n411), .A3(new_n484), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n567), .A2(new_n583), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n566), .A2(G200), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n333), .A2(new_n334), .A3(G20), .ZN(new_n592));
  XNOR2_X1  g0392(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n326), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G107), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n574), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n581), .B1(new_n597), .B2(new_n245), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n564), .A2(G190), .A3(new_n484), .A4(new_n565), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n591), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n434), .A2(new_n259), .ZN(new_n601));
  INV_X1    g0401(.A(new_n434), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n264), .A2(new_n602), .A3(new_n455), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n211), .B(G68), .C1(new_n333), .C2(new_n334), .ZN(new_n604));
  XOR2_X1   g0404(.A(KEYINPUT78), .B(KEYINPUT19), .Z(new_n605));
  NOR2_X1   g0405(.A1(new_n390), .A2(new_n462), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g0407(.A(KEYINPUT78), .B(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n211), .B1(new_n608), .B2(new_n402), .ZN(new_n609));
  INV_X1    g0409(.A(G87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n571), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n607), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n601), .B(new_n603), .C1(new_n612), .C2(new_n246), .ZN(new_n613));
  OAI211_X1 g0413(.A(G238), .B(new_n348), .C1(new_n333), .C2(new_n334), .ZN(new_n614));
  OAI211_X1 g0414(.A(G244), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n614), .B(new_n615), .C1(new_n253), .C2(new_n457), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n283), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n293), .A2(G45), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G250), .ZN(new_n619));
  OAI22_X1  g0419(.A1(new_n507), .A2(new_n618), .B1(new_n283), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n373), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n616), .B2(new_n283), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n411), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n613), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(G200), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n609), .A2(new_n611), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n254), .A2(G97), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n525), .A2(G68), .B1(new_n629), .B2(new_n608), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n245), .B1(new_n259), .B2(new_n434), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n547), .A2(G87), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(G190), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n627), .A2(new_n632), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n590), .A2(new_n600), .A3(new_n626), .A4(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n500), .A2(new_n558), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n453), .A2(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n453), .ZN(new_n639));
  INV_X1    g0439(.A(new_n490), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n549), .A2(new_n553), .ZN(new_n641));
  INV_X1    g0441(.A(new_n496), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n460), .A2(new_n470), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(G169), .A3(new_n487), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n495), .B1(new_n644), .B2(new_n491), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n550), .A2(new_n636), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n635), .A2(new_n626), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n567), .A2(new_n583), .A3(new_n589), .ZN(new_n650));
  XOR2_X1   g0450(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n635), .A2(new_n626), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT26), .B1(new_n653), .B2(new_n590), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n652), .A2(new_n626), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n639), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT89), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n379), .A2(new_n366), .A3(new_n376), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT18), .B1(new_n369), .B2(new_n374), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n416), .B1(new_n661), .B2(new_n446), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n359), .B1(new_n372), .B2(new_n299), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n369), .A2(new_n663), .A3(new_n361), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT17), .B1(new_n365), .B2(new_n366), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n660), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n451), .B1(new_n318), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n657), .A2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n394), .A2(new_n211), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n471), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n500), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n497), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT91), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n558), .ZN(new_n687));
  INV_X1    g0487(.A(new_n549), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n678), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n557), .B2(new_n678), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n641), .A2(new_n677), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n497), .A2(new_n677), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n207), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n611), .A2(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n214), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g0501(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n702));
  XNOR2_X1  g0502(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AOI211_X1 g0503(.A(new_n550), .B(new_n636), .C1(new_n497), .C2(new_n557), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n649), .A2(new_n650), .ZN(new_n705));
  INV_X1    g0505(.A(new_n651), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n707), .B(new_n626), .C1(KEYINPUT26), .C2(new_n705), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n677), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n677), .B1(new_n648), .B2(new_n655), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n558), .A2(new_n636), .ZN(new_n714));
  INV_X1    g0514(.A(new_n500), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(new_n678), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n566), .A2(new_n515), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n487), .A2(new_n411), .A3(new_n622), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT93), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT93), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n487), .A2(new_n720), .A3(new_n411), .A4(new_n622), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n717), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n588), .A2(new_n506), .A3(new_n513), .A4(new_n624), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n489), .ZN(new_n725));
  INV_X1    g0525(.A(new_n489), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n515), .A2(new_n622), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(KEYINPUT30), .A4(new_n588), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n677), .B1(new_n722), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT31), .B(new_n677), .C1(new_n722), .C2(new_n729), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n716), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n711), .A2(new_n713), .B1(new_n734), .B2(G330), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n703), .B1(new_n735), .B2(G1), .ZN(G364));
  XNOR2_X1  g0536(.A(new_n684), .B(KEYINPUT91), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n258), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n293), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n697), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n737), .B(new_n742), .C1(G330), .C2(new_n683), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n210), .B1(G20), .B2(new_n373), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n211), .A2(new_n411), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(new_n301), .A3(new_n299), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G20), .A3(new_n301), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n748), .A2(G311), .B1(new_n751), .B2(G329), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n211), .A2(new_n301), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(G179), .A3(new_n299), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n752), .B(new_n335), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n211), .B1(new_n749), .B2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n756), .B1(G294), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT95), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n411), .B2(G200), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n299), .A2(KEYINPUT95), .A3(G179), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n754), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n763), .A2(new_n211), .A3(G190), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n766), .A2(G303), .B1(new_n767), .B2(G283), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n211), .A2(new_n411), .A3(new_n299), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT94), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n301), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(G190), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G326), .A2(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n759), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n278), .B1(new_n747), .B2(new_n280), .ZN(new_n776));
  INV_X1    g0576(.A(new_n755), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(G58), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n767), .A2(G107), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  OR3_X1    g0581(.A1(new_n750), .A2(KEYINPUT32), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n758), .A2(G97), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT32), .B1(new_n750), .B2(new_n781), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n772), .B2(G68), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n766), .A2(G87), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n771), .A2(G50), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n780), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n745), .B1(new_n775), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n744), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n696), .A2(new_n335), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G355), .A2(new_n795), .B1(new_n457), .B2(new_n696), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n238), .A2(new_n477), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n696), .A2(new_n278), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n214), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n742), .B(new_n790), .C1(new_n794), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n793), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n683), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n743), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n440), .A2(new_n677), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n443), .A2(new_n446), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT99), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n807), .B(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n677), .B(new_n809), .C1(new_n648), .C2(new_n655), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n446), .A2(new_n678), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(new_n712), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n734), .A2(G330), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n741), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n744), .A2(new_n791), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n741), .B1(G77), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT96), .B(G283), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G303), .A2(new_n771), .B1(new_n772), .B2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n777), .A2(G294), .B1(new_n748), .B2(G116), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n278), .B1(new_n751), .B2(G311), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n824), .A2(new_n783), .A3(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n766), .A2(G107), .B1(new_n767), .B2(G87), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n777), .A2(G143), .B1(new_n748), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(new_n771), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  INV_X1    g0632(.A(new_n772), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n829), .B1(new_n830), .B2(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT97), .Z(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n767), .A2(G68), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n247), .B2(new_n765), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT98), .Z(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n278), .B1(new_n750), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G58), .B2(new_n758), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n836), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n828), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n820), .B1(new_n845), .B2(new_n744), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n792), .B2(new_n813), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n817), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  NOR2_X1   g0649(.A1(new_n738), .A2(new_n293), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n320), .B1(new_n321), .B2(KEYINPUT7), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n331), .B1(new_n851), .B2(new_n336), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT101), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT16), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n331), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT7), .ZN(new_n856));
  OAI21_X1  g0656(.A(G68), .B1(new_n592), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n321), .A2(new_n593), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT101), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n357), .B1(new_n861), .B2(new_n340), .ZN(new_n862));
  OAI211_X1 g0662(.A(KEYINPUT103), .B(new_n360), .C1(new_n862), .C2(new_n379), .ZN(new_n863));
  INV_X1    g0663(.A(new_n675), .ZN(new_n864));
  INV_X1    g0664(.A(new_n340), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n860), .B2(new_n854), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n864), .B1(new_n866), .B2(new_n357), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n374), .B1(new_n866), .B2(new_n357), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT103), .B1(new_n869), .B2(new_n360), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n369), .A2(KEYINPUT104), .A3(new_n374), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n369), .A2(new_n864), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n360), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n352), .A2(G169), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n341), .A2(new_n358), .B1(new_n876), .B2(new_n370), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n877), .B2(KEYINPUT104), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n384), .A2(new_n375), .A3(new_n380), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n881), .B(new_n867), .C1(new_n882), .C2(new_n666), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n375), .A2(new_n380), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT77), .B1(new_n877), .B2(KEYINPUT18), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n666), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n867), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT102), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n880), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n880), .B(KEYINPUT38), .C1(new_n883), .C2(new_n888), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT100), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n446), .A2(new_n677), .ZN(new_n895));
  INV_X1    g0695(.A(new_n809), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n712), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n398), .A2(new_n677), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n416), .A2(new_n420), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n898), .B1(new_n416), .B2(new_n420), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n894), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT105), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n889), .A2(new_n904), .A3(new_n890), .ZN(new_n905));
  INV_X1    g0705(.A(new_n901), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n899), .ZN(new_n907));
  OAI211_X1 g0707(.A(KEYINPUT100), .B(new_n907), .C1(new_n810), .C2(new_n895), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n893), .A2(new_n903), .A3(new_n905), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n660), .A2(new_n675), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n414), .A2(new_n415), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n398), .A3(new_n678), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n893), .B2(new_n905), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n369), .A2(new_n663), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n366), .A2(new_n675), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n917), .A2(new_n877), .A3(new_n918), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n919), .A2(new_n875), .B1(new_n874), .B2(new_n878), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT106), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n918), .B1(new_n660), .B2(new_n368), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT107), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n873), .A2(new_n360), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT37), .B1(new_n926), .B2(new_n877), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(KEYINPUT106), .C1(new_n878), .C2(new_n874), .ZN(new_n928));
  OAI211_X1 g0728(.A(KEYINPUT107), .B(new_n918), .C1(new_n660), .C2(new_n368), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n922), .A2(new_n925), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n890), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n892), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n915), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n916), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n911), .B1(new_n914), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n711), .A2(new_n453), .A3(new_n713), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n670), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G330), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n813), .B1(new_n900), .B2(new_n901), .ZN(new_n941));
  INV_X1    g0741(.A(new_n733), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n637), .B2(new_n678), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT108), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n730), .A2(new_n945), .A3(new_n731), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n941), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n893), .A2(new_n948), .A3(new_n905), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n716), .A2(new_n733), .A3(new_n944), .A4(new_n946), .ZN(new_n952));
  INV_X1    g0752(.A(new_n941), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n952), .A2(KEYINPUT40), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT109), .B1(new_n931), .B2(new_n892), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n931), .A2(KEYINPUT109), .A3(new_n892), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n453), .A2(new_n952), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n940), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n850), .B1(new_n939), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n939), .B2(new_n962), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n457), .B(new_n213), .C1(new_n574), .C2(KEYINPUT35), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(KEYINPUT35), .B2(new_n574), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT36), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n214), .A2(new_n280), .A3(new_n328), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n320), .A2(G50), .ZN(new_n969));
  OAI211_X1 g0769(.A(G1), .B(new_n258), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n964), .A2(new_n967), .A3(new_n970), .ZN(G367));
  INV_X1    g0771(.A(new_n798), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n794), .B1(new_n207), .B2(new_n434), .C1(new_n230), .C2(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(new_n741), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n632), .A2(new_n633), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n677), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n649), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n626), .B2(new_n976), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G143), .A2(new_n771), .B1(new_n772), .B2(G159), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n278), .B1(new_n755), .B2(new_n832), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n747), .A2(new_n247), .B1(new_n750), .B2(new_n831), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G68), .C2(new_n758), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n766), .A2(G58), .B1(new_n767), .B2(G77), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n766), .A2(G116), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT46), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n985), .A2(new_n986), .B1(new_n772), .B2(G294), .ZN(new_n987));
  INV_X1    g0787(.A(G311), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n987), .B1(new_n986), .B2(new_n985), .C1(new_n988), .C2(new_n830), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n767), .A2(G97), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n758), .A2(G107), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n777), .A2(G303), .B1(new_n748), .B2(new_n822), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n278), .B1(new_n751), .B2(G317), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n984), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT47), .Z(new_n996));
  OAI221_X1 g0796(.A(new_n974), .B1(new_n802), .B2(new_n978), .C1(new_n996), .C2(new_n745), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT112), .Z(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n697), .B(KEYINPUT41), .Z(new_n1000));
  NAND2_X1  g0800(.A1(new_n687), .A2(new_n693), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n690), .A2(new_n693), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n686), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n737), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n590), .B(new_n600), .C1(new_n598), .C2(new_n678), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n590), .B2(new_n678), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT110), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n694), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT44), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n694), .A2(new_n1009), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT45), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n686), .A3(new_n690), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n691), .A2(new_n1014), .A3(new_n1011), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1006), .A2(new_n1016), .A3(new_n735), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1000), .B1(new_n1018), .B2(new_n735), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n740), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1009), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n1001), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n590), .B1(new_n1021), .B2(new_n557), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1023), .A2(new_n1024), .B1(new_n678), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(KEYINPUT111), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n686), .A2(new_n690), .A3(new_n1009), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1030), .A2(new_n1032), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1030), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n1033), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1031), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n999), .B1(new_n1020), .B2(new_n1040), .ZN(G387));
  OR2_X1    g0841(.A1(new_n690), .A2(new_n802), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n795), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1043), .A2(new_n699), .B1(G107), .B2(new_n207), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n972), .B1(new_n227), .B2(G45), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n699), .B(new_n477), .C1(new_n320), .C2(new_n280), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT113), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT50), .B1(new_n251), .B2(G50), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n251), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1044), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n794), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n741), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G159), .A2(new_n771), .B1(new_n772), .B2(new_n252), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n747), .A2(new_n320), .B1(new_n750), .B2(new_n832), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n278), .B1(new_n755), .B2(new_n247), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n757), .A2(new_n434), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n766), .A2(G77), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1056), .A2(new_n990), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n767), .A2(G116), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n278), .B1(new_n751), .B2(G326), .ZN(new_n1064));
  INV_X1    g0864(.A(G294), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n765), .A2(new_n1065), .B1(new_n757), .B2(new_n821), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n777), .A2(G317), .B1(new_n748), .B2(G303), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n830), .B2(new_n753), .C1(new_n988), .C2(new_n833), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1063), .B(new_n1064), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1062), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1055), .B1(new_n1075), .B2(new_n744), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1006), .A2(new_n740), .B1(new_n1042), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1003), .A2(new_n1005), .A3(new_n735), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(KEYINPUT114), .A3(new_n697), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n735), .B2(new_n1006), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT114), .B1(new_n1078), .B2(new_n697), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(G393));
  NAND3_X1  g0882(.A1(new_n1017), .A2(new_n740), .A3(new_n1016), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1009), .A2(new_n802), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT115), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n794), .B1(new_n462), .B2(new_n207), .C1(new_n235), .C2(new_n972), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT116), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n742), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n771), .A2(G150), .B1(G159), .B2(new_n777), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n766), .A2(G68), .B1(new_n767), .B2(G87), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n757), .A2(new_n280), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n278), .B1(new_n747), .B2(new_n251), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(G143), .C2(new_n751), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1092), .B(new_n1095), .C1(new_n247), .C2(new_n833), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n771), .A2(G317), .B1(G311), .B2(new_n777), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n772), .A2(G303), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n335), .B1(new_n750), .B2(new_n753), .C1(new_n747), .C2(new_n1065), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G116), .B2(new_n758), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n766), .A2(new_n822), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1101), .A3(new_n779), .A4(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1091), .A2(new_n1096), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1089), .B1(new_n744), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1085), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1083), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1017), .A2(new_n1016), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1078), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1018), .A2(new_n1109), .A3(new_n697), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT117), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT117), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1018), .A2(new_n1109), .A3(new_n1112), .A4(new_n697), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1107), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(G390));
  INV_X1    g0915(.A(KEYINPUT120), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n771), .A2(G128), .B1(G132), .B2(new_n777), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT119), .Z(new_n1118));
  NOR2_X1   g0918(.A1(new_n757), .A2(new_n781), .ZN(new_n1119));
  INV_X1    g0919(.A(G125), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT54), .B(G143), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n278), .B1(new_n750), .B2(new_n1120), .C1(new_n747), .C2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1119), .B(new_n1122), .C1(G50), .C2(new_n767), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n831), .B2(new_n833), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n766), .A2(G150), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT53), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n787), .A2(new_n837), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n278), .B1(new_n751), .B2(G294), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n462), .B2(new_n747), .C1(new_n457), .C2(new_n755), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1128), .A2(new_n1093), .A3(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G107), .A2(new_n772), .B1(new_n771), .B2(G283), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1118), .A2(new_n1127), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n741), .B1(new_n252), .B2(new_n819), .C1(new_n1133), .C2(new_n745), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n892), .A2(KEYINPUT105), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n881), .B1(new_n385), .B2(new_n867), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n886), .A2(KEYINPUT102), .A3(new_n887), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT38), .B1(new_n1138), .B2(new_n880), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n905), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT39), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n933), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1134), .B1(new_n1143), .B2(new_n791), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n952), .A2(new_n953), .A3(G330), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n897), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n914), .B1(new_n1146), .B2(new_n907), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n916), .B2(new_n934), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n678), .B(new_n896), .C1(new_n704), .C2(new_n708), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n895), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n914), .B1(new_n1152), .B2(new_n907), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n956), .A3(new_n957), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1145), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT118), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1147), .B1(new_n1142), .B2(new_n933), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n734), .A2(G330), .A3(new_n813), .A4(new_n907), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1156), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1158), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n931), .A2(KEYINPUT109), .A3(new_n892), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n955), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1161), .B1(new_n1163), .B2(new_n1153), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1149), .A2(new_n1164), .A3(KEYINPUT118), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1155), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1144), .B1(new_n1166), .B2(new_n740), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n453), .A2(G330), .A3(new_n952), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n670), .A2(new_n937), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n813), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n902), .B1(new_n815), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1145), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1146), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1152), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n952), .A2(G330), .A3(new_n813), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1158), .C1(new_n1175), .C2(new_n907), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1169), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n697), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1145), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1154), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1157), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1149), .A2(new_n1164), .A3(KEYINPUT118), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT118), .B1(new_n1149), .B2(new_n1164), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1177), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1116), .B(new_n1167), .C1(new_n1178), .C2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1177), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n697), .A3(new_n1184), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1116), .B1(new_n1191), .B2(new_n1167), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1187), .A2(new_n1192), .ZN(G378));
  INV_X1    g0993(.A(new_n1169), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1184), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n951), .A2(G330), .A3(new_n958), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n304), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n311), .A2(KEYINPUT72), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n316), .B1(new_n315), .B2(new_n305), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n268), .A2(new_n864), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT55), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n451), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n318), .B2(new_n452), .ZN(new_n1205));
  XOR2_X1   g1005(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1206));
  AND3_X1   g1006(.A1(new_n1203), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1206), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1196), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT122), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n940), .B1(new_n1163), .B2(new_n954), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n951), .A3(new_n1209), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n936), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n910), .B(new_n909), .C1(new_n1143), .C2(new_n913), .ZN(new_n1216));
  AND4_X1   g1016(.A1(G330), .A2(new_n951), .A3(new_n1209), .A4(new_n958), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1209), .B1(new_n1213), .B2(new_n951), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1211), .A2(new_n936), .A3(new_n1214), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(KEYINPUT122), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1195), .A2(new_n1215), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n698), .B1(new_n1225), .B2(new_n1195), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1221), .A2(new_n740), .A3(new_n1215), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1210), .A2(new_n791), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G97), .A2(new_n772), .B1(new_n771), .B2(G116), .ZN(new_n1230));
  INV_X1    g1030(.A(G283), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n335), .B(new_n285), .C1(new_n750), .C2(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n428), .A2(new_n755), .B1(new_n747), .B2(new_n434), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(G68), .C2(new_n758), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n767), .A2(G58), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1230), .A2(new_n1061), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT58), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n335), .A2(new_n285), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G50), .B1(new_n253), .B2(new_n285), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1236), .A2(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n777), .A2(G128), .B1(new_n748), .B2(G137), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n832), .B2(new_n757), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1121), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n766), .B2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n1120), .B2(new_n830), .C1(new_n840), .C2(new_n833), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n767), .A2(G159), .ZN(new_n1247));
  AOI211_X1 g1047(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1240), .B1(new_n1237), .B2(new_n1236), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n744), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n742), .B1(new_n247), .B2(new_n818), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1229), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1228), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1227), .A2(new_n1257), .ZN(G375));
  AND3_X1   g1058(.A1(new_n1173), .A2(new_n1169), .A3(new_n1176), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1000), .B(KEYINPUT123), .Z(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1189), .A3(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n741), .B1(G68), .B2(new_n819), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G116), .A2(new_n772), .B1(new_n771), .B2(G294), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n278), .B1(new_n751), .B2(G303), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n428), .B2(new_n747), .C1(new_n1231), .C2(new_n755), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(new_n1059), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n766), .A2(G97), .B1(new_n767), .B2(G77), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1264), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n748), .A2(G150), .B1(new_n751), .B2(G128), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n831), .B2(new_n755), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G50), .B2(new_n758), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G132), .A2(new_n771), .B1(new_n772), .B2(new_n1243), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1272), .B(new_n1273), .C1(new_n781), .C2(new_n765), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1235), .A2(new_n278), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT124), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1269), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1263), .B1(new_n1277), .B2(new_n744), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n907), .B2(new_n792), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n739), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1262), .A2(new_n1282), .ZN(G381));
  OAI211_X1 g1083(.A(new_n804), .B(new_n1077), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(G390), .A2(G381), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1167), .B1(new_n1178), .B2(new_n1185), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1256), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(G387), .A2(G384), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1285), .A2(new_n1287), .A3(new_n1288), .A4(new_n1289), .ZN(G407));
  INV_X1    g1090(.A(G213), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(G343), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1288), .A2(new_n1287), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(G407), .A2(new_n1293), .A3(G213), .ZN(G409));
  INV_X1    g1094(.A(KEYINPUT60), .ZN(new_n1295));
  OAI21_X1  g1095(.A(KEYINPUT125), .B1(new_n1260), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1259), .A2(new_n1297), .A3(KEYINPUT60), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1189), .B(new_n697), .C1(KEYINPUT60), .C2(new_n1259), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(G384), .A3(new_n1282), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1300), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n848), .B1(new_n1304), .B2(new_n1281), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(G2897), .A3(new_n1292), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1292), .A2(G2897), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1303), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1286), .A2(KEYINPUT120), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1227), .A2(new_n1311), .A3(new_n1186), .A4(new_n1257), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1195), .A2(new_n1221), .A3(new_n1215), .A4(new_n1261), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n739), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1229), .B2(new_n1254), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1286), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1312), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1292), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1310), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT63), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1320), .B2(new_n1306), .ZN(new_n1323));
  AND2_X1   g1123(.A1(G387), .A2(new_n1114), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(G387), .A2(new_n1114), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1284), .ZN(new_n1326));
  AND2_X1   g1126(.A1(G393), .A2(G396), .ZN(new_n1327));
  OAI22_X1  g1127(.A1(new_n1324), .A2(new_n1325), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  OR2_X1    g1128(.A1(G387), .A2(new_n1114), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1327), .A2(new_n1326), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(G387), .A2(new_n1114), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1328), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1292), .B1(new_n1312), .B2(new_n1317), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1306), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1321), .A2(new_n1323), .A3(new_n1333), .A4(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1338), .B1(new_n1334), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1341), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1316), .B1(G378), .B2(new_n1288), .ZN(new_n1343));
  NOR4_X1   g1143(.A1(new_n1343), .A2(KEYINPUT62), .A3(new_n1292), .A4(new_n1306), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1340), .A2(new_n1342), .A3(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1337), .B1(new_n1345), .B2(new_n1333), .ZN(G405));
  NAND2_X1  g1146(.A1(new_n1335), .A2(KEYINPUT126), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1288), .A2(new_n1286), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1312), .ZN(new_n1349));
  AOI211_X1 g1149(.A(new_n1348), .B(new_n1349), .C1(new_n1332), .C2(new_n1328), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1328), .A2(new_n1332), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1348), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1351), .B1(new_n1352), .B2(new_n1312), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1347), .B1(new_n1350), .B2(new_n1353), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1333), .B1(new_n1349), .B2(new_n1348), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1351), .A2(new_n1312), .A3(new_n1352), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1355), .A2(KEYINPUT126), .A3(new_n1335), .A4(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1354), .A2(new_n1357), .ZN(G402));
endmodule


