

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G2104), .A2(n531), .ZN(n884) );
  XNOR2_X1 U555 ( .A(KEYINPUT104), .B(KEYINPUT32), .ZN(n746) );
  AND2_X1 U556 ( .A1(n787), .A2(n786), .ZN(n521) );
  AND2_X1 U557 ( .A1(n774), .A2(n773), .ZN(n522) );
  AND2_X1 U558 ( .A1(n1021), .A2(n834), .ZN(n523) );
  XNOR2_X1 U559 ( .A(n738), .B(KEYINPUT99), .ZN(n703) );
  INV_X1 U560 ( .A(n703), .ZN(n717) );
  INV_X1 U561 ( .A(KEYINPUT28), .ZN(n693) );
  INV_X1 U562 ( .A(KEYINPUT64), .ZN(n687) );
  XNOR2_X1 U563 ( .A(n688), .B(n687), .ZN(n724) );
  INV_X1 U564 ( .A(KEYINPUT98), .ZN(n727) );
  XNOR2_X1 U565 ( .A(n728), .B(n727), .ZN(n754) );
  AND2_X1 U566 ( .A1(n754), .A2(n753), .ZN(n755) );
  AND2_X1 U567 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U568 ( .A(n747), .B(n746), .ZN(n780) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NOR2_X1 U570 ( .A1(n821), .A2(n523), .ZN(n822) );
  NOR2_X1 U571 ( .A1(G651), .A2(n623), .ZN(n648) );
  BUF_X1 U572 ( .A(n685), .Z(G160) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n524), .Z(n891) );
  NAND2_X1 U574 ( .A1(G137), .A2(n891), .ZN(n526) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U576 ( .A1(G113), .A2(n885), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U578 ( .A(n527), .B(KEYINPUT68), .ZN(n537) );
  INV_X1 U579 ( .A(G2105), .ZN(n528) );
  AND2_X4 U580 ( .A1(n528), .A2(G2104), .ZN(n892) );
  NAND2_X1 U581 ( .A1(G101), .A2(n892), .ZN(n529) );
  XOR2_X1 U582 ( .A(n529), .B(KEYINPUT23), .Z(n530) );
  XNOR2_X1 U583 ( .A(n530), .B(KEYINPUT66), .ZN(n533) );
  INV_X1 U584 ( .A(G2105), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G125), .A2(n884), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n535) );
  INV_X1 U587 ( .A(KEYINPUT67), .ZN(n534) );
  XNOR2_X1 U588 ( .A(n535), .B(n534), .ZN(n536) );
  NOR2_X2 U589 ( .A1(n537), .A2(n536), .ZN(n685) );
  NAND2_X1 U590 ( .A1(G138), .A2(n891), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G102), .A2(n892), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G126), .A2(n884), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G114), .A2(n885), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U596 ( .A1(n543), .A2(n542), .ZN(G164) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U598 ( .A(G57), .ZN(G237) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U602 ( .A1(G89), .A2(n647), .ZN(n544) );
  XOR2_X1 U603 ( .A(KEYINPUT75), .B(n544), .Z(n545) );
  XNOR2_X1 U604 ( .A(n545), .B(KEYINPUT4), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  XNOR2_X1 U606 ( .A(KEYINPUT69), .B(G651), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n623), .A2(n549), .ZN(n651) );
  NAND2_X1 U608 ( .A1(G76), .A2(n651), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n548), .B(KEYINPUT5), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n648), .A2(G51), .ZN(n552) );
  NOR2_X1 U612 ( .A1(G543), .A2(n549), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT1), .B(n550), .Z(n655) );
  NAND2_X1 U614 ( .A1(G63), .A2(n655), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT6), .B(n553), .Z(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n556), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n557), .B(KEYINPUT10), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT72), .B(n558), .Z(n930) );
  NAND2_X1 U623 ( .A1(n930), .A2(G567), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  NAND2_X1 U625 ( .A1(n655), .A2(G56), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT14), .B(n560), .Z(n566) );
  NAND2_X1 U627 ( .A1(n647), .A2(G81), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G68), .A2(n651), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT13), .B(n564), .Z(n565) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n648), .A2(G43), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n1015) );
  INV_X1 U635 ( .A(G860), .ZN(n596) );
  OR2_X1 U636 ( .A1(n1015), .A2(n596), .ZN(G153) );
  NAND2_X1 U637 ( .A1(n648), .A2(G52), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G64), .A2(n655), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G90), .A2(n647), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G77), .A2(n651), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U644 ( .A1(n575), .A2(n574), .ZN(G171) );
  INV_X1 U645 ( .A(G171), .ZN(G301) );
  NAND2_X1 U646 ( .A1(n647), .A2(G92), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G66), .A2(n655), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n648), .A2(G54), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G79), .A2(n651), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U652 ( .A(n580), .B(KEYINPUT73), .Z(n581) );
  NOR2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n583), .Z(n584) );
  XNOR2_X1 U655 ( .A(KEYINPUT74), .B(n584), .ZN(n1005) );
  INV_X1 U656 ( .A(n1005), .ZN(n709) );
  NOR2_X1 U657 ( .A1(n709), .A2(G868), .ZN(n586) );
  INV_X1 U658 ( .A(G868), .ZN(n670) );
  NOR2_X1 U659 ( .A1(n670), .A2(G301), .ZN(n585) );
  NOR2_X1 U660 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U661 ( .A1(n647), .A2(G91), .ZN(n588) );
  NAND2_X1 U662 ( .A1(G65), .A2(n655), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U664 ( .A1(G53), .A2(n648), .ZN(n589) );
  XNOR2_X1 U665 ( .A(KEYINPUT71), .B(n589), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G78), .A2(n651), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(G299) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U670 ( .A1(G286), .A2(n670), .ZN(n594) );
  NOR2_X1 U671 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n597), .A2(n1005), .ZN(n598) );
  XNOR2_X1 U674 ( .A(n598), .B(KEYINPUT76), .ZN(n599) );
  XNOR2_X1 U675 ( .A(KEYINPUT16), .B(n599), .ZN(G148) );
  NOR2_X1 U676 ( .A1(G868), .A2(n1015), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n1005), .A2(G868), .ZN(n600) );
  NOR2_X1 U678 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U679 ( .A1(n602), .A2(n601), .ZN(G282) );
  XNOR2_X1 U680 ( .A(G2100), .B(KEYINPUT79), .ZN(n613) );
  NAND2_X1 U681 ( .A1(G123), .A2(n884), .ZN(n603) );
  XNOR2_X1 U682 ( .A(n603), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G135), .A2(n891), .ZN(n605) );
  NAND2_X1 U684 ( .A1(G111), .A2(n885), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G99), .A2(n892), .ZN(n606) );
  XNOR2_X1 U687 ( .A(KEYINPUT77), .B(n606), .ZN(n607) );
  NOR2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n983) );
  XOR2_X1 U690 ( .A(G2096), .B(KEYINPUT78), .Z(n611) );
  XNOR2_X1 U691 ( .A(n983), .B(n611), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U693 ( .A1(G559), .A2(n1005), .ZN(n667) );
  XNOR2_X1 U694 ( .A(n1015), .B(n667), .ZN(n614) );
  NOR2_X1 U695 ( .A1(n614), .A2(G860), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G93), .A2(n647), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G55), .A2(n648), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n651), .A2(G80), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT80), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G67), .A2(n655), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n669) );
  XOR2_X1 U704 ( .A(n622), .B(n669), .Z(G145) );
  NAND2_X1 U705 ( .A1(n623), .A2(G87), .ZN(n624) );
  XOR2_X1 U706 ( .A(KEYINPUT82), .B(n624), .Z(n625) );
  NOR2_X1 U707 ( .A1(n655), .A2(n625), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n648), .A2(G49), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n628) );
  XNOR2_X1 U711 ( .A(KEYINPUT81), .B(n628), .ZN(n629) );
  NOR2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U713 ( .A(KEYINPUT83), .B(n631), .ZN(G288) );
  NAND2_X1 U714 ( .A1(n651), .A2(G73), .ZN(n632) );
  XNOR2_X1 U715 ( .A(n632), .B(KEYINPUT2), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n647), .A2(G86), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G61), .A2(n655), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U719 ( .A(KEYINPUT84), .B(n635), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G48), .A2(n648), .ZN(n636) );
  XNOR2_X1 U721 ( .A(KEYINPUT85), .B(n636), .ZN(n637) );
  NOR2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G88), .A2(n647), .ZN(n642) );
  NAND2_X1 U725 ( .A1(G75), .A2(n651), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n648), .A2(G50), .ZN(n644) );
  NAND2_X1 U728 ( .A1(G62), .A2(n655), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U730 ( .A1(n646), .A2(n645), .ZN(G166) );
  NAND2_X1 U731 ( .A1(G85), .A2(n647), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G47), .A2(n648), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n651), .A2(G72), .ZN(n652) );
  XOR2_X1 U735 ( .A(KEYINPUT70), .B(n652), .Z(n653) );
  NOR2_X1 U736 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U737 ( .A1(G60), .A2(n655), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n657), .A2(n656), .ZN(G290) );
  INV_X1 U739 ( .A(G299), .ZN(n696) );
  XOR2_X1 U740 ( .A(n696), .B(G288), .Z(n665) );
  XOR2_X1 U741 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n658) );
  XNOR2_X1 U742 ( .A(G305), .B(n658), .ZN(n659) );
  XOR2_X1 U743 ( .A(n659), .B(KEYINPUT19), .Z(n661) );
  XNOR2_X1 U744 ( .A(G166), .B(KEYINPUT86), .ZN(n660) );
  XNOR2_X1 U745 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U746 ( .A(n669), .B(n662), .Z(n663) );
  XNOR2_X1 U747 ( .A(n663), .B(G290), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n1015), .B(n666), .ZN(n909) );
  XNOR2_X1 U750 ( .A(n667), .B(n909), .ZN(n668) );
  NAND2_X1 U751 ( .A1(n668), .A2(G868), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U762 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G96), .A2(n679), .ZN(n842) );
  NAND2_X1 U764 ( .A1(n842), .A2(G2106), .ZN(n683) );
  NAND2_X1 U765 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U766 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G108), .A2(n681), .ZN(n843) );
  NAND2_X1 U768 ( .A1(n843), .A2(G567), .ZN(n682) );
  NAND2_X1 U769 ( .A1(n683), .A2(n682), .ZN(n863) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U771 ( .A1(n863), .A2(n684), .ZN(n841) );
  NAND2_X1 U772 ( .A1(n841), .A2(G36), .ZN(G176) );
  XNOR2_X1 U773 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  NAND2_X1 U774 ( .A1(n685), .A2(G40), .ZN(n788) );
  INV_X1 U775 ( .A(n788), .ZN(n686) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n789) );
  NAND2_X1 U777 ( .A1(n686), .A2(n789), .ZN(n688) );
  INV_X1 U778 ( .A(n724), .ZN(n738) );
  NAND2_X1 U779 ( .A1(n703), .A2(G2072), .ZN(n689) );
  XOR2_X1 U780 ( .A(KEYINPUT27), .B(n689), .Z(n691) );
  NAND2_X1 U781 ( .A1(G1956), .A2(n717), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U783 ( .A(n692), .B(KEYINPUT101), .ZN(n695) );
  NOR2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n694) );
  XNOR2_X1 U785 ( .A(n694), .B(n693), .ZN(n715) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n713) );
  AND2_X1 U787 ( .A1(n724), .A2(G1996), .ZN(n698) );
  XNOR2_X1 U788 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n697) );
  XNOR2_X1 U789 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n738), .A2(G1341), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U792 ( .A1(n1015), .A2(n701), .ZN(n708) );
  NOR2_X1 U793 ( .A1(n709), .A2(n708), .ZN(n702) );
  XOR2_X1 U794 ( .A(n702), .B(KEYINPUT102), .Z(n707) );
  NAND2_X1 U795 ( .A1(n738), .A2(G1348), .ZN(n705) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n703), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U801 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U803 ( .A(n716), .B(KEYINPUT29), .ZN(n749) );
  NOR2_X1 U804 ( .A1(G1961), .A2(n724), .ZN(n720) );
  XOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .Z(n937) );
  NOR2_X1 U806 ( .A1(n937), .A2(n717), .ZN(n718) );
  XNOR2_X1 U807 ( .A(n718), .B(KEYINPUT100), .ZN(n719) );
  NOR2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n732) );
  NOR2_X1 U809 ( .A1(G301), .A2(n732), .ZN(n748) );
  INV_X1 U810 ( .A(G286), .ZN(n721) );
  OR2_X1 U811 ( .A1(n748), .A2(n721), .ZN(n722) );
  NOR2_X1 U812 ( .A1(n749), .A2(n722), .ZN(n737) );
  NOR2_X1 U813 ( .A1(n738), .A2(G2084), .ZN(n752) );
  INV_X1 U814 ( .A(G8), .ZN(n723) );
  OR2_X2 U815 ( .A1(n724), .A2(n723), .ZN(n726) );
  INV_X1 U816 ( .A(KEYINPUT97), .ZN(n725) );
  XNOR2_X1 U817 ( .A(n726), .B(n725), .ZN(n767) );
  NOR2_X1 U818 ( .A1(n767), .A2(G1966), .ZN(n728) );
  NAND2_X1 U819 ( .A1(G8), .A2(n754), .ZN(n729) );
  NOR2_X1 U820 ( .A1(n752), .A2(n729), .ZN(n730) );
  XOR2_X1 U821 ( .A(KEYINPUT30), .B(n730), .Z(n731) );
  NOR2_X1 U822 ( .A1(G168), .A2(n731), .ZN(n734) );
  AND2_X1 U823 ( .A1(G301), .A2(n732), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U825 ( .A(n735), .B(KEYINPUT31), .ZN(n750) );
  AND2_X1 U826 ( .A1(G286), .A2(n750), .ZN(n736) );
  NOR2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n743) );
  NOR2_X1 U828 ( .A1(n738), .A2(G2090), .ZN(n740) );
  INV_X1 U829 ( .A(n767), .ZN(n776) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n767), .ZN(n739) );
  NOR2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n741), .A2(G303), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U834 ( .A(KEYINPUT103), .B(n744), .Z(n745) );
  NAND2_X1 U835 ( .A1(n745), .A2(G8), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n751) );
  OR2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n756) );
  NAND2_X1 U838 ( .A1(n752), .A2(G8), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n756), .A2(n755), .ZN(n778) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n1018) );
  AND2_X1 U841 ( .A1(n778), .A2(n1018), .ZN(n758) );
  XNOR2_X1 U842 ( .A(G1981), .B(G305), .ZN(n1007) );
  INV_X1 U843 ( .A(n1007), .ZN(n757) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n764) );
  AND2_X1 U845 ( .A1(n764), .A2(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n759), .A2(n776), .ZN(n762) );
  AND2_X1 U847 ( .A1(n760), .A2(n762), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n780), .A2(n761), .ZN(n774) );
  INV_X1 U849 ( .A(n762), .ZN(n772) );
  INV_X1 U850 ( .A(n1018), .ZN(n765) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n1023) );
  OR2_X1 U853 ( .A1(n765), .A2(n1023), .ZN(n766) );
  OR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  INV_X1 U855 ( .A(n768), .ZN(n769) );
  NOR2_X1 U856 ( .A1(KEYINPUT33), .A2(n769), .ZN(n770) );
  OR2_X1 U857 ( .A1(n1007), .A2(n770), .ZN(n771) );
  OR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XNOR2_X1 U860 ( .A(n775), .B(KEYINPUT24), .ZN(n777) );
  AND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n782) );
  OR2_X1 U862 ( .A1(n782), .A2(n767), .ZN(n785) );
  AND2_X1 U863 ( .A1(n778), .A2(n785), .ZN(n779) );
  NAND2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n787) );
  INV_X1 U865 ( .A(G2090), .ZN(n990) );
  NAND2_X1 U866 ( .A1(G8), .A2(n990), .ZN(n781) );
  NOR2_X1 U867 ( .A1(n781), .A2(G303), .ZN(n783) );
  OR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n522), .A2(n521), .ZN(n823) );
  NOR2_X1 U871 ( .A1(n789), .A2(n788), .ZN(n834) );
  XNOR2_X1 U872 ( .A(KEYINPUT93), .B(KEYINPUT36), .ZN(n801) );
  NAND2_X1 U873 ( .A1(G140), .A2(n891), .ZN(n791) );
  NAND2_X1 U874 ( .A1(G104), .A2(n892), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U876 ( .A(n792), .B(KEYINPUT34), .ZN(n793) );
  XNOR2_X1 U877 ( .A(n793), .B(KEYINPUT91), .ZN(n799) );
  XNOR2_X1 U878 ( .A(KEYINPUT92), .B(KEYINPUT35), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G128), .A2(n884), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G116), .A2(n885), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U882 ( .A(n797), .B(n796), .ZN(n798) );
  NAND2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U884 ( .A(n801), .B(n800), .ZN(n898) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n832) );
  NOR2_X1 U886 ( .A1(n898), .A2(n832), .ZN(n981) );
  NAND2_X1 U887 ( .A1(n834), .A2(n981), .ZN(n830) );
  NAND2_X1 U888 ( .A1(G129), .A2(n884), .ZN(n803) );
  NAND2_X1 U889 ( .A1(G117), .A2(n885), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U891 ( .A1(n892), .A2(G105), .ZN(n804) );
  XOR2_X1 U892 ( .A(KEYINPUT38), .B(n804), .Z(n805) );
  NOR2_X1 U893 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n891), .A2(G141), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n808), .A2(n807), .ZN(n880) );
  NAND2_X1 U896 ( .A1(G1996), .A2(n880), .ZN(n809) );
  XNOR2_X1 U897 ( .A(n809), .B(KEYINPUT94), .ZN(n817) );
  NAND2_X1 U898 ( .A1(G119), .A2(n884), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G107), .A2(n885), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n811), .A2(n810), .ZN(n815) );
  NAND2_X1 U901 ( .A1(G131), .A2(n891), .ZN(n813) );
  NAND2_X1 U902 ( .A1(G95), .A2(n892), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n901) );
  NAND2_X1 U905 ( .A1(G1991), .A2(n901), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U907 ( .A(KEYINPUT95), .B(n818), .Z(n989) );
  NAND2_X1 U908 ( .A1(n989), .A2(n834), .ZN(n824) );
  NAND2_X1 U909 ( .A1(n830), .A2(n824), .ZN(n819) );
  XNOR2_X1 U910 ( .A(n819), .B(KEYINPUT96), .ZN(n821) );
  XNOR2_X1 U911 ( .A(G1986), .B(KEYINPUT90), .ZN(n820) );
  XNOR2_X1 U912 ( .A(n820), .B(G290), .ZN(n1021) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n837) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n880), .ZN(n992) );
  INV_X1 U915 ( .A(n824), .ZN(n827) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n901), .ZN(n986) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n986), .A2(n825), .ZN(n826) );
  NOR2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U920 ( .A1(n992), .A2(n828), .ZN(n829) );
  XNOR2_X1 U921 ( .A(n829), .B(KEYINPUT39), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U923 ( .A1(n898), .A2(n832), .ZN(n980) );
  NAND2_X1 U924 ( .A1(n833), .A2(n980), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U926 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U927 ( .A(n838), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n930), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U930 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U932 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XOR2_X1 U939 ( .A(G2096), .B(G2100), .Z(n845) );
  XNOR2_X1 U940 ( .A(KEYINPUT42), .B(G2678), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n849) );
  XNOR2_X1 U942 ( .A(KEYINPUT43), .B(n990), .ZN(n847) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U945 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U948 ( .A(KEYINPUT107), .B(G1981), .Z(n853) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1961), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U951 ( .A(n854), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U954 ( .A(G1976), .B(G1971), .Z(n858) );
  XNOR2_X1 U955 ( .A(G1956), .B(G1966), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U958 ( .A(KEYINPUT106), .B(G2474), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(G229) );
  INV_X1 U960 ( .A(n863), .ZN(G319) );
  NAND2_X1 U961 ( .A1(G124), .A2(n884), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n864), .B(KEYINPUT108), .ZN(n865) );
  XNOR2_X1 U963 ( .A(KEYINPUT44), .B(n865), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G100), .A2(n892), .ZN(n866) );
  XOR2_X1 U965 ( .A(KEYINPUT109), .B(n866), .Z(n867) );
  NAND2_X1 U966 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G136), .A2(n891), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G112), .A2(n885), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U970 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G130), .A2(n884), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G118), .A2(n885), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G142), .A2(n891), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G106), .A2(n892), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n883) );
  XNOR2_X1 U979 ( .A(G160), .B(n880), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n881), .B(n983), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n900) );
  XNOR2_X1 U982 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n890) );
  NAND2_X1 U983 ( .A1(G127), .A2(n884), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G115), .A2(n885), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n888), .B(KEYINPUT47), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n896) );
  NAND2_X1 U988 ( .A1(G139), .A2(n891), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G103), .A2(n892), .ZN(n893) );
  NAND2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n895) );
  NOR2_X1 U991 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U992 ( .A(KEYINPUT112), .B(n897), .Z(n976) );
  XNOR2_X1 U993 ( .A(n898), .B(n976), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n906) );
  XNOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n901), .B(G162), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U998 ( .A(G164), .B(n904), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n907), .ZN(n908) );
  XOR2_X1 U1001 ( .A(KEYINPUT113), .B(n908), .Z(G395) );
  XOR2_X1 U1002 ( .A(G301), .B(n1005), .Z(n910) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1004 ( .A(G286), .B(n911), .Z(n912) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n912), .ZN(G397) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n926) );
  XOR2_X1 U1009 ( .A(KEYINPUT105), .B(G2446), .Z(n916) );
  XNOR2_X1 U1010 ( .A(G2435), .B(G2438), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n923) );
  XOR2_X1 U1012 ( .A(G2451), .B(G2430), .Z(n918) );
  XNOR2_X1 U1013 ( .A(G2454), .B(G2427), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1015 ( .A(n919), .B(G2443), .Z(n921) );
  XNOR2_X1 U1016 ( .A(G1348), .B(G1341), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n924), .A2(G14), .ZN(n929) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n929), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n929), .ZN(G401) );
  INV_X1 U1027 ( .A(n930), .ZN(G223) );
  XNOR2_X1 U1028 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1038) );
  XOR2_X1 U1029 ( .A(G35), .B(G2090), .Z(n933) );
  XOR2_X1 U1030 ( .A(G2084), .B(G34), .Z(n931) );
  XNOR2_X1 U1031 ( .A(KEYINPUT54), .B(n931), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n947) );
  XOR2_X1 U1033 ( .A(G2067), .B(G26), .Z(n934) );
  NAND2_X1 U1034 ( .A1(n934), .A2(G28), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(G1996), .B(G32), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(G1991), .B(G25), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(G27), .B(n937), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(KEYINPUT53), .B(n944), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT118), .B(n945), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1046 ( .A(KEYINPUT55), .B(n948), .Z(n949) );
  NOR2_X1 U1047 ( .A1(G29), .A2(n949), .ZN(n1036) );
  XOR2_X1 U1048 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n956) );
  XNOR2_X1 U1049 ( .A(G1986), .B(G24), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(G22), .B(G1971), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(G1976), .B(KEYINPUT123), .ZN(n952) );
  XNOR2_X1 U1053 ( .A(n952), .B(G23), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(n956), .B(n955), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(G1961), .B(G5), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(G21), .B(G1966), .ZN(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n972) );
  XOR2_X1 U1060 ( .A(G4), .B(KEYINPUT122), .Z(n962) );
  XNOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT59), .ZN(n961) );
  XNOR2_X1 U1062 ( .A(n962), .B(n961), .ZN(n965) );
  XOR2_X1 U1063 ( .A(KEYINPUT121), .B(G1341), .Z(n963) );
  XNOR2_X1 U1064 ( .A(G19), .B(n963), .ZN(n964) );
  NOR2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(G1956), .B(G20), .ZN(n967) );
  XNOR2_X1 U1067 ( .A(G6), .B(G1981), .ZN(n966) );
  NOR2_X1 U1068 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1070 ( .A(KEYINPUT60), .B(n970), .ZN(n971) );
  NOR2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1072 ( .A(KEYINPUT61), .B(n973), .Z(n974) );
  NOR2_X1 U1073 ( .A1(G16), .A2(n974), .ZN(n1033) );
  XOR2_X1 U1074 ( .A(G164), .B(G2078), .Z(n975) );
  XNOR2_X1 U1075 ( .A(KEYINPUT116), .B(n975), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(n976), .B(G2072), .ZN(n977) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1078 ( .A(KEYINPUT50), .B(n979), .Z(n1000) );
  INV_X1 U1079 ( .A(n980), .ZN(n982) );
  NOR2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(G160), .B(G2084), .ZN(n984) );
  NAND2_X1 U1082 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n997) );
  INV_X1 U1085 ( .A(n989), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n990), .B(G162), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n993), .Z(n994) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT115), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1093 ( .A(KEYINPUT52), .B(n1001), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(KEYINPUT55), .A2(n1002), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(n1003), .B(KEYINPUT117), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1097 ( .A(G16), .B(KEYINPUT56), .ZN(n1029) );
  XOR2_X1 U1098 ( .A(G1348), .B(n1005), .Z(n1011) );
  XOR2_X1 U1099 ( .A(G1966), .B(G168), .Z(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1101 ( .A(KEYINPUT57), .B(n1008), .Z(n1009) );
  XNOR2_X1 U1102 ( .A(KEYINPUT119), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1027) );
  XOR2_X1 U1104 ( .A(G299), .B(G1956), .Z(n1012) );
  XNOR2_X1 U1105 ( .A(n1012), .B(KEYINPUT120), .ZN(n1014) );
  NAND2_X1 U1106 ( .A1(G1971), .A2(G303), .ZN(n1013) );
  NAND2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1108 ( .A(G1341), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NAND2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(G1961), .B(G301), .ZN(n1020) );
  NOR2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(G11), .ZN(n1035) );
  NOR2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1121 ( .A(n1038), .B(n1037), .ZN(n1039) );
  XOR2_X1 U1122 ( .A(KEYINPUT125), .B(n1039), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

