//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT75), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n190), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n195), .A2(new_n197), .A3(new_n198), .A4(G128), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT77), .B1(new_n204), .B2(G104), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT77), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G107), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n207), .B2(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(KEYINPUT3), .A3(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n207), .A2(G107), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n204), .A2(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n203), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n209), .A2(new_n213), .A3(new_n214), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n214), .B1(new_n209), .B2(new_n213), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n213), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n224), .A3(G101), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n195), .A2(new_n197), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G128), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n202), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n221), .B1(new_n225), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n195), .A2(new_n197), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT64), .B(G128), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n198), .B1(G143), .B2(new_n194), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n235), .B1(new_n239), .B2(new_n199), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT79), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n215), .A2(new_n241), .A3(new_n218), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n215), .B2(new_n218), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT80), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT80), .B(new_n240), .C1(new_n242), .C2(new_n243), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n234), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(G137), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(G137), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n251), .A2(new_n254), .A3(new_n257), .A4(new_n252), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n248), .A2(new_n260), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n259), .B(new_n234), .C1(new_n246), .C2(new_n247), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n193), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n193), .B1(new_n248), .B2(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n215), .A2(new_n218), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n239), .A2(new_n199), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n219), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n259), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  AOI211_X1 g088(.A(G469), .B(G902), .C1(new_n263), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n234), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n265), .A2(KEYINPUT79), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n215), .A2(new_n241), .A3(new_n218), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT80), .B1(new_n279), .B2(new_n240), .ZN(new_n280));
  INV_X1    g094(.A(new_n247), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n260), .B(new_n276), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n273), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n193), .B(KEYINPUT76), .Z(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n259), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n264), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n288), .A3(G469), .ZN(new_n289));
  NAND2_X1  g103(.A1(G469), .A2(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n188), .B1(new_n275), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n191), .A2(G952), .ZN(new_n293));
  NAND2_X1  g107(.A1(G234), .A2(G237), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(G902), .A3(G953), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT21), .B(G898), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g117(.A1(G116), .A2(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(G116), .A2(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT2), .A2(G113), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(KEYINPUT2), .A2(G113), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n304), .B(new_n305), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n310));
  INV_X1    g124(.A(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(G116), .A2(G119), .ZN(new_n313));
  NOR2_X1   g127(.A1(G116), .A2(G119), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n312), .B(new_n306), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n309), .A2(new_n315), .A3(KEYINPUT65), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT65), .B1(new_n309), .B2(new_n315), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n227), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT81), .B1(new_n318), .B2(new_n225), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n309), .A2(new_n315), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n309), .A2(new_n315), .A3(KEYINPUT65), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n226), .A2(G101), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n324), .A2(new_n326), .A3(new_n327), .A4(new_n227), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n329));
  INV_X1    g143(.A(G119), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G116), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n331), .A2(KEYINPUT82), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(KEYINPUT82), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n304), .A2(new_n305), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n311), .B1(new_n335), .B2(KEYINPUT5), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n307), .A2(new_n308), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n334), .A2(new_n336), .B1(new_n337), .B2(new_n335), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n242), .B2(new_n243), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n319), .A2(new_n328), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G122), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n319), .A2(new_n341), .A3(new_n328), .A4(new_n339), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(KEYINPUT6), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n231), .A2(G125), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n267), .B2(G125), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n191), .A2(G224), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n347), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n340), .A2(new_n351), .A3(new_n342), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n347), .B1(KEYINPUT86), .B2(new_n349), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n348), .A2(KEYINPUT7), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n347), .A2(KEYINPUT86), .A3(KEYINPUT7), .A4(new_n348), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(new_n344), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n266), .B1(new_n338), .B2(KEYINPUT84), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n338), .A2(KEYINPUT84), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n341), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n363), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(new_n360), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT85), .B1(new_n338), .B2(new_n266), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n364), .B(new_n366), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n359), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G210), .B1(G237), .B2(G902), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n353), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n353), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n303), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n237), .A2(G143), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n196), .A2(G128), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT13), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G134), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n250), .A3(new_n378), .ZN(new_n382));
  XNOR2_X1  g196(.A(G116), .B(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n204), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n204), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G122), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n204), .B1(new_n390), .B2(KEYINPUT14), .ZN(new_n391));
  AOI22_X1  g205(.A1(KEYINPUT94), .A2(new_n386), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(KEYINPUT94), .B2(new_n386), .ZN(new_n393));
  INV_X1    g207(.A(new_n382), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n250), .B1(new_n376), .B2(new_n378), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n385), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G217), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n187), .A2(new_n398), .A3(G953), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n385), .B(new_n399), .C1(new_n393), .C2(new_n396), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n397), .A2(new_n402), .A3(new_n400), .ZN(new_n405));
  INV_X1    g219(.A(G902), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT15), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n407), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G125), .ZN(new_n413));
  INV_X1    g227(.A(G125), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G140), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT16), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT71), .ZN(new_n417));
  XNOR2_X1  g231(.A(G125), .B(G140), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT71), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT16), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n414), .A2(KEYINPUT16), .A3(G140), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AND4_X1   g236(.A1(G146), .A2(new_n417), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n416), .B2(KEYINPUT71), .ZN(new_n424));
  AOI21_X1  g238(.A(G146), .B1(new_n424), .B2(new_n420), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT90), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n420), .A3(new_n422), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n194), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT90), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n424), .A2(G146), .A3(new_n420), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(G237), .A2(G953), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(G143), .A3(G214), .ZN(new_n433));
  AOI21_X1  g247(.A(G143), .B1(new_n432), .B2(G214), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  INV_X1    g250(.A(G237), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n191), .A3(G214), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n196), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n432), .A2(G143), .A3(G214), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n257), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n435), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n440), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT17), .A3(G131), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n426), .A2(new_n431), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT93), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n413), .A2(new_n415), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G146), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n418), .A2(new_n194), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(KEYINPUT18), .A2(G131), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n433), .B2(new_n434), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n439), .A2(new_n440), .A3(new_n452), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n446), .A2(new_n447), .A3(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G113), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT89), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n207), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n446), .A2(new_n458), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(KEYINPUT93), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n446), .A2(new_n463), .A3(new_n458), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT91), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT91), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n446), .A2(new_n468), .A3(new_n463), .A4(new_n458), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n459), .A2(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G475), .B1(new_n470), .B2(G902), .ZN(new_n471));
  NOR2_X1   g285(.A1(G475), .A2(G902), .ZN(new_n472));
  AND2_X1   g286(.A1(KEYINPUT92), .A2(KEYINPUT20), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n467), .A2(new_n469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n435), .A2(new_n441), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n448), .B(KEYINPUT19), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(new_n430), .C1(G146), .C2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n463), .B1(new_n479), .B2(new_n458), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(KEYINPUT92), .A2(KEYINPUT20), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n458), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n467), .A2(new_n469), .B1(new_n484), .B2(new_n462), .ZN(new_n485));
  INV_X1    g299(.A(new_n472), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n411), .A2(new_n471), .A3(new_n481), .A4(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n292), .A2(new_n375), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT32), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n316), .A2(new_n317), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n259), .A2(new_n232), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n250), .A2(G137), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n253), .A2(G134), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n258), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n267), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n258), .A2(new_n495), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n239), .B2(new_n199), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n231), .B1(new_n258), .B2(new_n256), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n324), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n498), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT67), .B1(new_n505), .B2(KEYINPUT28), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT67), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n507), .B(new_n499), .C1(new_n504), .C2(new_n498), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n500), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n437), .A2(new_n191), .A3(G210), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT27), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT27), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n432), .A2(new_n512), .A3(G210), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT26), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT26), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n515), .A2(G101), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G101), .B1(new_n515), .B2(new_n517), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n502), .B2(new_n503), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n492), .A2(new_n497), .A3(KEYINPUT30), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n324), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT31), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(KEYINPUT66), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n518), .A2(new_n519), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n528), .A3(new_n498), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT66), .A3(new_n526), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(KEYINPUT66), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n525), .A2(new_n528), .A3(new_n498), .A4(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n509), .A2(new_n521), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G472), .A2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n490), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n491), .A2(new_n492), .A3(new_n497), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n492), .A2(new_n497), .B1(new_n322), .B2(new_n323), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT28), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n507), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n505), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n520), .B1(new_n542), .B2(new_n500), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n529), .B(new_n531), .ZN(new_n544));
  OAI211_X1 g358(.A(KEYINPUT32), .B(new_n534), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n500), .A2(new_n520), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n505), .B2(KEYINPUT28), .ZN(new_n549));
  AOI21_X1  g363(.A(G902), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n546), .B1(new_n540), .B2(new_n541), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n525), .A2(new_n498), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n521), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n548), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n550), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G472), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n536), .A2(new_n545), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT68), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT68), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n536), .A2(new_n545), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(G217), .A2(G902), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n398), .B2(G234), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT69), .Z(new_n564));
  NOR2_X1   g378(.A1(new_n200), .A2(G119), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n330), .B2(G128), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT64), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G128), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n571), .A3(G119), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n566), .B(new_n568), .C1(new_n572), .C2(new_n567), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(G110), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n565), .B1(new_n237), .B2(G119), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT24), .B(G110), .Z(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n430), .B(new_n450), .C1(new_n574), .C2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n423), .A2(new_n425), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(G110), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n575), .B2(new_n576), .ZN(new_n582));
  AND4_X1   g396(.A1(new_n581), .A2(new_n576), .A3(new_n572), .A4(new_n566), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n578), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT22), .B(G137), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT72), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n576), .A2(new_n572), .A3(new_n566), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT70), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n575), .A2(new_n581), .A3(new_n576), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(new_n580), .C1(new_n423), .C2(new_n425), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n578), .A3(new_n589), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT25), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n564), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n596), .A2(new_n578), .A3(new_n589), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n589), .B1(new_n596), .B2(new_n578), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n406), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT25), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT73), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n598), .A2(new_n599), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(KEYINPUT25), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT73), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n564), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n564), .A2(G902), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n601), .B2(new_n602), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n605), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT74), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n605), .A2(KEYINPUT74), .A3(new_n609), .A4(new_n611), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n489), .A2(new_n561), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  NAND3_X1  g432(.A1(new_n471), .A2(new_n481), .A3(new_n487), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n353), .A2(new_n371), .A3(new_n372), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n301), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n373), .A2(new_n374), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n623), .B2(new_n621), .ZN(new_n624));
  INV_X1    g438(.A(new_n300), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n404), .A2(new_n405), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n401), .A2(KEYINPUT33), .A3(new_n403), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(G478), .A3(new_n406), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n407), .A2(new_n408), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND4_X1   g445(.A1(new_n619), .A2(new_n624), .A3(new_n625), .A4(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n533), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n534), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n533), .B2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n292), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n616), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  AOI21_X1  g455(.A(new_n302), .B1(new_n373), .B2(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n353), .A2(new_n371), .ZN(new_n643));
  INV_X1    g457(.A(new_n372), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n621), .A3(new_n620), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n407), .B(new_n409), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n648), .A2(new_n471), .A3(new_n481), .A4(new_n487), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n647), .A2(new_n300), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n638), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n589), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n585), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n610), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n605), .A2(new_n609), .A3(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n657), .A2(new_n634), .A3(new_n635), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n489), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  AND3_X1   g475(.A1(new_n642), .A2(new_n646), .A3(new_n657), .ZN(new_n662));
  INV_X1    g476(.A(new_n188), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n283), .A2(new_n284), .B1(new_n264), .B2(new_n287), .ZN(new_n664));
  OAI21_X1  g478(.A(G469), .B1(new_n664), .B2(G902), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n263), .A2(new_n274), .ZN(new_n666));
  INV_X1    g480(.A(G469), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n406), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n663), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n296), .B1(new_n298), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n649), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n662), .A2(new_n561), .A3(new_n669), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XOR2_X1   g488(.A(new_n671), .B(KEYINPUT39), .Z(new_n675));
  NAND2_X1  g489(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT98), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n676), .A2(KEYINPUT98), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n676), .A2(KEYINPUT98), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(KEYINPUT40), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT97), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n623), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT97), .B1(new_n373), .B2(new_n374), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n684), .A2(new_n685), .A3(KEYINPUT38), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT38), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n471), .A2(new_n481), .A3(new_n487), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n411), .ZN(new_n690));
  INV_X1    g504(.A(new_n552), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n521), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n406), .B1(new_n505), .B2(new_n520), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n536), .A2(new_n545), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n657), .A2(new_n302), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n690), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n679), .A2(new_n682), .A3(new_n688), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  INV_X1    g513(.A(new_n671), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n619), .A2(new_n631), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n662), .A2(new_n561), .A3(new_n669), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  AND2_X1   g517(.A1(new_n561), .A2(new_n616), .ZN(new_n704));
  INV_X1    g518(.A(new_n193), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n282), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n273), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n287), .B2(new_n282), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n406), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT99), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n668), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(KEYINPUT99), .A3(G469), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n663), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n632), .A2(new_n704), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND3_X1  g532(.A1(new_n704), .A2(new_n650), .A3(new_n715), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT100), .B(G116), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G18));
  NAND3_X1  g535(.A1(new_n642), .A2(new_n646), .A3(new_n657), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n560), .B2(new_n558), .ZN(new_n723));
  INV_X1    g537(.A(new_n488), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n663), .B(new_n300), .C1(new_n713), .C2(new_n714), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NAND2_X1  g541(.A1(new_n530), .A2(new_n532), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n539), .A2(new_n500), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n521), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n535), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n509), .A2(new_n521), .ZN(new_n732));
  AOI21_X1  g546(.A(G902), .B1(new_n732), .B2(new_n728), .ZN(new_n733));
  INV_X1    g547(.A(G472), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT101), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT101), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(G472), .C1(new_n533), .C2(G902), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n731), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n612), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n624), .A2(new_n690), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n713), .A2(new_n714), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n188), .A3(new_n625), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT102), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  AOI211_X1 g558(.A(new_n731), .B(new_n612), .C1(new_n735), .C2(new_n737), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n648), .A2(new_n642), .A3(new_n646), .A4(new_n619), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n725), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  AND3_X1   g563(.A1(new_n741), .A2(new_n624), .A3(new_n188), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n701), .A2(new_n657), .A3(new_n738), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n741), .A2(new_n624), .A3(new_n188), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n701), .A2(new_n657), .A3(new_n738), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT103), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  NAND3_X1  g572(.A1(new_n645), .A2(new_n620), .A3(new_n301), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n292), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n561), .A2(new_n616), .A3(new_n701), .A4(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n545), .B(KEYINPUT105), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n536), .A2(new_n556), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n612), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(KEYINPUT42), .A3(new_n701), .A4(new_n760), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G131), .ZN(G33));
  AND3_X1   g583(.A1(new_n561), .A2(new_n616), .A3(new_n760), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n672), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND2_X1  g586(.A1(new_n689), .A2(new_n631), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n636), .A2(new_n657), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(KEYINPUT44), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n759), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n664), .A2(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n664), .A2(KEYINPUT45), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(G469), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n290), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT46), .B1(new_n782), .B2(new_n290), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n668), .B(new_n783), .C1(new_n784), .C2(KEYINPUT106), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(KEYINPUT106), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n663), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n779), .A2(new_n788), .A3(new_n675), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  INV_X1    g607(.A(new_n787), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n188), .B1(new_n794), .B2(new_n785), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n797), .B(new_n188), .C1(new_n785), .C2(new_n794), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n561), .A2(new_n616), .A3(new_n759), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n701), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT107), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n412), .ZN(G42));
  NAND2_X1  g616(.A1(new_n774), .A2(new_n775), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n745), .A2(new_n296), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n688), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n302), .A3(new_n806), .A4(new_n715), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT50), .Z(new_n808));
  INV_X1    g622(.A(new_n695), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n759), .A2(new_n295), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n715), .A2(new_n616), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n619), .A3(new_n631), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n805), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n796), .A2(new_n798), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n741), .A2(new_n663), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n759), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n715), .A2(new_n774), .A3(new_n775), .A4(new_n810), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT114), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n735), .A2(new_n737), .ZN(new_n822));
  INV_X1    g636(.A(new_n731), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n822), .A2(new_n657), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n814), .A2(new_n819), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n814), .A2(new_n819), .A3(KEYINPUT51), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n821), .A2(new_n766), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT48), .Z(new_n831));
  NAND2_X1  g645(.A1(new_n619), .A2(new_n631), .ZN(new_n832));
  OAI221_X1 g646(.A(new_n293), .B1(new_n832), .B2(new_n811), .C1(new_n815), .C2(new_n754), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n829), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n657), .A2(new_n671), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT112), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n669), .A3(new_n695), .A4(new_n746), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n723), .B(new_n669), .C1(new_n672), .C2(new_n701), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT103), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n757), .A2(KEYINPUT52), .A3(new_n838), .A4(new_n839), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n704), .B(new_n715), .C1(new_n632), .C2(new_n650), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n748), .A2(new_n726), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT110), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n748), .A2(new_n847), .A3(KEYINPUT110), .A4(new_n726), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n778), .A2(new_n669), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT111), .B1(new_n755), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n824), .A2(new_n854), .A3(new_n701), .A4(new_n760), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n657), .A2(new_n700), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n852), .A2(new_n488), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n853), .A2(new_n855), .B1(new_n561), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n375), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n832), .A2(new_n649), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n616), .A2(new_n637), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n617), .A2(new_n861), .A3(new_n659), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n858), .A2(new_n768), .A3(new_n771), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n846), .A2(new_n850), .A3(new_n851), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n850), .A2(new_n851), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n863), .B1(new_n844), .B2(new_n845), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT53), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT54), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n748), .A2(new_n847), .A3(KEYINPUT53), .A4(new_n726), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n863), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n846), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT113), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n846), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT54), .B1(new_n865), .B2(new_n866), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n835), .A2(new_n881), .B1(G952), .B2(G953), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT49), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n741), .A2(new_n883), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n773), .A2(new_n612), .A3(new_n663), .A4(new_n302), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n884), .B1(new_n886), .B2(KEYINPUT108), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(KEYINPUT108), .B2(new_n886), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT109), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n695), .B1(new_n741), .B2(new_n883), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n806), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n882), .A2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n191), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n865), .A2(new_n866), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n878), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(G210), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n406), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n345), .A2(new_n352), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT115), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n350), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n894), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n903), .ZN(new_n905));
  AOI211_X1 g719(.A(KEYINPUT56), .B(new_n905), .C1(new_n896), .C2(new_n898), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT116), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n875), .A2(new_n877), .B1(new_n865), .B2(new_n866), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n908), .A2(new_n897), .A3(new_n406), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(KEYINPUT56), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT116), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n899), .A2(new_n903), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n894), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n907), .A2(new_n913), .ZN(G51));
  XOR2_X1   g728(.A(new_n290), .B(KEYINPUT57), .Z(new_n915));
  AND3_X1   g729(.A1(new_n846), .A2(new_n876), .A3(new_n873), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n876), .B1(new_n846), .B2(new_n873), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n918), .B2(new_n870), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT117), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT117), .B1(new_n878), .B2(new_n879), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n666), .ZN(new_n924));
  OR3_X1    g738(.A1(new_n908), .A2(new_n406), .A3(new_n782), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n893), .B1(new_n924), .B2(new_n925), .ZN(G54));
  NAND4_X1  g740(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n485), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n485), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n893), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n871), .B2(new_n880), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n627), .A2(new_n628), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n894), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n921), .A2(new_n922), .ZN(new_n936));
  INV_X1    g750(.A(new_n934), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n932), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(G63));
  XNOR2_X1  g753(.A(new_n562), .B(KEYINPUT60), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n597), .B(new_n591), .C1(new_n908), .C2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n655), .B(new_n942), .C1(new_n918), .C2(new_n870), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n894), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT118), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n945), .A3(new_n894), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(KEYINPUT61), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n878), .B2(new_n895), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n893), .B1(new_n948), .B2(new_n655), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n949), .B(new_n941), .C1(new_n945), .C2(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n947), .A2(new_n951), .ZN(G66));
  INV_X1    g766(.A(new_n299), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n953), .A2(G224), .A3(G953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n868), .A2(new_n862), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT119), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT119), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n868), .A2(new_n957), .A3(new_n862), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n954), .B1(new_n959), .B2(new_n191), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n901), .B1(G898), .B2(new_n191), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G69));
  AOI21_X1  g776(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT124), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n523), .A2(new_n524), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n478), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n860), .B(KEYINPUT120), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n675), .A3(new_n770), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n800), .A2(new_n792), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n673), .A2(new_n702), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n753), .B2(new_n756), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n698), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n973), .A2(new_n698), .A3(KEYINPUT62), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n971), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n968), .B1(new_n978), .B2(G953), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT121), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n792), .A2(new_n973), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT122), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT122), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n792), .A2(new_n983), .A3(new_n973), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n768), .A2(new_n771), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n788), .A2(new_n675), .A3(new_n746), .A4(new_n766), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n800), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n985), .A2(new_n991), .A3(new_n191), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n968), .B1(G900), .B2(G953), .ZN(new_n993));
  AOI22_X1  g807(.A1(new_n979), .A2(new_n980), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(KEYINPUT121), .B(new_n968), .C1(new_n978), .C2(G953), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n965), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n971), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n976), .A2(new_n977), .ZN(new_n998));
  AOI21_X1  g812(.A(G953), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n980), .B1(new_n999), .B2(new_n967), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n992), .A2(new_n993), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1000), .A2(new_n1001), .A3(new_n995), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1002), .A2(KEYINPUT124), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n964), .B1(new_n996), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n994), .A2(new_n965), .A3(new_n995), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(KEYINPUT124), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n963), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1004), .A2(new_n1007), .ZN(G72));
  NAND2_X1  g822(.A1(new_n691), .A2(new_n521), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT63), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n692), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1009), .B(new_n1013), .C1(new_n867), .C2(new_n870), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1012), .B1(new_n959), .B2(new_n978), .ZN(new_n1015));
  INV_X1    g829(.A(new_n692), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n956), .A2(new_n958), .A3(new_n985), .A4(new_n991), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1019), .B1(new_n1020), .B2(new_n1011), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT126), .ZN(new_n1022));
  OR3_X1    g836(.A1(new_n1021), .A2(new_n1022), .A3(new_n893), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1022), .B1(new_n1021), .B2(new_n893), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1017), .B1(new_n1023), .B2(new_n1024), .ZN(G57));
endmodule


