//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n202), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n217), .B(new_n220), .C1(new_n223), .C2(new_n225), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  XNOR2_X1  g0043(.A(KEYINPUT3), .B(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n244), .A2(G222), .A3(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n244), .A2(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G223), .ZN(new_n249));
  OAI221_X1 g0049(.A(new_n246), .B1(new_n247), .B2(new_n244), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  AND2_X1   g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(new_n221), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(new_n251), .B2(new_n221), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n256), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n255), .A2(G274), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G41), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n255), .A2(new_n257), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n253), .B(new_n266), .C1(new_n209), .C2(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n271), .A2(G179), .ZN(new_n272));
  OAI21_X1  g0072(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n273));
  INV_X1    g0073(.A(G150), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n222), .A2(G33), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n273), .B1(new_n274), .B2(new_n276), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT69), .B1(new_n205), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT69), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(new_n221), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n279), .A2(new_n284), .B1(new_n208), .B2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n281), .A2(new_n283), .A3(new_n221), .A4(new_n285), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n268), .A2(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G50), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n271), .A2(new_n293), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n272), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n271), .A2(G200), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n296), .B1(new_n297), .B2(new_n292), .C1(new_n298), .C2(new_n271), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT9), .B1(new_n287), .B2(new_n291), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT72), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n299), .A2(KEYINPUT10), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n295), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n244), .A2(G232), .A3(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n244), .A2(new_n245), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n209), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n252), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n267), .A2(G238), .A3(new_n269), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n266), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT13), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n309), .A2(new_n313), .A3(new_n266), .A4(new_n310), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT14), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(G169), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(G179), .A3(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n315), .B2(G169), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n275), .A2(G50), .B1(G20), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n247), .B2(new_n278), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n323), .A2(new_n284), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT11), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n285), .A2(G68), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n326), .A2(KEYINPUT73), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT12), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n326), .B2(KEYINPUT73), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n329), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n325), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n289), .A2(G68), .A3(new_n290), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n324), .B2(KEYINPUT11), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n319), .A2(new_n320), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n315), .A2(G200), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n332), .A2(new_n334), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n336), .B(new_n337), .C1(new_n298), .C2(new_n315), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G33), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n341), .A2(new_n343), .A3(G226), .A4(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n341), .A2(new_n343), .A3(G223), .A4(new_n245), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G87), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n347), .A2(new_n252), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n255), .A2(new_n257), .A3(G232), .A4(new_n269), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n255), .A2(G274), .A3(new_n257), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n260), .A2(new_n262), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n268), .B1(new_n351), .B2(G45), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(G169), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n347), .A2(new_n252), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n266), .A2(new_n355), .A3(G179), .A4(new_n349), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n244), .A2(new_n360), .A3(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n341), .A2(new_n343), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n362), .B2(new_n222), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n275), .A2(G159), .ZN(new_n365));
  INV_X1    g0165(.A(G58), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n321), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n367), .B2(new_n201), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n364), .A2(KEYINPUT16), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n360), .B1(new_n244), .B2(G20), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n362), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n321), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n365), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n375), .A3(new_n284), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n277), .B1(new_n268), .B2(G20), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n289), .A2(new_n377), .B1(new_n286), .B2(new_n277), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n354), .A2(KEYINPUT74), .A3(new_n356), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n359), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT18), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n348), .B2(new_n353), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n266), .A2(new_n355), .A3(new_n298), .A4(new_n349), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n386), .A2(new_n376), .A3(new_n378), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n386), .A2(new_n376), .A3(KEYINPUT75), .A4(new_n378), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT17), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n359), .A2(new_n379), .A3(new_n392), .A4(new_n380), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n382), .A2(new_n388), .A3(new_n391), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n277), .A2(new_n276), .B1(new_n222), .B2(new_n247), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT70), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT15), .B(G87), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n398), .B(new_n399), .C1(new_n278), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n284), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n290), .A2(G77), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n288), .A2(new_n403), .B1(G77), .B2(new_n285), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G244), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n266), .B1(new_n270), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n244), .A2(G232), .A3(new_n245), .ZN(new_n410));
  INV_X1    g0210(.A(G107), .ZN(new_n411));
  INV_X1    g0211(.A(G238), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n410), .B1(new_n411), .B2(new_n244), .C1(new_n248), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n252), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n406), .B1(G200), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n298), .B2(new_n415), .ZN(new_n417));
  AOI21_X1  g0217(.A(G169), .B1(new_n409), .B2(new_n414), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n404), .B1(new_n401), .B2(new_n284), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT71), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT71), .ZN(new_n421));
  INV_X1    g0221(.A(new_n414), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n293), .B1(new_n422), .B2(new_n408), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n406), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G179), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n409), .A2(new_n425), .A3(new_n414), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n417), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n304), .A2(new_n340), .A3(new_n395), .A4(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n341), .A2(new_n343), .A3(G238), .A4(new_n245), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n341), .A2(new_n343), .A3(G244), .A4(G1698), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G116), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n252), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n264), .A2(G1), .A3(G274), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n268), .A2(G45), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n211), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n267), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n293), .ZN(new_n440));
  NAND3_X1  g0240(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n441), .A2(new_n222), .ZN(new_n442));
  INV_X1    g0242(.A(G97), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n210), .A2(new_n443), .A3(new_n411), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT81), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(G87), .A2(G97), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(KEYINPUT81), .A3(new_n411), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n442), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n341), .A2(new_n343), .A3(new_n222), .A4(G68), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT19), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n278), .B2(new_n443), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n284), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n400), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(new_n285), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n281), .A2(new_n221), .A3(new_n283), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n280), .A2(G1), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n458), .A2(new_n285), .A3(new_n455), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n454), .A2(new_n457), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n434), .A2(new_n438), .A3(new_n425), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n288), .A2(new_n459), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G87), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n454), .A3(new_n457), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n383), .B1(new_n434), .B2(new_n438), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n439), .A2(new_n298), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n440), .A2(new_n464), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT5), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n436), .B1(new_n351), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT79), .B1(new_n476), .B2(G41), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT79), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n474), .A2(KEYINPUT78), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n474), .A2(KEYINPUT78), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n478), .B(new_n259), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n475), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G257), .A3(new_n267), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n341), .A2(new_n343), .A3(G244), .A4(new_n245), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT77), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n244), .A2(G244), .A3(new_n245), .A4(new_n486), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n244), .A2(G250), .A3(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n252), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n258), .A2(new_n481), .A3(new_n477), .A4(new_n475), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n483), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n293), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n497), .A2(new_n443), .A3(G107), .ZN(new_n498));
  XNOR2_X1  g0298(.A(G97), .B(G107), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n500), .A2(new_n222), .B1(new_n247), .B2(new_n276), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n411), .B1(new_n371), .B2(new_n372), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n284), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(G97), .B1(new_n288), .B2(new_n459), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT76), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n285), .A2(new_n443), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n483), .A2(new_n493), .A3(new_n425), .A4(new_n494), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n496), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n495), .A2(new_n383), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n475), .A2(new_n477), .A3(new_n481), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n258), .B1(new_n492), .B2(new_n252), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n298), .A3(new_n483), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT80), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n512), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n499), .A2(new_n497), .ZN(new_n520));
  INV_X1    g0320(.A(new_n498), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(G20), .B1(G77), .B2(new_n275), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n361), .B2(new_n363), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n458), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n509), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n525), .B1(new_n507), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(G200), .B1(new_n515), .B2(new_n483), .ZN(new_n528));
  AND4_X1   g0328(.A1(new_n298), .A2(new_n483), .A3(new_n493), .A4(new_n494), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n496), .A2(new_n510), .A3(new_n511), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT80), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n519), .A2(new_n532), .ZN(new_n533));
  OR3_X1    g0333(.A1(new_n432), .A2(KEYINPUT84), .A3(G20), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT84), .B1(new_n432), .B2(G20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n411), .A2(G20), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT23), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT23), .B1(new_n411), .B2(G20), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n534), .B(new_n535), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n244), .A2(new_n222), .A3(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n244), .A2(new_n222), .A3(G87), .A4(new_n542), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT24), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n284), .B1(new_n546), .B2(KEYINPUT24), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n288), .A2(new_n411), .A3(new_n459), .ZN(new_n550));
  INV_X1    g0350(.A(G13), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(G1), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n222), .A2(G107), .ZN(new_n553));
  OR2_X1    g0353(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n554));
  NAND2_X1  g0354(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n552), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n536), .A2(G1), .A3(new_n551), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n555), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(KEYINPUT86), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT86), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n550), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n548), .A2(new_n549), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n482), .A2(G264), .A3(new_n267), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n244), .A2(G257), .A3(G1698), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G294), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n565), .B(new_n566), .C1(new_n307), .C2(new_n211), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n252), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n494), .A3(new_n568), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n569), .A2(G179), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n293), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n563), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n559), .B(KEYINPUT86), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n544), .A2(new_n545), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n540), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n284), .A3(new_n547), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n564), .A2(new_n568), .A3(G190), .A4(new_n494), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n569), .A2(G200), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n573), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n293), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n482), .A2(G270), .A3(new_n267), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n342), .A2(G33), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n588));
  OAI21_X1  g0388(.A(G303), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n341), .A2(new_n343), .A3(G264), .A4(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n341), .A2(new_n343), .A3(G257), .A4(new_n245), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n252), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n482), .B2(new_n350), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n585), .B1(new_n586), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n482), .A2(G270), .A3(new_n267), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(G179), .A3(new_n494), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n465), .A2(G116), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n286), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(G20), .B1(G33), .B2(G283), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n280), .A2(G97), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n602), .A2(new_n603), .B1(G20), .B2(new_n600), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n284), .A2(KEYINPUT20), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT20), .B1(new_n284), .B2(new_n604), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n599), .B(new_n601), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n596), .A2(new_n494), .A3(new_n593), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(G169), .A3(new_n607), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n598), .A2(new_n607), .B1(new_n609), .B2(new_n584), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(G200), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n514), .A2(new_n258), .B1(new_n252), .B2(new_n592), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(G190), .A3(new_n596), .ZN(new_n613));
  INV_X1    g0413(.A(new_n607), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n583), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n585), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n612), .B2(new_n596), .ZN(new_n618));
  AND4_X1   g0418(.A1(G179), .A2(new_n596), .A3(new_n494), .A4(new_n593), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n607), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n609), .A2(new_n584), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n583), .A2(new_n620), .A3(new_n615), .A4(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n582), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  NOR4_X1   g0423(.A1(new_n429), .A2(new_n473), .A3(new_n533), .A4(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n429), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n293), .B1(new_n612), .B2(new_n596), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT21), .B1(new_n626), .B2(new_n607), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n614), .B1(new_n595), .B2(new_n597), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT89), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT89), .B1(new_n620), .B2(new_n621), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n572), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n580), .A2(new_n530), .A3(new_n531), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n439), .A2(G200), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n445), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT81), .B1(new_n447), .B2(new_n411), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n450), .B(new_n452), .C1(new_n638), .C2(new_n442), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n456), .B1(new_n639), .B2(new_n284), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n635), .A2(new_n640), .A3(new_n466), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(KEYINPUT88), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT88), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n471), .B1(new_n469), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n440), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n439), .A2(KEYINPUT87), .A3(new_n293), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n462), .A2(new_n463), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n642), .A2(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n634), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n632), .A2(new_n633), .A3(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n563), .A2(new_n571), .A3(new_n570), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n629), .B1(new_n627), .B2(new_n628), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n620), .A2(KEYINPUT89), .A3(new_n621), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n649), .B1(new_n646), .B2(new_n647), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n470), .B1(new_n641), .B2(KEYINPUT88), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n469), .A2(new_n643), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(new_n531), .A3(new_n530), .A4(new_n580), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT90), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n512), .A2(new_n472), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n657), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT91), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n496), .A2(new_n510), .A3(new_n666), .A4(new_n511), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n531), .A2(KEYINPUT91), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n660), .A2(new_n665), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n652), .A2(new_n662), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n625), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n376), .A2(new_n378), .B1(new_n354), .B2(new_n356), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n427), .A2(KEYINPUT92), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT92), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n420), .A2(new_n424), .A3(new_n676), .A4(new_n426), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n678), .A2(new_n335), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n389), .B(KEYINPUT17), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n338), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n674), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n302), .A2(new_n303), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n295), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n672), .A2(new_n684), .ZN(G369));
  NAND2_X1  g0485(.A1(new_n552), .A2(new_n222), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n616), .A2(new_n622), .B1(new_n614), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n654), .A2(new_n655), .A3(new_n607), .A4(new_n691), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT93), .ZN(new_n698));
  INV_X1    g0498(.A(new_n580), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n692), .B1(new_n573), .B2(new_n577), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n572), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n653), .A2(new_n692), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n697), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n703), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT93), .B1(new_n696), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n610), .A2(new_n691), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n701), .A2(new_n708), .B1(new_n653), .B2(new_n692), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n218), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n351), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G1), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n638), .A2(new_n600), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n714), .A2(new_n715), .B1(new_n224), .B2(new_n713), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n717));
  XNOR2_X1  g0517(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n671), .A2(new_n692), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n610), .A2(new_n572), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n651), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n657), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n660), .A2(new_n667), .A3(new_n668), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT26), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n723), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .A3(new_n692), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n472), .B(new_n692), .C1(new_n519), .C2(new_n532), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT96), .B1(new_n623), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n620), .A2(new_n615), .A3(new_n621), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT82), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n610), .A2(new_n583), .A3(new_n615), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n581), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT96), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n518), .B1(new_n512), .B2(new_n517), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n530), .A2(KEYINPUT80), .A3(new_n531), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n473), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n737), .A2(new_n738), .A3(new_n741), .A4(new_n692), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n733), .A2(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n252), .A2(new_n433), .B1(new_n267), .B2(new_n437), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G179), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n495), .A2(new_n608), .A3(new_n569), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n564), .A2(new_n744), .A3(new_n568), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n495), .A2(new_n597), .A3(new_n747), .A4(KEYINPUT30), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n495), .A2(new_n747), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(new_n750), .B2(new_n619), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n746), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT95), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n692), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n746), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n483), .A2(new_n493), .A3(new_n494), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n564), .A2(new_n744), .A3(new_n568), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT30), .B1(new_n758), .B2(new_n597), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n750), .A2(new_n749), .A3(new_n619), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT31), .B1(new_n754), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT31), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n692), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n752), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n731), .B1(new_n743), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n730), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n718), .B1(new_n769), .B2(G1), .ZN(G364));
  NAND2_X1  g0570(.A1(new_n222), .A2(G13), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n268), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n712), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n697), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G330), .B2(new_n695), .ZN(new_n777));
  INV_X1    g0577(.A(new_n775), .ZN(new_n778));
  OAI21_X1  g0578(.A(G20), .B1(KEYINPUT99), .B2(G169), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(KEYINPUT99), .A2(G169), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n221), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n425), .A2(new_n383), .A3(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n443), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n222), .A2(new_n425), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n298), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n222), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(new_n298), .A3(G200), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n791), .A2(new_n208), .B1(new_n793), .B2(new_n411), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n789), .A2(G190), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n787), .B(new_n794), .C1(G68), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G159), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT32), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n800), .A2(KEYINPUT32), .B1(new_n803), .B2(G87), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n788), .A2(new_n797), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n244), .B1(new_n805), .B2(new_n247), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n788), .A2(G190), .A3(new_n383), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(G58), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n796), .A2(new_n801), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n362), .B1(new_n805), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(G329), .C2(new_n799), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n790), .A2(G326), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n795), .A2(new_n817), .B1(new_n803), .B2(G303), .ZN(new_n818));
  INV_X1    g0618(.A(new_n793), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G283), .B1(new_n785), .B2(G294), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n815), .A2(new_n816), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n783), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n782), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n711), .A2(new_n600), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT98), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n362), .B1(new_n828), .B2(G355), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(G355), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n711), .A2(new_n244), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(G45), .B2(new_n224), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n242), .A2(G45), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n827), .B1(new_n711), .B2(new_n830), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n778), .B(new_n822), .C1(new_n826), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n825), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n695), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n777), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  NOR2_X1   g0639(.A1(new_n419), .A2(new_n692), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n675), .A2(new_n677), .A3(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n417), .B(new_n427), .C1(new_n419), .C2(new_n692), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n428), .A2(new_n692), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n719), .A2(new_n844), .B1(new_n671), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(new_n768), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n768), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(new_n778), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n782), .A2(new_n823), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n775), .B1(G77), .B2(new_n851), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n793), .A2(new_n210), .B1(new_n798), .B2(new_n813), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT100), .Z(new_n854));
  OAI21_X1  g0654(.A(new_n362), .B1(new_n805), .B2(new_n600), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G294), .B2(new_n808), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n787), .B1(G283), .B2(new_n795), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n790), .A2(G303), .B1(new_n803), .B2(G107), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n854), .A2(new_n856), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n793), .A2(new_n321), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n244), .B1(new_n798), .B2(new_n861), .C1(new_n208), .C2(new_n802), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(G58), .C2(new_n785), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT101), .ZN(new_n864));
  INV_X1    g0664(.A(new_n805), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n808), .A2(G143), .B1(new_n865), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  INV_X1    g0667(.A(new_n795), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n866), .B1(new_n791), .B2(new_n867), .C1(new_n274), .C2(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT34), .Z(new_n870));
  OAI21_X1  g0670(.A(new_n859), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n852), .B1(new_n871), .B2(new_n782), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n843), .B2(new_n824), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n849), .A2(new_n873), .ZN(G384));
  OR2_X1    g0674(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n223), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  OR3_X1    g0678(.A1(new_n224), .A2(new_n247), .A3(new_n367), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n208), .A2(G68), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n268), .B(G13), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n671), .A2(new_n845), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n427), .A2(new_n691), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n386), .A2(new_n376), .A3(new_n378), .ZN(new_n890));
  INV_X1    g0690(.A(new_n689), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n379), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n381), .A2(new_n889), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n358), .A2(new_n357), .B1(new_n376), .B2(new_n378), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n392), .B1(new_n894), .B2(new_n380), .ZN(new_n895));
  INV_X1    g0695(.A(new_n393), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n892), .B1(new_n897), .B2(new_n680), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n379), .A2(new_n357), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n892), .A3(new_n890), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n888), .B(new_n893), .C1(new_n898), .C2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n892), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n394), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n893), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT38), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n337), .A2(new_n692), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n335), .A2(new_n338), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n335), .B2(new_n338), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n887), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n674), .A2(new_n891), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n883), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n902), .A2(new_n906), .A3(KEYINPUT39), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT103), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n387), .B2(new_n673), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n899), .A2(KEYINPUT103), .A3(new_n890), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(new_n892), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n905), .B1(KEYINPUT37), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n892), .B1(new_n680), .B2(new_n674), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n888), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT39), .B1(new_n924), .B2(new_n906), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n917), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n335), .A2(new_n691), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n885), .B1(new_n671), .B2(new_n845), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n912), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n907), .ZN(new_n932));
  INV_X1    g0732(.A(new_n915), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(KEYINPUT102), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n916), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n721), .A2(new_n729), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n684), .B1(new_n936), .B2(new_n429), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n691), .B1(new_n761), .B2(KEYINPUT95), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n753), .B(new_n755), .C1(new_n759), .C2(new_n760), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n939), .A2(new_n764), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n763), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n743), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n924), .A2(new_n906), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n843), .B1(new_n910), .B2(new_n911), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT40), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n945), .B1(new_n743), .B2(new_n942), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT40), .B1(new_n902), .B2(new_n906), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n429), .B1(new_n743), .B2(new_n942), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n731), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n938), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n268), .B2(new_n772), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n938), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n882), .B1(new_n957), .B2(new_n958), .ZN(G367));
  OR2_X1    g0759(.A1(new_n730), .A2(new_n768), .ZN(new_n960));
  INV_X1    g0760(.A(new_n709), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n530), .B(new_n531), .C1(new_n527), .C2(new_n692), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n512), .A2(new_n691), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n961), .A2(KEYINPUT109), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT109), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n709), .B2(new_n964), .ZN(new_n968));
  XNOR2_X1  g0768(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n966), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(new_n966), .B2(new_n968), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n961), .A2(KEYINPUT44), .A3(new_n965), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n709), .B2(new_n964), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(KEYINPUT110), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT110), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n978), .B(new_n975), .C1(new_n709), .C2(new_n964), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n707), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n703), .B(new_n708), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(new_n696), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n960), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n712), .B(KEYINPUT41), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n773), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n964), .B(KEYINPUT105), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n990), .A2(new_n653), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n692), .B1(new_n991), .B2(new_n512), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT42), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n703), .A2(new_n708), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n965), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n703), .A2(KEYINPUT42), .A3(new_n708), .A4(new_n964), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n467), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n660), .B1(new_n999), .B2(new_n692), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n657), .A2(new_n467), .A3(new_n691), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(KEYINPUT43), .B2(new_n1002), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n998), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT107), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n992), .A2(new_n997), .A3(new_n1005), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT106), .Z(new_n1010));
  INV_X1    g0810(.A(new_n707), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n990), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1008), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n989), .A2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n234), .A2(new_n711), .A3(new_n244), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n826), .B1(new_n218), .B2(new_n400), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n775), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(G159), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n868), .A2(new_n1022), .B1(new_n802), .B2(new_n366), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G68), .B2(new_n785), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n807), .A2(new_n274), .B1(new_n805), .B2(new_n208), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n362), .B(new_n1025), .C1(G137), .C2(new_n799), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n790), .A2(G143), .B1(new_n819), .B2(G77), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n244), .B1(new_n799), .B2(G317), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n443), .B2(new_n793), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT112), .Z(new_n1031));
  AOI22_X1  g0831(.A1(new_n865), .A2(G283), .B1(G107), .B2(new_n785), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT111), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n803), .A2(G116), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT46), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G311), .A2(new_n790), .B1(new_n808), .B2(G303), .ZN(new_n1037));
  INV_X1    g0837(.A(G294), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1036), .B(new_n1037), .C1(new_n1038), .C2(new_n868), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1028), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT47), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1021), .B1(new_n1041), .B2(new_n782), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1000), .A2(new_n825), .A3(new_n1001), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1018), .A2(new_n1044), .ZN(G387));
  AOI22_X1  g0845(.A1(new_n808), .A2(G317), .B1(new_n865), .B2(G303), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n791), .B2(new_n811), .C1(new_n813), .C2(new_n868), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n803), .A2(G294), .B1(new_n785), .B2(G283), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT49), .Z(new_n1053));
  AOI21_X1  g0853(.A(new_n244), .B1(new_n799), .B2(G326), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n600), .B2(new_n793), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n786), .A2(new_n400), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G50), .B2(new_n808), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT114), .Z(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT113), .B(G150), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n244), .B1(new_n798), .B2(new_n1060), .C1(new_n321), .C2(new_n805), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n868), .A2(new_n277), .B1(new_n443), .B2(new_n793), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n791), .A2(new_n1022), .B1(new_n802), .B2(new_n247), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n782), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n231), .A2(new_n264), .A3(new_n244), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n277), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT50), .B1(new_n277), .B2(G50), .ZN(new_n1068));
  AOI21_X1  g0868(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n715), .B1(new_n1070), .B2(new_n362), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n218), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n826), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G107), .B2(new_n711), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n778), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1065), .B(new_n1075), .C1(new_n703), .C2(new_n836), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n712), .B1(new_n960), .B2(new_n985), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n769), .A2(new_n986), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1076), .B1(new_n773), .B2(new_n985), .C1(new_n1077), .C2(new_n1078), .ZN(G393));
  NOR2_X1   g0879(.A1(new_n960), .A2(new_n985), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n713), .B1(new_n983), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1080), .B2(new_n983), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n983), .A2(new_n774), .ZN(new_n1083));
  INV_X1    g0883(.A(G283), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n802), .A2(new_n1084), .B1(new_n798), .B2(new_n811), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT115), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n362), .B1(new_n805), .B2(new_n1038), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G107), .B2(new_n819), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n795), .A2(G303), .B1(G116), .B2(new_n785), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G317), .A2(new_n790), .B1(new_n808), .B2(G311), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G150), .A2(new_n790), .B1(new_n808), .B2(G159), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT51), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n786), .A2(new_n247), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G50), .B2(new_n795), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n805), .A2(new_n277), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n362), .B1(new_n799), .B2(G143), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n803), .A2(G68), .B1(new_n819), .B2(G87), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1092), .A2(new_n1094), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n782), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n239), .A2(new_n831), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1073), .B1(G97), .B2(new_n711), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n778), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(new_n990), .C2(new_n836), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1082), .A2(new_n1083), .A3(new_n1108), .ZN(G390));
  NAND2_X1  g0909(.A1(new_n743), .A2(new_n767), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(G330), .A3(new_n843), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n731), .B1(new_n743), .B2(new_n942), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1111), .A2(new_n912), .B1(new_n946), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1110), .A2(G330), .A3(new_n843), .A4(new_n913), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n728), .A2(new_n692), .A3(new_n843), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1115), .A2(new_n886), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n913), .B1(new_n1112), .B2(new_n843), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1113), .A2(new_n930), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n943), .A2(G330), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n429), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n937), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n928), .B1(new_n924), .B2(new_n906), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1116), .B2(new_n912), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n928), .B1(new_n887), .B2(new_n913), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n926), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1120), .A2(new_n945), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1125), .B(new_n1114), .C1(new_n1126), .C2(new_n926), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1119), .A2(new_n1129), .A3(new_n1130), .A4(new_n1122), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n712), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1129), .A2(new_n774), .A3(new_n1130), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT116), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n807), .A2(new_n861), .B1(new_n805), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n362), .B(new_n1138), .C1(G125), .C2(new_n799), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n802), .A2(new_n1060), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n795), .A2(G137), .B1(new_n819), .B2(G50), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n786), .A2(new_n1022), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G128), .B2(new_n790), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n805), .A2(new_n443), .B1(new_n798), .B2(new_n1038), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n244), .B(new_n1146), .C1(G116), .C2(new_n808), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n795), .A2(G107), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1097), .B1(G283), .B2(new_n790), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n860), .B1(G87), .B2(new_n803), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n783), .B1(new_n1145), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n778), .B(new_n1152), .C1(new_n277), .C2(new_n850), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n926), .B2(new_n824), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1135), .A2(new_n1136), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1136), .B1(new_n1135), .B2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1134), .B1(new_n1155), .B2(new_n1156), .ZN(G378));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n292), .A2(new_n891), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n304), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n304), .A2(new_n1160), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1159), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1161), .A3(new_n1158), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n952), .B2(G330), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n947), .A2(KEYINPUT40), .B1(new_n949), .B2(new_n950), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1169), .A2(new_n731), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n935), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1169), .B2(new_n731), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n915), .B1(new_n931), .B2(new_n907), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1174), .A2(KEYINPUT102), .B1(new_n928), .B2(new_n926), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n951), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT40), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n949), .B2(new_n944), .ZN(new_n1178));
  OAI211_X1 g0978(.A(G330), .B(new_n1167), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1173), .A2(new_n1175), .A3(new_n1179), .A4(new_n916), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n774), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1170), .A2(new_n823), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n775), .B1(G50), .B2(new_n851), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n263), .B2(new_n362), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n807), .A2(new_n411), .B1(new_n805), .B2(new_n400), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n263), .B(new_n362), .C1(new_n1084), .C2(new_n798), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n793), .A2(new_n366), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G116), .B2(new_n790), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n795), .A2(G97), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n803), .A2(G77), .B1(new_n785), .B2(G68), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1189), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1186), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n808), .A2(G128), .B1(new_n865), .B2(G137), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n802), .B2(new_n1137), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n790), .A2(G125), .B1(G150), .B2(new_n785), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT117), .Z(new_n1201));
  AOI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(G132), .C2(new_n795), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT59), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1197), .B1(new_n1022), .B2(new_n793), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1196), .B1(new_n1195), .B2(new_n1194), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1184), .B1(new_n1206), .B2(new_n782), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1183), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1182), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1117), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1118), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n731), .B(new_n844), .C1(new_n743), .C2(new_n767), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1212), .A2(new_n913), .B1(new_n1120), .B2(new_n945), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1210), .A2(new_n1211), .B1(new_n1213), .B2(new_n887), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1122), .B1(new_n1131), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1180), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1173), .A2(new_n1179), .B1(new_n1175), .B2(new_n916), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n713), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT118), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1172), .A2(new_n1221), .A3(new_n1180), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1219), .B1(new_n1133), .B2(new_n1122), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1217), .A2(KEYINPUT118), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1209), .B1(new_n1220), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(G375));
  OR2_X1    g1027(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n988), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1123), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n912), .A2(new_n823), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT119), .Z(new_n1232));
  AOI21_X1  g1032(.A(new_n778), .B1(new_n321), .B2(new_n850), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n244), .B1(new_n799), .B2(G303), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n411), .B2(new_n805), .C1(new_n1084), .C2(new_n807), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1057), .B(new_n1235), .C1(G77), .C2(new_n819), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n600), .A2(new_n868), .B1(new_n791), .B2(new_n1038), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G97), .B2(new_n803), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n786), .A2(new_n208), .B1(new_n802), .B2(new_n1022), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G132), .B2(new_n790), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n362), .B1(new_n799), .B2(G128), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n867), .B2(new_n807), .C1(new_n274), .C2(new_n805), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n868), .A2(new_n1137), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1242), .A2(new_n1190), .A3(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1236), .A2(new_n1238), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1232), .B(new_n1233), .C1(new_n783), .C2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1214), .B2(new_n773), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1230), .A2(new_n1248), .ZN(G381));
  INV_X1    g1049(.A(G390), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n989), .A2(new_n1017), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1253), .A2(G375), .A3(G378), .A4(G381), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT120), .Z(G407));
  INV_X1    g1055(.A(G378), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1226), .A2(new_n1256), .A3(new_n690), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(G407), .A2(G213), .A3(new_n1257), .ZN(G409));
  XNOR2_X1  g1058(.A(G393), .B(new_n838), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(G387), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1259), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(new_n1251), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1250), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1251), .B2(KEYINPUT124), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1265), .B(G390), .C1(new_n1251), .C2(new_n1262), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1123), .A2(KEYINPUT60), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1228), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT122), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1268), .A2(KEYINPUT122), .A3(new_n1228), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n713), .B1(new_n1273), .B2(KEYINPUT60), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1271), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G384), .A2(KEYINPUT123), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1248), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(G213), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(G343), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1275), .A2(new_n1248), .ZN(new_n1283));
  XOR2_X1   g1083(.A(G384), .B(KEYINPUT123), .Z(new_n1284));
  OAI211_X1 g1084(.A(new_n1278), .B(new_n1282), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1275), .A2(new_n1248), .A3(new_n1277), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1284), .B1(new_n1275), .B2(new_n1248), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1281), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1181), .A2(new_n774), .B1(new_n1183), .B2(new_n1207), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1172), .A2(new_n1180), .B1(new_n1133), .B2(new_n1122), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n712), .B1(new_n1291), .B2(KEYINPUT57), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G378), .B(new_n1290), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT121), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1220), .A2(new_n1225), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1297), .A2(KEYINPUT121), .A3(G378), .A4(new_n1290), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1222), .A2(new_n774), .A3(new_n1224), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1299), .B(new_n1208), .C1(new_n988), .C2(new_n1218), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1296), .A2(new_n1298), .B1(new_n1256), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1289), .B1(new_n1301), .B2(new_n1280), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1256), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1280), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1278), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1267), .B(new_n1302), .C1(new_n1308), .C2(KEYINPUT62), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1264), .B(new_n1266), .C1(new_n1309), .C2(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1278), .B(KEYINPUT63), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT125), .B1(new_n1305), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT125), .ZN(new_n1315));
  NOR4_X1   g1115(.A1(new_n1301), .A2(new_n1315), .A3(new_n1280), .A4(new_n1312), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1301), .A2(new_n1280), .A3(new_n1306), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1302), .B(new_n1318), .C1(new_n1319), .C2(KEYINPUT63), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1317), .A2(new_n1320), .A3(KEYINPUT126), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1302), .A2(new_n1318), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT63), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1298), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT121), .B1(new_n1226), .B2(G378), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1304), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1280), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n1329), .A3(new_n1313), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1315), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1305), .A2(KEYINPUT125), .A3(new_n1313), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1322), .B1(new_n1325), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1311), .B1(new_n1321), .B2(new_n1334), .ZN(G405));
  NAND2_X1  g1135(.A1(G375), .A2(new_n1256), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1303), .A2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1307), .B1(new_n1337), .B2(KEYINPUT127), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1338), .B1(KEYINPUT127), .B2(new_n1337), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1337), .A2(KEYINPUT127), .A3(new_n1306), .ZN(new_n1341));
  OR3_X1    g1141(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1340), .B1(new_n1339), .B2(new_n1341), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(G402));
endmodule


