//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT70), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT71), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(new_n457), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT72), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT72), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT73), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n471), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT73), .A4(KEYINPUT3), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT72), .B(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT3), .B(G2104), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G125), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT75), .Z(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(new_n474), .B2(new_n475), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT74), .Z(new_n496));
  AOI211_X1 g071(.A(new_n493), .B(new_n496), .C1(G136), .C2(new_n476), .ZN(G162));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR4_X1   g073(.A1(new_n484), .A2(KEYINPUT4), .A3(new_n498), .A4(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n472), .B1(new_n478), .B2(KEYINPUT3), .ZN(new_n500));
  AND4_X1   g075(.A1(KEYINPUT73), .A2(new_n467), .A3(new_n469), .A4(KEYINPUT3), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n491), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n499), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(G126), .B(G2105), .C1(new_n500), .C2(new_n501), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n503), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  XOR2_X1   g087(.A(new_n512), .B(KEYINPUT76), .Z(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(new_n514), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G166));
  AOI22_X1  g098(.A1(new_n517), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n514), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n520), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n526), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n526), .B2(new_n530), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n518), .A2(new_n535), .B1(new_n520), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n511), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(new_n514), .A2(G56), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n511), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n517), .A2(new_n514), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n517), .A2(G543), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT79), .B(G43), .Z(new_n548));
  AOI22_X1  g123(.A1(G81), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n543), .A2(new_n544), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT80), .Z(G188));
  NAND2_X1  g134(.A1(new_n547), .A2(G53), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT9), .Z(new_n561));
  AOI22_X1  g136(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n511), .B1(new_n518), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  OAI21_X1  g144(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT81), .Z(new_n571));
  AOI22_X1  g146(.A1(G87), .A2(new_n546), .B1(new_n547), .B2(G49), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n546), .A2(G86), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n547), .A2(G48), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n511), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n518), .A2(new_n581), .B1(new_n520), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n511), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n546), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n525), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n547), .B2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT82), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n589), .B1(new_n598), .B2(new_n588), .ZN(G284));
  AOI21_X1  g174(.A(new_n589), .B1(new_n598), .B2(new_n588), .ZN(G321));
  NOR2_X1   g175(.A1(G286), .A2(new_n588), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n588), .B2(new_n565), .ZN(G297));
  AOI21_X1  g177(.A(new_n601), .B1(new_n588), .B2(new_n565), .ZN(G280));
  XNOR2_X1  g178(.A(KEYINPUT83), .B(G559), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(G860), .B2(new_n605), .ZN(G148));
  NAND2_X1  g181(.A1(new_n552), .A2(new_n588), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n597), .A2(new_n604), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n588), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n479), .A2(new_n483), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n476), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n494), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n491), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(G2096), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT85), .ZN(G156));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT86), .Z(new_n638));
  OAI21_X1  g213(.A(G14), .B1(new_n635), .B2(new_n636), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT17), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT88), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  INV_X1    g224(.A(new_n642), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n649), .B(new_n646), .C1(new_n650), .C2(new_n644), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n644), .A3(new_n645), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n648), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n662), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n664), .B(new_n666), .C1(new_n659), .C2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n675), .A2(G23), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(G288), .B2(G16), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT33), .ZN(new_n678));
  INV_X1    g253(.A(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(G22), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n675), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT92), .Z(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(G1971), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(G1971), .ZN(new_n685));
  NOR2_X1   g260(.A1(G6), .A2(G16), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n579), .B2(G16), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n680), .A2(new_n684), .A3(new_n685), .A4(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT34), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT90), .B(G29), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G25), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n476), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n494), .A2(G119), .ZN(new_n696));
  OR2_X1    g271(.A1(G95), .A2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G107), .C2(new_n491), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT91), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n586), .A2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G16), .B2(G24), .ZN(new_n708));
  INV_X1    g283(.A(G1986), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n709), .B2(new_n708), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n691), .A2(new_n704), .A3(new_n705), .A4(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n675), .A2(G4), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n598), .B2(new_n675), .ZN(new_n717));
  INV_X1    g292(.A(G1348), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n692), .A2(G35), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT101), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n692), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT29), .B(G2090), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n494), .A2(G129), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT26), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n479), .A2(G105), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n476), .A2(G141), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(G32), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G1996), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT24), .B(G34), .ZN(new_n739));
  AOI22_X1  g314(.A1(G160), .A2(G29), .B1(new_n692), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n737), .A2(new_n738), .B1(G2084), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G5), .A2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT98), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G301), .B2(new_n675), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT99), .ZN(new_n747));
  NOR2_X1   g322(.A1(G16), .A2(G19), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n553), .B2(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G1341), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G11), .Z(new_n751));
  NOR2_X1   g326(.A1(new_n620), .A2(new_n692), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n735), .B1(new_n753), .B2(G28), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT97), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n755), .A2(KEYINPUT97), .B1(new_n753), .B2(G28), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n751), .B(new_n752), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n476), .A2(G139), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n491), .A2(G103), .A3(G2104), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n483), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n759), .B(new_n762), .C1(new_n491), .C2(new_n763), .ZN(new_n764));
  MUX2_X1   g339(.A(G33), .B(new_n764), .S(G29), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G2072), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n747), .A2(new_n750), .A3(new_n758), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n675), .A2(G20), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT23), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n565), .B2(new_n675), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  OAI22_X1  g346(.A1(new_n749), .A2(G1341), .B1(G2072), .B2(new_n765), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n767), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n719), .A2(new_n724), .A3(new_n741), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT96), .B1(G16), .B2(G21), .ZN(new_n775));
  NAND2_X1  g350(.A1(G168), .A2(G16), .ZN(new_n776));
  MUX2_X1   g351(.A(KEYINPUT96), .B(new_n775), .S(new_n776), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1966), .ZN(new_n778));
  NOR2_X1   g353(.A1(G164), .A2(new_n692), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G27), .B2(new_n692), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n692), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n476), .A2(G140), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n494), .A2(G128), .ZN(new_n788));
  OR2_X1    g363(.A1(G104), .A2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n789), .B(G2104), .C1(G116), .C2(new_n491), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n787), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n786), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2067), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n778), .A2(new_n782), .A3(new_n783), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n744), .A2(new_n745), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n796), .B1(G2084), .B2(new_n740), .C1(new_n737), .C2(new_n738), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT100), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n774), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n714), .A2(new_n715), .A3(new_n799), .ZN(G150));
  INV_X1    g375(.A(G150), .ZN(G311));
  NAND2_X1  g376(.A1(new_n598), .A2(G559), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT38), .Z(new_n803));
  INV_X1    g378(.A(G93), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT102), .B(G55), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n518), .A2(new_n804), .B1(new_n520), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT103), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(new_n511), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n552), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n552), .A2(new_n810), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n803), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT39), .ZN(new_n816));
  AOI21_X1  g391(.A(G860), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n810), .A2(G860), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(G145));
  INV_X1    g396(.A(KEYINPUT40), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n823));
  INV_X1    g398(.A(new_n499), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT104), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n504), .A2(new_n826), .A3(new_n508), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n504), .B2(new_n508), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n792), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n476), .A2(G142), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n494), .A2(G130), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n491), .A2(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n830), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n733), .B(new_n764), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n699), .B(new_n613), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n488), .B(new_n620), .Z(new_n841));
  XNOR2_X1  g416(.A(G162), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n836), .A2(new_n839), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT105), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT106), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n842), .B1(new_n840), .B2(new_n843), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(G37), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n847), .B1(new_n846), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n822), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n846), .A2(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT106), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(KEYINPUT40), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n852), .A2(new_n856), .ZN(G395));
  NAND2_X1  g432(.A1(new_n810), .A2(new_n588), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n608), .B(new_n814), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n565), .A2(new_n596), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n565), .A2(new_n596), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n862), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n860), .A2(new_n866), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n871), .A2(new_n872), .B1(new_n860), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n865), .B1(new_n859), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(G305), .B(G288), .ZN(new_n876));
  XOR2_X1   g451(.A(G166), .B(new_n586), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT42), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n875), .B(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n858), .B1(new_n880), .B2(new_n588), .ZN(G295));
  OAI21_X1  g456(.A(new_n858), .B1(new_n880), .B2(new_n588), .ZN(G331));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n883));
  AOI21_X1  g458(.A(G171), .B1(G286), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(G286), .A2(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n814), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n812), .B2(new_n813), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n884), .A3(new_n888), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n874), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n893), .A2(new_n889), .A3(new_n863), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n878), .ZN(new_n896));
  AOI21_X1  g471(.A(G37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n890), .A2(new_n891), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT110), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n868), .A2(new_n870), .A3(new_n873), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(KEYINPUT41), .B2(new_n863), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n898), .A2(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n890), .A2(new_n891), .A3(new_n864), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT110), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n878), .B(new_n902), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n897), .A2(new_n906), .A3(KEYINPUT43), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n892), .B2(new_n894), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n893), .A2(new_n889), .ZN(new_n910));
  OAI211_X1 g485(.A(KEYINPUT109), .B(new_n904), .C1(new_n910), .C2(new_n874), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n878), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT43), .B1(new_n912), .B2(new_n897), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n897), .A2(new_n906), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n912), .B2(new_n897), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n914), .B1(new_n918), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g494(.A(G1384), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT45), .B1(new_n829), .B2(new_n920), .ZN(new_n921));
  AND4_X1   g496(.A1(G40), .A2(new_n477), .A3(new_n487), .A4(new_n480), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(G1996), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT46), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n792), .B(G2067), .Z(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n734), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT47), .Z(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT127), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n733), .B(G1996), .Z(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n926), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n699), .B(new_n703), .Z(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(new_n923), .ZN(new_n935));
  INV_X1    g510(.A(new_n923), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n709), .A3(new_n586), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n935), .B1(KEYINPUT48), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(KEYINPUT48), .B2(new_n938), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n703), .ZN(new_n941));
  OAI22_X1  g516(.A1(new_n932), .A2(new_n941), .B1(G2067), .B2(new_n792), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n936), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n930), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n929), .A2(KEYINPUT127), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(G288), .A2(new_n679), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT115), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n829), .A2(new_n920), .A3(new_n922), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT114), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n950), .A2(new_n951), .A3(G8), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n950), .B2(G8), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT52), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT52), .B1(G288), .B2(new_n679), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n949), .B(new_n956), .C1(new_n952), .C2(new_n953), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT118), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n950), .A2(G8), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT114), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n950), .A2(new_n951), .A3(G8), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(G1981), .B1(new_n576), .B2(new_n578), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n577), .A2(new_n511), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT116), .B(G1981), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n964), .A2(new_n574), .A3(new_n575), .A4(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(KEYINPUT117), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(KEYINPUT117), .B2(new_n963), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n968), .B(KEYINPUT49), .C1(KEYINPUT117), .C2(new_n963), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n958), .B1(new_n962), .B2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n973), .B(new_n958), .C1(new_n952), .C2(new_n953), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n955), .B(new_n957), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  NOR2_X1   g553(.A1(G166), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(G166), .B2(new_n978), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n829), .B2(new_n920), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n920), .B1(new_n503), .B2(new_n509), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n922), .B1(new_n988), .B2(KEYINPUT50), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n987), .A2(new_n989), .A3(G2090), .ZN(new_n990));
  INV_X1    g565(.A(G1971), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT111), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n829), .A2(KEYINPUT45), .A3(new_n920), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n988), .A2(new_n996), .A3(new_n992), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(new_n922), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n990), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n985), .B1(new_n999), .B2(new_n978), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT120), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(new_n985), .C1(new_n999), .C2(new_n978), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n977), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT45), .B(new_n920), .C1(new_n503), .C2(new_n509), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n922), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G126), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n1008), .B(new_n491), .C1(new_n474), .C2(new_n475), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT104), .B1(new_n1009), .B2(new_n507), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n504), .A2(new_n826), .A3(new_n508), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n503), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n992), .B1(new_n1012), .B2(G1384), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1966), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G2084), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n922), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n986), .B1(new_n1012), .B2(G1384), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT50), .B(new_n920), .C1(new_n503), .C2(new_n509), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(G8), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G168), .A2(new_n978), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(KEYINPUT51), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  INV_X1    g599(.A(G1966), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n921), .B2(new_n1006), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1016), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT50), .B1(new_n829), .B2(new_n920), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1018), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1024), .B(G8), .C1(new_n1031), .C2(G286), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1022), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(KEYINPUT125), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT125), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1035), .B(new_n1022), .C1(new_n1026), .C2(new_n1030), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1023), .B(new_n1032), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n998), .B2(G2078), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(G2078), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1007), .A2(new_n1013), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n922), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n745), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(G171), .B(KEYINPUT54), .Z(new_n1045));
  AND2_X1   g620(.A1(new_n997), .A2(new_n922), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(new_n781), .A3(new_n995), .A4(new_n994), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1047), .A2(new_n1038), .B1(new_n745), .B2(new_n1042), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n491), .B1(new_n486), .B2(KEYINPUT126), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(KEYINPUT126), .B2(new_n486), .ZN(new_n1050));
  AND4_X1   g625(.A1(G40), .A2(new_n481), .A3(new_n1040), .A4(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n995), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1045), .B1(new_n1052), .B2(new_n1013), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1044), .A2(new_n1045), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1037), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n998), .A2(new_n991), .ZN(new_n1056));
  INV_X1    g631(.A(G2090), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(new_n922), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(G8), .A3(new_n984), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT113), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n978), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n984), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1004), .A2(new_n1055), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1046), .A2(new_n995), .A3(new_n994), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n564), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n565), .B(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1956), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n987), .B2(new_n989), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n950), .A2(G2067), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1042), .B2(new_n718), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n596), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1075), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT61), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1075), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(new_n1076), .ZN(new_n1087));
  INV_X1    g662(.A(new_n596), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1088), .B(new_n1081), .C1(new_n1042), .C2(new_n718), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT60), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1082), .A2(new_n1091), .A3(new_n1088), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1087), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1085), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1075), .A2(KEYINPUT124), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1078), .A3(new_n1079), .A4(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT58), .B(G1341), .Z(new_n1098));
  NAND2_X1  g673(.A1(new_n950), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n998), .B2(G1996), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n553), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT59), .B(new_n553), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1093), .A2(new_n1097), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1066), .B1(new_n1084), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1110));
  INV_X1    g685(.A(new_n977), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1020), .A2(G286), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1065), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n977), .A2(KEYINPUT119), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n947), .B(KEYINPUT115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n960), .B2(new_n961), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n957), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n973), .B1(new_n952), .B2(new_n953), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n975), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1115), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1112), .B(KEYINPUT63), .C1(new_n1062), .C2(new_n984), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1113), .A2(new_n1114), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n974), .A2(new_n976), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1131), .A2(KEYINPUT119), .A3(new_n1119), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1121), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1131), .A2(G1976), .A3(G288), .ZN(new_n1135));
  INV_X1    g710(.A(new_n967), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n962), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1037), .A2(KEYINPUT62), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1033), .B(KEYINPUT125), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n1023), .A4(new_n1032), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1048), .B2(new_n1041), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1110), .A2(new_n1065), .A3(new_n1111), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1134), .B(new_n1137), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1109), .A2(new_n1129), .A3(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n586), .B(G1986), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n923), .B1(new_n934), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n946), .B1(new_n1146), .B2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g724(.A1(new_n640), .A2(G229), .A3(new_n464), .A4(G227), .ZN(new_n1151));
  OAI21_X1  g725(.A(new_n1151), .B1(new_n916), .B2(new_n917), .ZN(new_n1152));
  NOR2_X1   g726(.A1(new_n850), .A2(new_n851), .ZN(new_n1153));
  NOR2_X1   g727(.A1(new_n1152), .A2(new_n1153), .ZN(G308));
  OAI221_X1 g728(.A(new_n1151), .B1(new_n850), .B2(new_n851), .C1(new_n917), .C2(new_n916), .ZN(G225));
endmodule


