//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1176, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G107), .ZN(new_n204));
  INV_X1    g0004(.A(G264), .ZN(new_n205));
  INV_X1    g0005(.A(G116), .ZN(new_n206));
  INV_X1    g0006(.A(G270), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT64), .B(G77), .Z(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G244), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n208), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n203), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR2_X1   g0029(.A1(G58), .A2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n226), .A2(new_n229), .A3(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n207), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  OAI21_X1  g0051(.A(G20), .B1(new_n231), .B2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n233), .A2(G33), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n252), .B1(new_n253), .B2(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n234), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n258), .A2(new_n260), .B1(new_n222), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n261), .B2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT67), .A2(G223), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT67), .A2(G223), .ZN(new_n275));
  OAI21_X1  g0075(.A(G1698), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n279), .B(new_n280), .C1(new_n214), .C2(new_n273), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G41), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n261), .B(G274), .C1(new_n286), .C2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(new_n280), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n281), .B(new_n287), .C1(new_n223), .C2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT68), .B(G200), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n267), .A2(new_n268), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n293), .B1(new_n268), .B2(new_n267), .C1(new_n294), .C2(new_n291), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G226), .A2(G1698), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n218), .B2(G1698), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n273), .A2(new_n298), .B1(G33), .B2(G97), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n287), .B1(new_n290), .B2(new_n210), .C1(new_n299), .C2(new_n288), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT13), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT13), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n300), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G190), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n255), .A2(new_n222), .B1(new_n233), .B2(G68), .ZN(new_n306));
  INV_X1    g0106(.A(G77), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n256), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n260), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT11), .ZN(new_n310));
  OR3_X1    g0110(.A1(new_n262), .A2(KEYINPUT12), .A3(G68), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT12), .B1(new_n262), .B2(G68), .ZN(new_n312));
  AOI22_X1  g0112(.A1(G68), .A2(new_n265), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n302), .A2(new_n305), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT14), .B1(new_n304), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT70), .B1(new_n301), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT14), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n301), .A2(new_n320), .A3(G169), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT70), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n304), .A2(new_n322), .A3(G179), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n317), .A2(new_n319), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n314), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n315), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n291), .A2(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n291), .A2(new_n316), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n267), .A3(new_n328), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n296), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT71), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT71), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n271), .A3(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(G223), .A2(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n223), .A2(G1698), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n334), .A2(new_n270), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G87), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n280), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n290), .A2(new_n218), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n342), .A3(new_n287), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G200), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n334), .A2(new_n270), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(new_n233), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n331), .A2(new_n333), .B1(KEYINPUT3), .B2(new_n269), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT7), .B1(new_n348), .B2(G20), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n349), .A3(G68), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n217), .A2(new_n209), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n351), .B2(new_n230), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n254), .A2(G159), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n350), .A2(KEYINPUT16), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n273), .B2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n270), .A2(new_n272), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n346), .A2(KEYINPUT72), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n233), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n209), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n357), .B1(new_n363), .B2(new_n354), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n356), .A2(new_n260), .A3(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n340), .A2(G190), .A3(new_n287), .A4(new_n342), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n257), .A2(new_n262), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n265), .B2(new_n257), .ZN(new_n368));
  AND4_X1   g0168(.A1(new_n344), .A2(new_n365), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT17), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n365), .A2(new_n344), .A3(new_n366), .A4(new_n368), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n365), .A2(new_n368), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n343), .A2(G169), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n340), .A2(new_n342), .A3(G179), .A4(new_n287), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT18), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n374), .A2(KEYINPUT18), .A3(new_n377), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n370), .B(new_n373), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  XOR2_X1   g0181(.A(KEYINPUT8), .B(G58), .Z(new_n382));
  AOI22_X1  g0182(.A1(G20), .A2(new_n214), .B1(new_n382), .B2(new_n254), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n256), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n260), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n265), .A2(G77), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n386), .B(new_n387), .C1(new_n214), .C2(new_n262), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G238), .A2(G1698), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n273), .B(new_n389), .C1(new_n218), .C2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(new_n280), .C1(G107), .C2(new_n273), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n288), .A2(new_n215), .A3(new_n289), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n287), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(G190), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n292), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n316), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n388), .B(new_n398), .C1(G179), .C2(new_n393), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g0200(.A(new_n400), .B(KEYINPUT69), .Z(new_n401));
  AND3_X1   g0201(.A1(new_n330), .A2(new_n381), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G244), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(G1698), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n334), .A2(new_n270), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT74), .B(KEYINPUT4), .Z(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G283), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(KEYINPUT4), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G250), .A2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n273), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n280), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT5), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n283), .A2(new_n285), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G45), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(G1), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(G257), .A3(new_n288), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n261), .A2(G45), .A3(G274), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT75), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT75), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n427), .A3(new_n424), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n415), .A2(new_n426), .A3(new_n318), .A4(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n406), .A2(new_n407), .B1(new_n412), .B2(new_n273), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n288), .B1(new_n430), .B2(new_n409), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n316), .B1(new_n431), .B2(new_n425), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n204), .B1(new_n359), .B2(new_n362), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT6), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n434), .A2(new_n219), .A3(G107), .ZN(new_n435));
  XNOR2_X1  g0235(.A(G97), .B(G107), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n437), .A2(new_n233), .B1(new_n307), .B2(new_n255), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n260), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n261), .A2(G33), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n262), .A2(new_n440), .A3(new_n234), .A4(new_n259), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G97), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G97), .B2(new_n263), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT73), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n442), .B(KEYINPUT73), .C1(G97), .C2(new_n263), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n429), .A2(new_n432), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n429), .A2(new_n432), .A3(KEYINPUT77), .A4(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n415), .A2(new_n426), .A3(new_n428), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G200), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT76), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n431), .A2(new_n294), .A3(new_n425), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n448), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(KEYINPUT76), .A3(G200), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n334), .A2(new_n233), .A3(G68), .A4(new_n270), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT19), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n256), .B2(new_n219), .ZN(new_n464));
  NOR2_X1   g0264(.A1(G97), .A2(G107), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n211), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n463), .A2(new_n269), .A3(new_n219), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(G20), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n462), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n260), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n384), .A2(new_n263), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n384), .B(KEYINPUT79), .ZN(new_n472));
  INV_X1    g0272(.A(new_n441), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n419), .A2(new_n212), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n288), .B1(new_n476), .B2(new_n423), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n269), .A2(new_n206), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G238), .A2(G1698), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n404), .B2(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n348), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n318), .B(new_n477), .C1(new_n481), .C2(new_n288), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT78), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n334), .A2(new_n480), .A3(new_n270), .ZN(new_n484));
  INV_X1    g0284(.A(new_n478), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n280), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT78), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(new_n318), .A4(new_n477), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n477), .B1(new_n481), .B2(new_n288), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n316), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n475), .A2(new_n483), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n292), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n469), .A2(new_n260), .B1(new_n263), .B2(new_n384), .ZN(new_n494));
  OAI211_X1 g0294(.A(G190), .B(new_n477), .C1(new_n481), .C2(new_n288), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n473), .A2(G87), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n453), .A2(new_n461), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT80), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n212), .A2(new_n277), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n348), .B(new_n501), .C1(G257), .C2(new_n277), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G294), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n288), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n421), .A2(new_n288), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n205), .ZN(new_n506));
  INV_X1    g0306(.A(new_n424), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n316), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n318), .ZN(new_n511));
  INV_X1    g0311(.A(new_n260), .ZN(new_n512));
  NOR4_X1   g0312(.A1(new_n360), .A2(KEYINPUT22), .A3(G20), .A4(new_n211), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n334), .A2(new_n233), .A3(G87), .A4(new_n270), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT81), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT22), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n513), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT23), .B1(new_n204), .B2(G20), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n204), .A2(KEYINPUT23), .A3(G20), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n521), .A2(new_n522), .B1(new_n478), .B2(new_n233), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT24), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n513), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT22), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n517), .B1(new_n514), .B2(KEYINPUT22), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n530), .A3(new_n523), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n512), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT25), .B1(new_n263), .B2(new_n204), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n204), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n535), .B1(new_n473), .B2(G107), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n510), .B(new_n511), .C1(new_n532), .C2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n529), .A2(new_n530), .A3(new_n523), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n530), .B1(new_n529), .B2(new_n523), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n260), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n508), .A2(G190), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n509), .A2(G200), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n541), .A2(new_n536), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT80), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n453), .A2(new_n461), .A3(new_n546), .A4(new_n498), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n421), .A2(G270), .A3(new_n288), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n220), .A2(new_n277), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n348), .B(new_n549), .C1(G264), .C2(new_n277), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n360), .A2(G303), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n424), .B(new_n548), .C1(new_n552), .C2(new_n288), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n473), .A2(G116), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n409), .B(new_n233), .C1(G33), .C2(new_n219), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n555), .B(new_n260), .C1(new_n233), .C2(G116), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT20), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n554), .B1(G116), .B2(new_n262), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n553), .A2(G169), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n553), .A2(new_n318), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n560), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n553), .A2(KEYINPUT21), .A3(G169), .A4(new_n560), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n553), .A2(G200), .ZN(new_n568));
  INV_X1    g0368(.A(new_n560), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n294), .C2(new_n553), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n500), .A2(new_n545), .A3(new_n547), .A4(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n403), .A2(new_n573), .ZN(G372));
  INV_X1    g0374(.A(new_n329), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n374), .A2(new_n377), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT18), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n374), .A2(KEYINPUT18), .A3(new_n377), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n315), .A2(new_n399), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n325), .B2(new_n324), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n371), .B(KEYINPUT17), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n575), .B1(new_n585), .B2(new_n296), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n475), .A2(new_n491), .A3(new_n482), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n497), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n449), .A2(new_n588), .A3(KEYINPUT26), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n451), .A2(new_n498), .A3(new_n452), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(KEYINPUT26), .ZN(new_n591));
  INV_X1    g0391(.A(new_n588), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n511), .B1(G169), .B2(new_n508), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n541), .B2(new_n536), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n594), .B2(new_n567), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n544), .A2(new_n453), .A3(new_n461), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n587), .B(new_n591), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n586), .B1(new_n403), .B2(new_n598), .ZN(G369));
  INV_X1    g0399(.A(G13), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n600), .A2(G20), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n261), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n602), .A2(KEYINPUT27), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(KEYINPUT27), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(G213), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G343), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n569), .A2(new_n608), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n567), .A2(new_n571), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n567), .A2(new_n609), .ZN(new_n611));
  OAI21_X1  g0411(.A(G330), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n607), .B1(new_n532), .B2(new_n537), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n538), .A2(new_n544), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT82), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n538), .A2(new_n544), .A3(new_n613), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n594), .A2(new_n607), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n612), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n567), .A2(new_n608), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n615), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n594), .A2(new_n608), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n620), .A2(new_n624), .ZN(G399));
  INV_X1    g0425(.A(new_n227), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n286), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G1), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n465), .A2(new_n211), .A3(new_n206), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n629), .A2(new_n630), .B1(new_n232), .B2(new_n628), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT28), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT30), .ZN(new_n633));
  AOI211_X1 g0433(.A(new_n425), .B(new_n431), .C1(KEYINPUT83), .C2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n490), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n504), .A2(new_n506), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n564), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n508), .A2(new_n635), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(new_n318), .A3(new_n454), .A4(new_n553), .ZN(new_n642));
  NOR4_X1   g0442(.A1(new_n553), .A2(new_n318), .A3(new_n504), .A4(new_n506), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n643), .A2(new_n635), .A3(new_n638), .A4(new_n634), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n607), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT31), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(KEYINPUT31), .A3(new_n607), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n648), .B(new_n649), .C1(new_n573), .C2(new_n607), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G330), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n597), .A2(new_n608), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT29), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n590), .A2(KEYINPUT26), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n654), .B(new_n587), .C1(new_n595), .C2(new_n596), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n449), .A2(new_n588), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(KEYINPUT26), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n608), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT29), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n651), .A2(new_n653), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT84), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT84), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n651), .A2(new_n653), .A3(new_n659), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n632), .B1(new_n664), .B2(G1), .ZN(G364));
  NAND2_X1  g0465(.A1(new_n612), .A2(KEYINPUT85), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n610), .A2(new_n611), .ZN(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n666), .B(new_n669), .Z(new_n670));
  NAND2_X1  g0470(.A1(new_n601), .A2(G45), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n628), .A2(G1), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n234), .B1(G20), .B2(new_n316), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n233), .A2(G179), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n292), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G190), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G283), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n360), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT88), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT88), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n683), .A2(new_n294), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(KEYINPUT33), .B(G317), .ZN(new_n686));
  NOR2_X1   g0486(.A1(G190), .A2(G200), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n676), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n685), .A2(new_n686), .B1(G329), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n683), .A2(G190), .A3(new_n684), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G326), .ZN(new_n693));
  INV_X1    g0493(.A(G311), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n233), .A2(new_n318), .A3(KEYINPUT87), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT87), .B1(new_n233), .B2(new_n318), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(new_n696), .A3(new_n687), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n690), .B(new_n693), .C1(new_n694), .C2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n294), .A2(G200), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n695), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  AOI211_X1 g0500(.A(new_n681), .B(new_n698), .C1(G322), .C2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G294), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n318), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G20), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G303), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n677), .A2(new_n294), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI221_X1 g0508(.A(new_n701), .B1(new_n702), .B2(new_n705), .C1(new_n706), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(G87), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n679), .B2(new_n204), .ZN(new_n711));
  INV_X1    g0511(.A(new_n700), .ZN(new_n712));
  INV_X1    g0512(.A(new_n214), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n217), .B1(new_n713), .B2(new_n697), .ZN(new_n714));
  AOI211_X1 g0514(.A(new_n711), .B(new_n714), .C1(G50), .C2(new_n692), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n704), .A2(G97), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT89), .B(G159), .Z(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n688), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT32), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n360), .B1(new_n685), .B2(G68), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n715), .A2(new_n716), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n675), .B1(new_n709), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT86), .Z(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n674), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n273), .A2(G355), .A3(new_n227), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n247), .A2(G45), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n348), .A2(new_n626), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G45), .B2(new_n232), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n729), .B1(G116), .B2(new_n227), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n723), .B1(new_n728), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n667), .A2(new_n727), .ZN(new_n735));
  INV_X1    g0535(.A(new_n672), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n673), .A2(new_n737), .ZN(G396));
  NAND2_X1  g0538(.A1(new_n651), .A2(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n388), .A2(new_n607), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n397), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n399), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n399), .A2(new_n607), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n597), .A2(new_n608), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT94), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n597), .A2(KEYINPUT94), .A3(new_n745), .A4(new_n608), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n748), .A2(new_n749), .B1(new_n652), .B2(new_n744), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n739), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n651), .B(KEYINPUT95), .Z(new_n752));
  OAI211_X1 g0552(.A(new_n672), .B(new_n751), .C1(new_n752), .C2(new_n750), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n674), .A2(new_n724), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT90), .Z(new_n755));
  OAI21_X1  g0555(.A(new_n736), .B1(new_n755), .B2(G77), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT91), .Z(new_n757));
  OAI21_X1  g0557(.A(new_n716), .B1(new_n679), .B2(new_n211), .ZN(new_n758));
  INV_X1    g0558(.A(new_n685), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n680), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n691), .A2(new_n706), .B1(new_n694), .B2(new_n688), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n360), .B1(new_n697), .B2(new_n206), .ZN(new_n762));
  NOR4_X1   g0562(.A1(new_n758), .A2(new_n760), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n702), .B2(new_n712), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(G107), .B2(new_n707), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT92), .B(G143), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n700), .A2(new_n766), .B1(new_n685), .B2(G150), .ZN(new_n767));
  INV_X1    g0567(.A(G137), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n767), .B1(new_n768), .B2(new_n691), .C1(new_n697), .C2(new_n718), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT93), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT34), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n348), .B1(new_n705), .B2(new_n217), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n222), .A2(new_n708), .B1(new_n679), .B2(new_n209), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(G132), .C2(new_n689), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n765), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n757), .B1(new_n745), .B2(new_n726), .C1(new_n675), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n753), .A2(new_n776), .ZN(G384));
  INV_X1    g0577(.A(new_n605), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n374), .B1(new_n377), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT37), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(new_n780), .A3(new_n371), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n350), .A2(new_n355), .ZN(new_n782));
  NOR2_X1   g0582(.A1(KEYINPUT98), .A2(KEYINPUT16), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n350), .B(new_n355), .C1(KEYINPUT98), .C2(KEYINPUT16), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n784), .A2(new_n260), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n605), .B1(new_n786), .B2(new_n368), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n786), .A2(new_n368), .B1(new_n375), .B2(new_n376), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n787), .A2(new_n788), .A3(new_n369), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n781), .B1(new_n789), .B2(new_n780), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n380), .A2(new_n787), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n790), .A2(new_n791), .A3(KEYINPUT38), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT38), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n374), .A2(new_n778), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n583), .B2(new_n580), .ZN(new_n795));
  AND3_X1   g0595(.A1(new_n779), .A2(new_n780), .A3(new_n371), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n780), .B1(new_n779), .B2(new_n371), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n793), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n792), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT99), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n314), .A2(new_n608), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n324), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT97), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT97), .ZN(new_n806));
  INV_X1    g0606(.A(new_n803), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n326), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n808), .B2(new_n804), .ZN(new_n809));
  AND3_X1   g0609(.A1(new_n650), .A2(new_n745), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n802), .A2(KEYINPUT40), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n787), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n786), .A2(new_n368), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n377), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n812), .A2(new_n814), .A3(new_n371), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n796), .B1(KEYINPUT37), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n812), .B1(new_n583), .B2(new_n580), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n793), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n792), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n650), .A2(new_n819), .A3(new_n809), .A4(new_n745), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT40), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT100), .Z(new_n824));
  NAND2_X1  g0624(.A1(new_n402), .A2(new_n650), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G330), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT39), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n800), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n324), .A2(new_n325), .A3(new_n608), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(new_n828), .C2(new_n819), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n578), .A2(new_n579), .A3(new_n605), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n743), .B(KEYINPUT96), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n748), .B2(new_n749), .ZN(new_n836));
  INV_X1    g0636(.A(new_n809), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n834), .B1(new_n819), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n653), .A2(new_n659), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n402), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n586), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n839), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n827), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n261), .B2(new_n601), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT35), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n233), .B(new_n234), .C1(new_n437), .C2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(G116), .C1(new_n846), .C2(new_n437), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT36), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n232), .A2(new_n351), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n850), .A2(new_n713), .B1(G50), .B2(new_n209), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(G1), .A3(new_n600), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n845), .A2(new_n849), .A3(new_n852), .ZN(G367));
  INV_X1    g0653(.A(new_n622), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n453), .A2(new_n461), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT42), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n448), .A2(new_n607), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n449), .A2(new_n608), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n594), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n607), .B1(new_n862), .B2(new_n453), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT43), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n608), .B1(new_n496), .B2(new_n494), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n587), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n592), .B2(new_n865), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT101), .Z(new_n868));
  OAI22_X1  g0668(.A1(new_n857), .A2(new_n863), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n620), .A2(new_n861), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n864), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n869), .B(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n627), .B(KEYINPUT41), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n861), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n624), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT44), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT44), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n624), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n622), .A2(new_n623), .A3(new_n861), .ZN(new_n883));
  XOR2_X1   g0683(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n622), .A2(new_n623), .A3(new_n861), .A4(new_n884), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n620), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n612), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n618), .A2(new_n619), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n621), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n892), .B2(new_n854), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n612), .B(new_n622), .C1(new_n891), .C2(new_n621), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI211_X1 g0695(.A(KEYINPUT44), .B(new_n861), .C1(new_n622), .C2(new_n623), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n880), .B1(new_n624), .B2(new_n877), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n886), .A2(new_n887), .ZN(new_n899));
  INV_X1    g0699(.A(new_n620), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n664), .A2(new_n889), .A3(new_n895), .A4(new_n901), .ZN(new_n902));
  AOI211_X1 g0702(.A(KEYINPUT103), .B(new_n876), .C1(new_n902), .C2(new_n664), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT103), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n889), .A2(new_n901), .ZN(new_n905));
  INV_X1    g0705(.A(new_n895), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n664), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n904), .B1(new_n907), .B2(new_n875), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n671), .A2(G1), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n874), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n766), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n222), .A2(new_n697), .B1(new_n691), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n704), .A2(G68), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n712), .B2(new_n253), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n914), .B(new_n916), .C1(new_n685), .C2(new_n717), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n273), .B1(new_n679), .B2(new_n713), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT104), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n918), .A2(new_n919), .B1(G137), .B2(new_n689), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n921), .B1(new_n919), .B2(new_n918), .C1(new_n217), .C2(new_n708), .ZN(new_n922));
  INV_X1    g0722(.A(G317), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n688), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT46), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n708), .A2(new_n925), .A3(new_n206), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n348), .B1(new_n685), .B2(G294), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n927), .B1(new_n680), .B2(new_n697), .C1(new_n706), .C2(new_n712), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n926), .B(new_n928), .C1(G107), .C2(new_n704), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n925), .B1(new_n708), .B2(new_n206), .ZN(new_n930));
  AOI22_X1  g0730(.A1(G311), .A2(new_n692), .B1(new_n678), .B2(G97), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n922), .B1(new_n924), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n674), .ZN(new_n935));
  INV_X1    g0735(.A(new_n731), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n728), .B1(new_n227), .B2(new_n384), .C1(new_n243), .C2(new_n936), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n935), .A2(new_n736), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n868), .A2(new_n727), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT105), .B1(new_n912), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n664), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n900), .B1(new_n898), .B2(new_n899), .ZN(new_n944));
  NOR4_X1   g0744(.A1(new_n888), .A2(new_n896), .A3(new_n897), .A4(new_n620), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n943), .B1(new_n946), .B2(new_n895), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT103), .B1(new_n947), .B2(new_n876), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n907), .A2(new_n904), .A3(new_n875), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(new_n911), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n873), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT105), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n940), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n942), .A2(new_n953), .ZN(G387));
  AOI21_X1  g0754(.A(new_n628), .B1(new_n664), .B2(new_n895), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(new_n664), .C2(new_n895), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n382), .A2(new_n222), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT50), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n209), .A2(new_n307), .ZN(new_n961));
  NOR4_X1   g0761(.A1(new_n960), .A2(G45), .A3(new_n961), .A4(new_n630), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n731), .B1(new_n240), .B2(new_n418), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n273), .A2(new_n630), .A3(new_n227), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n227), .A2(G107), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n728), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n348), .B1(new_n697), .B2(new_n209), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n707), .A2(new_n214), .B1(G150), .B2(new_n689), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT106), .Z(new_n970));
  AOI211_X1 g0770(.A(new_n968), .B(new_n970), .C1(G159), .C2(new_n692), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n685), .A2(new_n382), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G50), .A2(new_n700), .B1(new_n678), .B2(G97), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n472), .A2(new_n704), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G317), .A2(new_n700), .B1(new_n685), .B2(G311), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n692), .A2(G322), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(new_n706), .C2(new_n697), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT48), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n680), .B2(new_n705), .C1(new_n702), .C2(new_n708), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT49), .Z(new_n981));
  AOI21_X1  g0781(.A(new_n348), .B1(G326), .B2(new_n689), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n679), .B2(new_n206), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n975), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT107), .Z(new_n985));
  OAI21_X1  g0785(.A(new_n967), .B1(new_n985), .B2(new_n675), .ZN(new_n986));
  INV_X1    g0786(.A(new_n727), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n891), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n986), .A2(new_n672), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n910), .B2(new_n895), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n958), .A2(new_n990), .ZN(G393));
  INV_X1    g0791(.A(KEYINPUT109), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n944), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n905), .B2(new_n992), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n664), .A2(new_n895), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n627), .B(new_n902), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n679), .A2(new_n204), .B1(new_n697), .B2(new_n702), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n273), .B(new_n998), .C1(G322), .C2(new_n689), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n712), .A2(new_n694), .B1(new_n923), .B2(new_n691), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT52), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(new_n680), .C2(new_n708), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G303), .B2(new_n685), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n206), .B2(new_n705), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT110), .ZN(new_n1005));
  INV_X1    g0805(.A(G159), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n712), .A2(new_n1006), .B1(new_n253), .B2(new_n691), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT51), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n348), .B1(new_n688), .B2(new_n913), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n705), .A2(new_n307), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G68), .C2(new_n707), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n685), .A2(G50), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n697), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1013), .A2(new_n382), .B1(new_n678), .B2(G87), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n675), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n861), .A2(new_n987), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n728), .B1(new_n219), .B2(new_n227), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n250), .B2(new_n731), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n1016), .A2(new_n672), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n994), .B2(new_n910), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n997), .A2(new_n1021), .ZN(G390));
  NAND3_X1  g0822(.A1(new_n402), .A2(G330), .A3(new_n650), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n841), .A2(new_n586), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n650), .A2(G330), .A3(new_n745), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n837), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n650), .A2(G330), .A3(new_n809), .A4(new_n745), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n608), .B(new_n745), .C1(new_n655), .C2(new_n657), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n835), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n836), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1027), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT111), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(KEYINPUT111), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n829), .B1(new_n828), .B2(new_n819), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n748), .A2(new_n749), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n1029), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n809), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1039), .B1(new_n1042), .B2(new_n830), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n830), .B1(new_n1030), .B2(new_n837), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n800), .B(KEYINPUT99), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1036), .B(new_n1037), .C1(new_n1043), .C2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1038), .B1(new_n838), .B2(new_n831), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n802), .B(new_n830), .C1(new_n837), .C2(new_n1030), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1048), .A2(KEYINPUT111), .A3(new_n1035), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1034), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1047), .A2(new_n1034), .A3(new_n1050), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n627), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n910), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT54), .B(G143), .Z(new_n1057));
  AOI22_X1  g0857(.A1(new_n1013), .A2(new_n1057), .B1(new_n704), .B2(G159), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n768), .B2(new_n759), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT112), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n707), .A2(G150), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT53), .Z(new_n1062));
  AOI21_X1  g0862(.A(new_n360), .B1(new_n700), .B2(G132), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G125), .B2(new_n689), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n692), .A2(G128), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n222), .C2(new_n679), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT113), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n679), .A2(new_n209), .B1(new_n697), .B2(new_n219), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G294), .B2(new_n689), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n206), .B2(new_n712), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1010), .B(new_n1071), .C1(G283), .C2(new_n692), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n685), .A2(G107), .ZN(new_n1073));
  AND4_X1   g0873(.A1(new_n360), .A2(new_n1072), .A3(new_n710), .A4(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n674), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n755), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n672), .B1(new_n1076), .B2(new_n257), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1075), .B(new_n1077), .C1(new_n1039), .C2(new_n726), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT114), .B1(new_n1056), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n911), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT114), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1078), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1054), .B1(new_n1079), .B2(new_n1083), .ZN(G378));
  NAND4_X1  g0884(.A1(new_n650), .A2(KEYINPUT40), .A3(new_n809), .A4(new_n745), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n822), .B(G330), .C1(new_n1045), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n296), .A2(new_n329), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1087), .B(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n267), .A2(new_n778), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1090), .B(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n811), .A2(new_n1093), .A3(G330), .A4(new_n822), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1095), .A2(new_n839), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n839), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n841), .A2(new_n586), .A3(new_n1023), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1051), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT57), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1099), .B(KEYINPUT57), .C1(new_n1051), .C2(new_n1100), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n627), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n839), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1095), .A2(new_n839), .A3(new_n1096), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n910), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT116), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1094), .A2(new_n726), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n283), .A2(new_n285), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n345), .B(new_n1113), .C1(new_n708), .C2(new_n713), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n915), .B1(new_n680), .B2(new_n688), .C1(new_n712), .C2(new_n204), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n472), .B2(new_n1013), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n217), .B2(new_n679), .C1(new_n206), .C2(new_n691), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1114), .B(new_n1117), .C1(G97), .C2(new_n685), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT58), .Z(new_n1119));
  NAND2_X1  g0919(.A1(new_n269), .A2(new_n282), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT115), .ZN(new_n1121));
  AOI211_X1 g0921(.A(G50), .B(new_n1121), .C1(new_n1113), .C2(new_n345), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G137), .A2(new_n1013), .B1(new_n692), .B2(G125), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n707), .A2(new_n1057), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n700), .A2(G128), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n685), .A2(G132), .B1(G150), .B2(new_n704), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT59), .Z(new_n1128));
  NAND2_X1  g0928(.A1(new_n689), .A2(G124), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1121), .B(new_n1129), .C1(new_n679), .C2(new_n718), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1122), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n675), .B1(new_n1119), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n755), .A2(G50), .ZN(new_n1134));
  OR4_X1    g0934(.A1(new_n672), .A2(new_n1112), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1110), .A2(new_n1111), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1111), .B1(new_n1110), .B2(new_n1135), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1105), .A2(new_n1138), .ZN(G375));
  NOR3_X1   g0939(.A1(new_n809), .A2(G13), .A3(G33), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n679), .A2(new_n307), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G107), .A2(new_n1013), .B1(new_n700), .B2(G283), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n206), .B2(new_n759), .C1(new_n706), .C2(new_n688), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(G97), .C2(new_n707), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n692), .A2(G294), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n360), .A3(new_n974), .A4(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT118), .Z(new_n1147));
  NOR2_X1   g0947(.A1(new_n679), .A2(new_n217), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G150), .A2(new_n1013), .B1(new_n700), .B2(G137), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1006), .B2(new_n708), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(G50), .C2(new_n704), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n685), .A2(new_n1057), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n692), .A2(G132), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n345), .B1(G128), .B2(new_n689), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n675), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n755), .A2(G68), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1140), .A2(new_n672), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1041), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1031), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n910), .B(KEYINPUT117), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1158), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n875), .B1(new_n1161), .B2(new_n1024), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1034), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(G381));
  INV_X1    g0966(.A(G390), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n942), .A2(new_n953), .A3(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n958), .A2(new_n737), .A3(new_n673), .A4(new_n990), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1168), .A2(G384), .A3(G381), .A4(new_n1169), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT119), .Z(new_n1171));
  NOR2_X1   g0971(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1054), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1105), .A2(new_n1138), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(G407));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n606), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(G407), .A2(G213), .A3(new_n1176), .ZN(G409));
  INV_X1    g0977(.A(KEYINPUT61), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1160), .A2(new_n1100), .A3(KEYINPUT60), .A4(new_n1031), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1034), .A2(new_n627), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT60), .B1(new_n1181), .B2(new_n1100), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1163), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(G384), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(G384), .B(new_n1163), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n606), .A2(G213), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT120), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT121), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1185), .A2(new_n1192), .A3(new_n1186), .A4(new_n1189), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(G2897), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1191), .A2(G2897), .A3(new_n1188), .A4(new_n1193), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1105), .A2(G378), .A3(new_n1138), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1099), .A2(new_n1162), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1135), .B(new_n1200), .C1(new_n1101), .C2(new_n876), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1173), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1188), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1178), .B1(new_n1198), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n1207));
  AND4_X1   g1007(.A1(new_n1187), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1204), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT124), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n1169), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n952), .B1(new_n951), .B2(new_n940), .ZN(new_n1216));
  AOI211_X1 g1016(.A(KEYINPUT105), .B(new_n941), .C1(new_n950), .C2(new_n873), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1216), .A2(new_n1217), .A3(G390), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1167), .B1(new_n951), .B2(new_n940), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1215), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n912), .A2(new_n941), .A3(G390), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1221), .A2(new_n1215), .A3(new_n1219), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1213), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1215), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1219), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1168), .B2(new_n1226), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1227), .A2(KEYINPUT123), .A3(new_n1222), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1212), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1220), .A2(new_n1213), .A3(new_n1223), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT123), .B1(new_n1227), .B2(new_n1222), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(KEYINPUT124), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1211), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1204), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT63), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1203), .A2(new_n1236), .A3(new_n1206), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1234), .B(new_n1235), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT125), .B1(new_n1233), .B2(new_n1240), .ZN(new_n1241));
  OR3_X1    g1041(.A1(new_n1204), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1230), .A2(new_n1231), .A3(KEYINPUT124), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT124), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT125), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n1239), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1241), .A2(new_n1247), .ZN(G405));
  OAI21_X1  g1048(.A(KEYINPUT127), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G375), .A2(new_n1173), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1199), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(KEYINPUT126), .A3(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1206), .B(KEYINPUT126), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n1250), .A3(new_n1199), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1249), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1224), .A2(new_n1228), .A3(KEYINPUT127), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1256), .B(new_n1257), .ZN(G402));
endmodule


