//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936;
  XOR2_X1   g000(.A(KEYINPUT67), .B(G119), .Z(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(G116), .B2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G113), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  AND4_X1   g012(.A1(new_n194), .A2(new_n196), .A3(new_n198), .A4(G128), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n197), .B2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n196), .A2(new_n198), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(KEYINPUT65), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n199), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(G134), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n214), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n214), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n214), .A2(G137), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n212), .A2(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n209), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT0), .A4(G128), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n203), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n216), .A2(new_n218), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n227), .B1(new_n229), .B2(new_n219), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n193), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n234), .B(new_n237), .C1(new_n224), .C2(new_n230), .ZN(new_n238));
  INV_X1    g052(.A(new_n199), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n202), .A2(new_n203), .A3(new_n200), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT65), .B1(new_n206), .B2(new_n207), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n219), .A2(new_n222), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n227), .ZN(new_n245));
  INV_X1    g059(.A(new_n219), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n217), .B1(new_n216), .B2(new_n218), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n244), .A2(new_n248), .A3(new_n235), .A4(new_n236), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n192), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n233), .B1(new_n251), .B2(KEYINPUT68), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT31), .ZN(new_n253));
  NOR2_X1   g067(.A1(G237), .A2(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G210), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n255), .B(KEYINPUT27), .Z(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(G101), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n256), .B(new_n257), .Z(new_n258));
  AOI21_X1  g072(.A(new_n193), .B1(new_n238), .B2(new_n249), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n252), .A2(new_n253), .A3(new_n258), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT70), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n232), .B1(new_n259), .B2(new_n260), .ZN(new_n264));
  AOI211_X1 g078(.A(KEYINPUT68), .B(new_n193), .C1(new_n238), .C2(new_n249), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n253), .A4(new_n258), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n270), .A2(new_n258), .A3(new_n261), .A4(new_n232), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n252), .A2(new_n273), .A3(new_n258), .A4(new_n261), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(KEYINPUT31), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n258), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n231), .B(new_n192), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n233), .A2(KEYINPUT28), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n269), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n287));
  OR3_X1    g101(.A1(new_n279), .A2(new_n276), .A3(new_n280), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n276), .B1(new_n264), .B2(new_n265), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n288), .B2(new_n290), .ZN(new_n293));
  OAI21_X1  g107(.A(G472), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n284), .A2(new_n295), .A3(new_n285), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n287), .A2(new_n294), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n187), .B2(G128), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n189), .A2(new_n201), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n187), .B2(new_n201), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n302), .B2(new_n299), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT24), .B(G110), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  OAI22_X1  g119(.A1(new_n303), .A2(G110), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G125), .B(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT16), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n309), .A2(KEYINPUT16), .A3(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(G146), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n195), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n303), .A2(G110), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n302), .A2(new_n305), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n308), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n195), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n311), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT73), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT22), .B(G137), .ZN(new_n326));
  INV_X1    g140(.A(G953), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n327), .A2(G221), .A3(G234), .ZN(new_n328));
  XOR2_X1   g142(.A(new_n326), .B(new_n328), .Z(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n320), .B2(new_n321), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n332), .A3(new_n292), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n331), .B1(new_n325), .B2(new_n329), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT25), .A3(new_n292), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G217), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(G234), .B2(new_n292), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(G902), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT74), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G107), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G104), .ZN(new_n348));
  NOR2_X1   g162(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G104), .ZN(new_n353));
  OAI22_X1  g167(.A1(new_n353), .A2(G107), .B1(KEYINPUT75), .B2(KEYINPUT3), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(G107), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G101), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n351), .ZN(new_n358));
  OAI211_X1 g172(.A(G104), .B(new_n347), .C1(new_n358), .C2(new_n349), .ZN(new_n359));
  INV_X1    g173(.A(G101), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n354), .A4(new_n355), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n361), .A3(KEYINPUT4), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n363), .B(G101), .C1(new_n352), .C2(new_n356), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n190), .A2(new_n191), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT83), .B1(new_n188), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n187), .A2(new_n367), .A3(new_n370), .A4(G116), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(G113), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n190), .A2(new_n367), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n366), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n348), .A2(new_n355), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n361), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n361), .B2(new_n377), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n193), .A2(new_n365), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G122), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI221_X1 g198(.A(new_n382), .B1(new_n374), .B2(new_n380), .C1(new_n193), .C2(new_n365), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT6), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n209), .A2(new_n309), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n245), .B2(new_n309), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n227), .A2(KEYINPUT84), .A3(G125), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n327), .A2(G224), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n393), .B(new_n394), .Z(new_n395));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT7), .B1(new_n394), .B2(KEYINPUT85), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(KEYINPUT85), .B2(new_n394), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n389), .A2(new_n391), .A3(new_n392), .A4(new_n398), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(KEYINPUT86), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(KEYINPUT86), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n190), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n366), .B1(new_n372), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n361), .A2(new_n377), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n382), .B(KEYINPUT8), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(new_n409), .C1(new_n407), .C2(new_n374), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n394), .A2(KEYINPUT7), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n393), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n402), .A2(new_n410), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n385), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n400), .A2(new_n401), .B1(new_n393), .B2(new_n412), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n411), .B1(new_n416), .B2(new_n410), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n396), .B(new_n292), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G210), .B1(G237), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n410), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT87), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n414), .A3(new_n385), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n424), .A2(new_n292), .A3(new_n419), .A4(new_n396), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G214), .B1(G237), .B2(G902), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT81), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  INV_X1    g245(.A(G227), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(G953), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n431), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT10), .B(new_n242), .C1(new_n378), .C2(new_n379), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n194), .B1(G143), .B2(new_n195), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n201), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n205), .A2(KEYINPUT76), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n203), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n361), .B(new_n377), .C1(new_n441), .C2(new_n199), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT10), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n362), .A2(new_n245), .A3(new_n364), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n436), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n247), .B2(new_n246), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n246), .A2(new_n247), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n436), .A2(new_n448), .A3(new_n444), .A4(new_n445), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n435), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n435), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT79), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT79), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n454), .A3(new_n435), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n209), .A2(new_n406), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n448), .B1(new_n442), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(KEYINPUT12), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n459));
  AOI211_X1 g273(.A(new_n459), .B(new_n448), .C1(new_n442), .C2(new_n456), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n453), .A2(new_n455), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n451), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G469), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n292), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT78), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n449), .A2(new_n435), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n447), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n449), .B1(new_n458), .B2(new_n460), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n434), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n466), .B1(new_n471), .B2(new_n464), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n447), .A2(new_n467), .B1(new_n469), .B2(new_n434), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT78), .B(G469), .C1(new_n473), .C2(G902), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G221), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT9), .B(G234), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n478), .B2(new_n292), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT80), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n483), .A3(new_n480), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n430), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n318), .ZN(new_n486));
  INV_X1    g300(.A(G237), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n327), .A3(G214), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n197), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n254), .A2(G143), .A3(G214), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT17), .A3(G131), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(G131), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n486), .B(new_n492), .C1(KEYINPUT17), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(KEYINPUT18), .A3(G131), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT89), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n491), .B1(KEYINPUT18), .B2(G131), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n307), .B(KEYINPUT90), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G146), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n497), .B1(new_n499), .B2(new_n312), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(G113), .B(G122), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(new_n353), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n307), .A2(KEYINPUT19), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n307), .B(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n507), .B2(KEYINPUT19), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n311), .B(new_n493), .C1(new_n508), .C2(G146), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n503), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT91), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n501), .A2(new_n509), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n503), .ZN(new_n515));
  NOR2_X1   g329(.A1(G475), .A2(G902), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n513), .B1(new_n514), .B2(new_n503), .ZN(new_n520));
  NOR3_X1   g334(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n197), .A2(G128), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n201), .A2(G143), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(new_n214), .ZN(new_n527));
  XNOR2_X1  g341(.A(G116), .B(G122), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G107), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G116), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT14), .A3(G122), .ZN(new_n533));
  OAI211_X1 g347(.A(G107), .B(new_n533), .C1(new_n529), .C2(KEYINPUT14), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n527), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n201), .A2(G143), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n536), .B1(new_n537), .B2(KEYINPUT13), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n524), .A2(KEYINPUT93), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n540), .A3(new_n525), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n541), .A2(KEYINPUT94), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n541), .A2(KEYINPUT94), .B1(KEYINPUT13), .B2(new_n537), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n214), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n526), .A2(new_n214), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n528), .A2(new_n347), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n545), .B1(new_n530), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n535), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n477), .A2(new_n339), .A3(G953), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n535), .B(new_n549), .C1(new_n544), .C2(new_n547), .ZN(new_n552));
  AOI21_X1  g366(.A(G902), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT15), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(G478), .ZN(new_n556));
  INV_X1    g370(.A(G478), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n553), .A2(KEYINPUT15), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G475), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n503), .B1(new_n494), .B2(new_n501), .ZN(new_n561));
  OR3_X1    g375(.A1(new_n504), .A2(new_n561), .A3(KEYINPUT92), .ZN(new_n562));
  AOI21_X1  g376(.A(G902), .B1(new_n561), .B2(KEYINPUT92), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n523), .A2(new_n559), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G952), .ZN(new_n567));
  AOI211_X1 g381(.A(G953), .B(new_n567), .C1(G234), .C2(G237), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT21), .B(G898), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT95), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n292), .B(new_n327), .C1(G234), .C2(G237), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n298), .A2(new_n346), .A3(new_n485), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G101), .ZN(G3));
  AOI21_X1  g390(.A(new_n345), .B1(new_n482), .B2(new_n484), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n282), .A2(new_n292), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n578), .A2(G472), .B1(new_n283), .B2(new_n282), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n430), .A2(new_n573), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n517), .A2(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(new_n564), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n551), .A2(new_n552), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n551), .A2(KEYINPUT96), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT33), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n551), .B(new_n552), .C1(KEYINPUT96), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(G478), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n557), .A2(new_n292), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n553), .B2(new_n557), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n581), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n580), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT34), .B(G104), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  AOI21_X1  g411(.A(KEYINPUT97), .B1(new_n517), .B2(new_n518), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n517), .B2(new_n518), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n517), .A2(new_n518), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n564), .B1(new_n600), .B2(KEYINPUT97), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n559), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n581), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n580), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n329), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n320), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n343), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n341), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n485), .A2(new_n574), .A3(new_n579), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT37), .B(G110), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G12));
  XOR2_X1   g430(.A(KEYINPUT98), .B(G900), .Z(new_n617));
  AOI21_X1  g431(.A(new_n568), .B1(new_n572), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n604), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n428), .B1(new_n421), .B2(new_n425), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n475), .A2(new_n483), .A3(new_n480), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n483), .B1(new_n475), .B2(new_n480), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n621), .B(new_n613), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n298), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G128), .ZN(G30));
  AND2_X1   g441(.A1(new_n421), .A2(new_n425), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT38), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n523), .A2(new_n565), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n429), .A3(new_n603), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n613), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n272), .A2(new_n274), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n277), .A2(new_n258), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n292), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n287), .A2(new_n296), .A3(new_n297), .A4(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n639), .A2(KEYINPUT99), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n622), .A2(new_n623), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n618), .B(KEYINPUT39), .Z(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT40), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n639), .A2(KEYINPUT99), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT100), .B(G143), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G45));
  NAND2_X1  g463(.A1(new_n593), .A2(new_n619), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n298), .A2(new_n625), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  NAND2_X1  g467(.A1(new_n463), .A2(new_n292), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(G469), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n463), .B(new_n292), .C1(KEYINPUT101), .C2(new_n464), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n479), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n298), .A2(new_n594), .A3(new_n346), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT41), .B(G113), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G15));
  AND2_X1   g476(.A1(new_n298), .A2(new_n346), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n663), .A2(new_n605), .A3(new_n659), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n532), .ZN(G18));
  AND2_X1   g479(.A1(new_n659), .A2(new_n621), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n298), .A2(new_n574), .A3(new_n613), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G119), .ZN(G21));
  INV_X1    g482(.A(new_n573), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n656), .A2(new_n480), .A3(new_n669), .A4(new_n657), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n628), .A2(new_n670), .A3(new_n631), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n341), .A2(new_n672), .A3(new_n344), .ZN(new_n673));
  INV_X1    g487(.A(new_n340), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n335), .B2(new_n337), .ZN(new_n675));
  INV_X1    g489(.A(new_n344), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT103), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n578), .A2(G472), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n283), .B(KEYINPUT102), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n282), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n671), .A2(new_n678), .A3(new_n679), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G122), .ZN(G24));
  AND2_X1   g497(.A1(new_n679), .A2(new_n681), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n613), .A3(new_n651), .A4(new_n666), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G125), .ZN(G27));
  NOR2_X1   g500(.A1(new_n426), .A2(new_n428), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n465), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n471), .A2(new_n464), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n480), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n650), .A2(KEYINPUT42), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n346), .A2(new_n298), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n688), .A2(new_n650), .A3(new_n691), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n297), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT32), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n284), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n282), .A2(KEYINPUT104), .A3(KEYINPUT32), .A4(new_n283), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n697), .A2(new_n699), .A3(new_n294), .A4(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n701), .A2(new_n702), .A3(new_n678), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n701), .B2(new_n678), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n695), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n694), .B1(new_n705), .B2(KEYINPUT42), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G131), .ZN(G33));
  NAND3_X1  g521(.A1(new_n663), .A2(new_n620), .A3(new_n692), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n711));
  INV_X1    g525(.A(new_n592), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n583), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n592), .A2(KEYINPUT106), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n583), .A2(KEYINPUT43), .A3(new_n712), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n716), .A2(KEYINPUT107), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(KEYINPUT107), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n613), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n579), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(KEYINPUT44), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT108), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n473), .A2(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n473), .A2(KEYINPUT45), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(G469), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(G469), .A2(G902), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT46), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n689), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n727), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n479), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n731), .A2(new_n643), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n687), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(KEYINPUT44), .B2(new_n721), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n723), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G137), .ZN(G39));
  AND2_X1   g550(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n737));
  NOR2_X1   g551(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n731), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n731), .B2(new_n738), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n651), .A2(new_n345), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n740), .A2(new_n298), .A3(new_n688), .A4(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(G140), .Z(G42));
  NAND2_X1  g557(.A1(new_n658), .A2(KEYINPUT49), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n630), .A2(new_n479), .A3(new_n428), .A4(new_n592), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n678), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  OAI221_X1 g560(.A(new_n629), .B1(KEYINPUT49), .B2(new_n658), .C1(new_n746), .C2(KEYINPUT110), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(KEYINPUT110), .B2(new_n746), .ZN(new_n748));
  INV_X1    g562(.A(new_n638), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n703), .A2(new_n704), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n719), .A2(new_n568), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n687), .A2(new_n659), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT48), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(new_n678), .A3(new_n684), .ZN(new_n758));
  INV_X1    g572(.A(new_n666), .ZN(new_n759));
  OAI211_X1 g573(.A(G952), .B(new_n327), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n346), .A2(new_n749), .A3(new_n568), .A4(new_n754), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n593), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n629), .A2(new_n428), .A3(new_n659), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT116), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n758), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT50), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n583), .A3(new_n592), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n684), .A2(new_n613), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n755), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n758), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n656), .A2(new_n479), .A3(new_n657), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n740), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n774), .A3(new_n687), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n740), .B(KEYINPUT114), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n773), .B(KEYINPUT115), .Z(new_n778));
  AOI211_X1 g592(.A(new_n688), .B(new_n758), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n771), .A2(new_n779), .ZN(new_n780));
  OAI221_X1 g594(.A(new_n763), .B1(new_n771), .B2(new_n776), .C1(new_n780), .C2(KEYINPUT51), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n592), .B1(new_n582), .B2(new_n564), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n566), .A2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n621), .A3(new_n669), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n577), .A2(new_n785), .A3(new_n579), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n614), .A2(new_n786), .A3(new_n682), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n575), .A3(new_n660), .A4(new_n667), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n664), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n613), .A2(new_n559), .A3(new_n602), .A4(new_n619), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n641), .A3(new_n688), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n769), .A2(new_n695), .B1(new_n791), .B2(new_n298), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n708), .A2(new_n792), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n628), .A2(new_n691), .A3(new_n631), .A4(new_n618), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n638), .A2(new_n633), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n626), .A2(new_n652), .A3(new_n795), .A4(new_n685), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(KEYINPUT111), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n789), .A2(new_n706), .A3(new_n793), .A4(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n796), .A2(new_n797), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n796), .A2(new_n797), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT111), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n782), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n800), .B2(new_n801), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n626), .A2(new_n652), .A3(new_n685), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(KEYINPUT52), .A3(new_n795), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n796), .A2(new_n797), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(KEYINPUT112), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n789), .A2(new_n706), .A3(new_n793), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n803), .B1(new_n812), .B2(new_n782), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT54), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n807), .A2(new_n815), .A3(new_n808), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n811), .A2(KEYINPUT53), .A3(new_n816), .A4(new_n798), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n789), .A2(new_n706), .A3(new_n793), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n805), .B2(new_n809), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n817), .B(new_n818), .C1(new_n820), .C2(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n814), .A2(KEYINPUT113), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n813), .A2(new_n823), .A3(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n781), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(G952), .A2(G953), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n750), .B1(new_n825), .B2(new_n826), .ZN(G75));
  NAND2_X1  g641(.A1(new_n567), .A2(G953), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT118), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT119), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n395), .B(KEYINPUT55), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n810), .B2(new_n811), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n799), .A2(new_n802), .A3(new_n782), .ZN(new_n835));
  OAI211_X1 g649(.A(G210), .B(G902), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n386), .A2(new_n388), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT117), .Z(new_n839));
  AND3_X1   g653(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n833), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n837), .ZN(new_n843));
  INV_X1    g657(.A(new_n839), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n832), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n831), .B1(new_n842), .B2(new_n847), .ZN(G51));
  INV_X1    g662(.A(new_n829), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n812), .A2(new_n782), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n292), .B1(new_n850), .B2(new_n817), .ZN(new_n851));
  INV_X1    g665(.A(new_n726), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n851), .A2(KEYINPUT120), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT120), .B1(new_n851), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n818), .B1(new_n850), .B2(new_n817), .ZN(new_n856));
  INV_X1    g670(.A(new_n821), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n727), .B(KEYINPUT57), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n463), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n849), .B1(new_n855), .B2(new_n860), .ZN(G54));
  NAND3_X1  g675(.A1(new_n851), .A2(KEYINPUT58), .A3(G475), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n511), .A3(new_n515), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n511), .A2(new_n515), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n851), .A2(KEYINPUT58), .A3(G475), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n849), .B1(new_n863), .B2(new_n865), .ZN(G60));
  AND2_X1   g680(.A1(new_n586), .A2(new_n588), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n590), .B(KEYINPUT59), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n830), .B1(new_n858), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n868), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n822), .A2(new_n824), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n867), .B2(new_n872), .ZN(G63));
  OAI21_X1  g687(.A(new_n817), .B1(new_n820), .B2(KEYINPUT53), .ZN(new_n874));
  NAND2_X1  g688(.A1(G217), .A2(G902), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT60), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n336), .B(KEYINPUT121), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n874), .A2(new_n611), .A3(new_n876), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n830), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n879), .A2(KEYINPUT61), .A3(new_n830), .A4(new_n880), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(G66));
  AOI21_X1  g699(.A(new_n327), .B1(new_n570), .B2(G224), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT122), .ZN(new_n887));
  INV_X1    g701(.A(new_n789), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(new_n327), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n839), .B1(G898), .B2(new_n327), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT123), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n889), .B(new_n891), .ZN(G69));
  NAND2_X1  g706(.A1(new_n647), .A2(new_n806), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT62), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n742), .B1(new_n723), .B2(new_n734), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n687), .A2(new_n784), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n663), .A2(new_n642), .A3(new_n643), .A4(new_n896), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT124), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(G953), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n250), .B(new_n508), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(G900), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n905), .B2(new_n327), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n628), .A2(new_n631), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n751), .A2(new_n907), .A3(new_n732), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n895), .A2(new_n708), .A3(new_n806), .A4(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n706), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n906), .B1(new_n911), .B2(new_n327), .ZN(new_n912));
  OAI21_X1  g726(.A(G953), .B1(new_n432), .B2(new_n905), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n903), .B2(KEYINPUT125), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n904), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n904), .B2(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(G72));
  NAND2_X1  g731(.A1(new_n266), .A2(new_n276), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT126), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n266), .A2(new_n276), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(G472), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT63), .Z(new_n923));
  OAI21_X1  g737(.A(new_n829), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n900), .A2(new_n920), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n911), .A2(new_n919), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n927), .B2(new_n789), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n272), .A2(new_n289), .A3(new_n274), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n813), .A2(new_n923), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(KEYINPUT127), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n924), .ZN(new_n932));
  AOI22_X1  g746(.A1(new_n900), .A2(new_n920), .B1(new_n911), .B2(new_n919), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n930), .B(new_n932), .C1(new_n933), .C2(new_n888), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n931), .A2(new_n936), .ZN(G57));
endmodule


