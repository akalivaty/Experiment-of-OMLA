//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G77), .A2(G244), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G87), .A2(G250), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT66), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  AND3_X1   g0022(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n223));
  AOI21_X1  g0023(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n209), .B(new_n222), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G270), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT67), .B(G264), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n234), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT69), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  INV_X1    g0045(.A(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT68), .B(G87), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(new_n257), .B2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n203), .A2(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G150), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n226), .A2(G33), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n260), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n256), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n202), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n259), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT9), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n259), .A2(new_n266), .A3(new_n272), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(KEYINPUT71), .A3(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(G223), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n278), .A2(G1698), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G222), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n283), .B(new_n285), .C1(new_n286), .C2(new_n281), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n223), .B2(new_n224), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(new_n292), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n296), .B2(new_n292), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G226), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n291), .A2(G190), .A3(new_n295), .A4(new_n302), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n291), .A2(new_n295), .A3(new_n302), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n274), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT74), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n271), .A2(new_n308), .A3(new_n273), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n308), .B1(new_n271), .B2(new_n273), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT75), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT75), .ZN(new_n315));
  NOR4_X1   g0115(.A1(new_n310), .A2(new_n315), .A3(KEYINPUT10), .A4(new_n312), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n307), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n304), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(new_n270), .C1(G169), .C2(new_n304), .ZN(new_n320));
  INV_X1    g0120(.A(new_n263), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n264), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n256), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n268), .A2(new_n286), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n258), .A2(G77), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n284), .A2(G232), .B1(G107), .B2(new_n278), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n280), .A2(G238), .A3(new_n282), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n294), .B1(new_n331), .B2(new_n290), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n301), .A2(G244), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n328), .B1(new_n334), .B2(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n333), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(G179), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT73), .ZN(new_n339));
  INV_X1    g0139(.A(new_n328), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n334), .C2(new_n305), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n305), .B1(new_n332), .B2(new_n333), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT73), .B1(new_n342), .B2(new_n328), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT72), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n334), .A2(new_n345), .A3(G190), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT72), .B1(new_n336), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n338), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT76), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G33), .A3(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT3), .ZN(new_n356));
  INV_X1    g0156(.A(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n358), .A2(new_n359), .B1(new_n236), .B2(G1698), .ZN(new_n360));
  INV_X1    g0160(.A(G226), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n279), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n355), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n295), .B1(new_n363), .B2(new_n289), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n299), .A2(new_n300), .A3(new_n219), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT13), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n362), .B1(G232), .B2(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n367));
  INV_X1    g0167(.A(new_n355), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n294), .B1(new_n369), .B2(new_n290), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  INV_X1    g0171(.A(new_n300), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(G238), .A3(new_n298), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n366), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n370), .A2(KEYINPUT77), .A3(new_n371), .A4(new_n373), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(G200), .A3(new_n377), .ZN(new_n378));
  NOR4_X1   g0178(.A1(new_n202), .A2(KEYINPUT78), .A3(G20), .A4(G33), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT78), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n261), .B2(G50), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n382), .B1(new_n226), .B2(G68), .C1(new_n286), .C2(new_n264), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n256), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT11), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT11), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(new_n386), .A3(new_n256), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n258), .A2(G68), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n268), .A2(KEYINPUT12), .A3(new_n218), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT12), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n267), .B2(G68), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT79), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n388), .A2(new_n394), .A3(new_n389), .A4(new_n391), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n385), .A2(new_n387), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n366), .A2(new_n374), .A3(G190), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n378), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n376), .A2(G169), .A3(new_n377), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n401), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n376), .A2(G169), .A3(new_n377), .A4(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n366), .A2(new_n374), .A3(G179), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n396), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n398), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n317), .A2(new_n320), .A3(new_n350), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n358), .A2(new_n226), .A3(new_n359), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n226), .A4(new_n359), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n218), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G58), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n218), .ZN(new_n417));
  OAI21_X1  g0217(.A(G20), .B1(new_n417), .B2(new_n201), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n261), .A2(G159), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n410), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT7), .B1(new_n278), .B2(new_n226), .ZN(new_n422));
  INV_X1    g0222(.A(new_n414), .ZN(new_n423));
  OAI21_X1  g0223(.A(G68), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n420), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(new_n426), .A3(new_n256), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n263), .A2(new_n268), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n258), .A2(new_n321), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT81), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n427), .A2(new_n432), .A3(new_n428), .A4(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n296), .A2(G232), .A3(new_n292), .ZN(new_n435));
  NOR2_X1   g0235(.A1(G223), .A2(G1698), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n358), .B2(new_n359), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n361), .A2(G1698), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n437), .A2(new_n438), .B1(G33), .B2(G87), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n435), .B(new_n295), .C1(new_n439), .C2(new_n289), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT82), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n440), .A2(new_n441), .A3(G179), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n438), .B1(G223), .B2(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G87), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n289), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n435), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n445), .A2(new_n446), .A3(new_n294), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT82), .B1(new_n447), .B2(G169), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n318), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n442), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n434), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT18), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n440), .A2(G200), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n440), .A2(new_n347), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n454), .B2(new_n456), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT18), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n434), .A2(new_n462), .A3(new_n450), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n409), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT85), .B(G116), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n226), .A3(G33), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n226), .A2(G107), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n468), .B(KEYINPUT23), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n226), .B(G87), .C1(new_n276), .C2(new_n277), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n470), .A2(KEYINPUT22), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(KEYINPUT22), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n467), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT24), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n470), .B(KEYINPUT22), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n476), .A2(KEYINPUT24), .A3(new_n467), .A4(new_n469), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n256), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n357), .A2(G1), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n256), .A2(new_n268), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G107), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n267), .A2(G107), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n482), .B(KEYINPUT25), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  INV_X1    g0286(.A(G41), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT5), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT5), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G41), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n293), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(G264), .A3(new_n296), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G250), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT88), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n281), .A2(KEYINPUT88), .A3(G250), .A4(new_n279), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n281), .A2(G257), .A3(G1698), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G294), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n492), .B(new_n494), .C1(new_n501), .C2(new_n290), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G169), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n318), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n484), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n281), .A2(new_n226), .A3(G68), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n264), .B2(new_n246), .ZN(new_n510));
  AOI21_X1  g0310(.A(G20), .B1(new_n355), .B2(KEYINPUT19), .ZN(new_n511));
  NOR3_X1   g0311(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n508), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n513), .A2(new_n256), .B1(new_n268), .B2(new_n323), .ZN(new_n514));
  INV_X1    g0314(.A(new_n323), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n480), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n466), .A2(G33), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n219), .A2(new_n279), .ZN(new_n518));
  INV_X1    g0318(.A(G244), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G1698), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n518), .B(new_n520), .C1(new_n276), .C2(new_n277), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n289), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n257), .A2(G45), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT84), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n257), .A2(KEYINPUT84), .A3(G45), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n525), .A2(G250), .A3(new_n296), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n523), .A2(new_n293), .ZN(new_n529));
  OR3_X1    g0329(.A1(new_n522), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n514), .A2(new_n516), .B1(new_n530), .B2(new_n504), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n522), .A2(new_n528), .A3(new_n529), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n318), .ZN(new_n533));
  NOR4_X1   g0333(.A1(new_n522), .A2(new_n528), .A3(new_n347), .A4(new_n529), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(G200), .B2(new_n530), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n513), .A2(new_n256), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n323), .A2(new_n268), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n480), .A2(G87), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n531), .A2(new_n533), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n501), .A2(new_n290), .ZN(new_n541));
  INV_X1    g0341(.A(new_n492), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n541), .A2(new_n347), .A3(new_n542), .A4(new_n493), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n502), .B2(G200), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n544), .A2(new_n481), .A3(new_n483), .A4(new_n478), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n507), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n479), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n225), .A2(new_n267), .A3(new_n255), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G116), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n548), .A2(new_n549), .B1(new_n267), .B2(new_n466), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(KEYINPUT85), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G116), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(new_n226), .C1(G33), .C2(new_n246), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n256), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT20), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n225), .A2(new_n255), .B1(new_n554), .B2(G20), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n550), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G257), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n564));
  OAI211_X1 g0364(.A(G264), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n358), .A2(G303), .A3(new_n359), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n290), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n491), .A2(G270), .A3(new_n296), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT86), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n491), .A2(KEYINPUT86), .A3(G270), .A4(new_n296), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n568), .A2(new_n542), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(KEYINPUT21), .A3(G169), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n492), .B1(new_n567), .B2(new_n290), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n575), .A2(G179), .A3(new_n571), .A4(new_n572), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n563), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n573), .A2(G200), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n575), .A2(G190), .A3(new_n571), .A4(new_n572), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(new_n563), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT87), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n573), .A2(G169), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n563), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n466), .A2(new_n267), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n480), .B2(G116), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT20), .B1(new_n561), .B2(new_n557), .ZN(new_n590));
  AND4_X1   g0390(.A1(KEYINPUT20), .A2(new_n555), .A3(new_n256), .A4(new_n557), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(G169), .A3(new_n573), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n583), .B1(new_n593), .B2(new_n584), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n578), .B(new_n582), .C1(new_n587), .C2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n491), .A2(G257), .A3(new_n296), .ZN(new_n596));
  OAI211_X1 g0396(.A(G244), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT4), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n556), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n596), .B1(new_n602), .B2(new_n290), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n542), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  INV_X1    g0405(.A(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(KEYINPUT6), .A3(G97), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n246), .A2(new_n606), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G97), .A2(G107), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n607), .B1(new_n610), .B2(KEYINPUT6), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G20), .ZN(new_n612));
  OAI21_X1  g0412(.A(G107), .B1(new_n422), .B2(new_n423), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n261), .A2(G77), .ZN(new_n614));
  XOR2_X1   g0414(.A(new_n614), .B(KEYINPUT83), .Z(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n616), .A2(new_n256), .B1(new_n246), .B2(new_n268), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n480), .A2(G97), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n603), .A2(G190), .A3(new_n542), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n605), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n616), .A2(new_n256), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n268), .A2(new_n246), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n622), .A3(new_n618), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n604), .A2(new_n504), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n603), .A2(new_n318), .A3(new_n542), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n546), .A2(new_n595), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n465), .A2(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n406), .A2(new_n407), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n335), .A2(new_n337), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n398), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n461), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n450), .A2(new_n430), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(new_n462), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT90), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n634), .A2(KEYINPUT90), .A3(new_n636), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n317), .A3(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(new_n320), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT89), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n532), .B2(new_n305), .ZN(new_n644));
  INV_X1    g0444(.A(new_n534), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n530), .A2(KEYINPUT89), .A3(G200), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n539), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n531), .A2(new_n533), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n649), .A2(KEYINPUT26), .A3(new_n626), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  INV_X1    g0451(.A(new_n626), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n540), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n584), .B1(new_n585), .B2(new_n563), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT87), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n577), .B1(new_n656), .B2(new_n586), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n507), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n620), .A2(new_n626), .A3(new_n647), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n545), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n654), .A2(new_n660), .A3(new_n648), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n465), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n642), .A2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(G13), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G20), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n257), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT91), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT27), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(G213), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n592), .ZN(new_n674));
  MUX2_X1   g0474(.A(new_n657), .B(new_n595), .S(new_n674), .Z(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n484), .A2(new_n673), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n507), .B(new_n545), .C1(new_n678), .C2(KEYINPUT93), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n678), .A2(KEYINPUT93), .ZN(new_n680));
  OR3_X1    g0480(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT94), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT94), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n673), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n507), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n677), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n507), .A2(new_n673), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n657), .A2(new_n673), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n683), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  AND2_X1   g0492(.A1(new_n512), .A2(new_n549), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n207), .A2(new_n487), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n228), .B2(new_n694), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT95), .ZN(new_n698));
  INV_X1    g0498(.A(new_n648), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n620), .A2(new_n626), .A3(new_n647), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n657), .B2(new_n507), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n701), .B2(new_n545), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n673), .B1(new_n702), .B2(new_n654), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n698), .B1(new_n703), .B2(KEYINPUT29), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT26), .B1(new_n649), .B2(new_n626), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n652), .A2(new_n540), .A3(new_n651), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n660), .A2(new_n648), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .A3(new_n685), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n661), .A2(new_n685), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(KEYINPUT95), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n704), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n507), .A2(new_n540), .A3(new_n545), .ZN(new_n713));
  AOI211_X1 g0513(.A(new_n577), .B(new_n581), .C1(new_n656), .C2(new_n586), .ZN(new_n714));
  INV_X1    g0514(.A(new_n627), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n715), .A4(new_n685), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  AND4_X1   g0517(.A1(new_n568), .A2(new_n542), .A3(new_n571), .A4(new_n572), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(G179), .A3(new_n532), .A4(new_n603), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n717), .B1(new_n719), .B2(new_n503), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n603), .A2(new_n532), .ZN(new_n721));
  INV_X1    g0521(.A(new_n576), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n721), .A2(KEYINPUT30), .A3(new_n722), .A4(new_n502), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n494), .B1(new_n501), .B2(new_n290), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n542), .B1(new_n724), .B2(new_n603), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n318), .A3(new_n573), .A4(new_n530), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n720), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n727), .A2(new_n673), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n716), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(KEYINPUT31), .ZN(new_n731));
  OAI21_X1  g0531(.A(G330), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n712), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n697), .B1(new_n733), .B2(G1), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT96), .ZN(G364));
  NAND2_X1  g0535(.A1(new_n665), .A2(G45), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n694), .A2(G1), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n677), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G330), .B2(new_n676), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n278), .A2(new_n207), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT97), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n243), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G45), .B2(new_n228), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n281), .A2(new_n207), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n745), .B1(G116), .B2(new_n207), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n225), .B1(G20), .B2(new_n504), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT100), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n226), .A2(new_n318), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G200), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n755), .B1(new_n757), .B2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n757), .A2(new_n755), .A3(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT33), .B(G317), .Z(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n347), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n318), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n281), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n305), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G20), .A3(new_n347), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G283), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n756), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT98), .B1(new_n226), .B2(new_n318), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G311), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n770), .A2(G20), .A3(G190), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  INV_X1    g0582(.A(G329), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n776), .A2(G20), .A3(new_n318), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n781), .A2(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n775), .A2(new_n777), .A3(new_n764), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n757), .A2(new_n347), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n785), .B(new_n788), .C1(G326), .C2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n769), .A2(new_n773), .A3(new_n780), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n766), .A2(G97), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n761), .B2(new_n218), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT101), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n779), .A2(G77), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n771), .A2(new_n606), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n281), .B1(new_n786), .B2(new_n416), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(G50), .C2(new_n789), .ZN(new_n798));
  INV_X1    g0598(.A(new_n784), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT99), .B(G159), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n781), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n801), .A2(KEYINPUT32), .B1(new_n802), .B2(G87), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n794), .A2(new_n795), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n801), .A2(KEYINPUT32), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n791), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n737), .B(new_n754), .C1(new_n806), .C2(new_n749), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT102), .ZN(new_n808));
  INV_X1    g0608(.A(new_n752), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n676), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n740), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NAND3_X1  g0612(.A1(new_n661), .A2(new_n350), .A3(new_n685), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n338), .A2(new_n685), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n344), .A2(new_n349), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n673), .A2(new_n328), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n815), .B1(new_n818), .B2(new_n631), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n813), .B1(new_n703), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n732), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n737), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n344), .A2(new_n349), .B1(new_n328), .B2(new_n673), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n814), .B1(new_n824), .B2(new_n338), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n750), .ZN(new_n826));
  INV_X1    g0626(.A(new_n761), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G283), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n802), .A2(G107), .B1(new_n799), .B2(G311), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n779), .A2(new_n466), .ZN(new_n830));
  AND4_X1   g0630(.A1(new_n792), .A2(new_n828), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n786), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G294), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n789), .A2(G303), .B1(new_n772), .B2(G87), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n831), .A2(new_n278), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n779), .A2(new_n800), .B1(G137), .B2(new_n789), .ZN(new_n836));
  INV_X1    g0636(.A(G143), .ZN(new_n837));
  INV_X1    g0637(.A(G150), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n837), .B2(new_n786), .C1(new_n761), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT34), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n771), .A2(new_n218), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n767), .A2(new_n416), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(G132), .C2(new_n799), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n281), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n781), .A2(new_n202), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n835), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n749), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n749), .A2(new_n750), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n286), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n826), .A2(new_n738), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n823), .A2(new_n850), .ZN(G384));
  NAND2_X1  g0651(.A1(new_n430), .A2(KEYINPUT106), .ZN(new_n852));
  INV_X1    g0652(.A(new_n671), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT106), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n427), .A2(new_n854), .A3(new_n428), .A4(new_n429), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n852), .A2(new_n450), .A3(new_n855), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n455), .A2(new_n457), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n454), .B2(new_n456), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n434), .B2(new_n450), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n434), .A2(new_n853), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n462), .B1(new_n434), .B2(new_n450), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n447), .A2(KEYINPUT82), .A3(new_n318), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n441), .B1(new_n440), .B2(new_n504), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n440), .A2(G179), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI211_X1 g0671(.A(KEYINPUT18), .B(new_n871), .C1(new_n431), .C2(new_n433), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n458), .A2(new_n460), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n867), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n866), .B(KEYINPUT38), .C1(new_n874), .C2(new_n856), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n455), .A2(new_n457), .B1(new_n450), .B2(new_n430), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n864), .A2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .B1(new_n863), .B2(new_n864), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n864), .B1(new_n636), .B2(new_n461), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT109), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n630), .A2(new_n685), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n407), .A2(new_n673), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n630), .A2(new_n633), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n408), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n885), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n727), .A2(KEYINPUT108), .A3(new_n673), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT31), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT108), .B1(new_n727), .B2(new_n673), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n819), .B1(new_n730), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n875), .A2(new_n881), .A3(KEYINPUT109), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n884), .A2(new_n898), .A3(KEYINPUT40), .A4(new_n899), .ZN(new_n900));
  XOR2_X1   g0700(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n901));
  NOR2_X1   g0701(.A1(new_n867), .A2(new_n872), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n856), .B1(new_n902), .B2(new_n461), .ZN(new_n903));
  AOI22_X1  g0703(.A1(KEYINPUT37), .A2(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n903), .A2(new_n876), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n856), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n464), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n907), .B2(new_n866), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n727), .A2(new_n673), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n893), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n628), .B2(new_n685), .ZN(new_n912));
  INV_X1    g0712(.A(new_n895), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n893), .A3(new_n892), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n825), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n885), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n408), .A2(new_n889), .A3(new_n886), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n889), .B1(new_n408), .B2(new_n886), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n901), .B1(new_n909), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n900), .A2(new_n921), .A3(G330), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n912), .A2(new_n914), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n465), .A2(G330), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n900), .A2(new_n921), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n465), .A2(new_n923), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n636), .A2(new_n853), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n891), .B1(new_n814), .B2(new_n813), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n876), .B1(new_n903), .B2(new_n904), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n875), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n929), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n882), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n630), .A2(new_n673), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n931), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n928), .B(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n704), .A2(new_n465), .A3(new_n708), .A4(new_n711), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n642), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n257), .B2(new_n665), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n549), .B1(new_n611), .B2(KEYINPUT35), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n946), .B(new_n227), .C1(KEYINPUT35), .C2(new_n611), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT36), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n218), .A2(KEYINPUT103), .A3(G50), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT103), .B1(new_n218), .B2(G50), .ZN(new_n950));
  OAI21_X1  g0750(.A(G77), .B1(new_n416), .B2(new_n218), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n949), .B(new_n950), .C1(new_n228), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(G1), .A3(new_n664), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT104), .Z(new_n954));
  NAND3_X1  g0754(.A1(new_n945), .A2(new_n948), .A3(new_n954), .ZN(G367));
  NAND2_X1  g0755(.A1(new_n673), .A2(new_n623), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n715), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n652), .A2(new_n673), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n688), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n685), .A2(new_n539), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n699), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n649), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT110), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n961), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n683), .A2(new_n690), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT42), .B1(new_n968), .B2(new_n957), .ZN(new_n969));
  INV_X1    g0769(.A(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT42), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n689), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n969), .B1(new_n626), .B2(new_n673), .C1(new_n972), .C2(new_n957), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n967), .B(new_n975), .Z(new_n976));
  XOR2_X1   g0776(.A(new_n694), .B(KEYINPUT41), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n691), .A2(new_n959), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n691), .A2(new_n959), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n688), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n984), .A2(new_n985), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n968), .B1(new_n687), .B2(new_n690), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(new_n677), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n733), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT111), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(KEYINPUT111), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n978), .B1(new_n995), .B2(new_n733), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n736), .A2(G1), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n976), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n827), .A2(new_n800), .B1(G137), .B2(new_n799), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n278), .B1(new_n772), .B2(G77), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n789), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n999), .B(new_n1000), .C1(new_n837), .C2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n767), .A2(new_n218), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n786), .A2(new_n838), .B1(new_n416), .B2(new_n781), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n779), .A2(G50), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n771), .A2(new_n246), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OR3_X1    g0808(.A1(new_n781), .A2(new_n554), .A3(KEYINPUT46), .ZN(new_n1009));
  OAI21_X1  g0809(.A(KEYINPUT46), .B1(new_n781), .B2(new_n549), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1009), .A2(new_n1010), .B1(new_n779), .B2(G283), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n763), .B2(new_n761), .ZN(new_n1012));
  INV_X1    g0812(.A(G317), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n278), .B1(new_n1013), .B2(new_n784), .C1(new_n786), .C2(new_n782), .ZN(new_n1014));
  INV_X1    g0814(.A(G311), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1001), .A2(new_n1015), .B1(new_n767), .B2(new_n606), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1005), .A2(new_n1006), .B1(new_n1008), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT47), .Z(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n749), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n964), .A2(new_n809), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n234), .A2(new_n742), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1022), .B(new_n753), .C1(new_n207), .C2(new_n323), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n738), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n998), .A2(new_n1024), .ZN(G387));
  AOI22_X1  g0825(.A1(new_n779), .A2(G303), .B1(G322), .B2(new_n789), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n1013), .B2(new_n786), .C1(new_n761), .C2(new_n1015), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  INV_X1    g0828(.A(G283), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n767), .C1(new_n763), .C2(new_n781), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT49), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n281), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n799), .A2(G326), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n772), .A2(new_n466), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n786), .A2(new_n202), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n827), .A2(new_n321), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n278), .B1(new_n789), .B2(G159), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT114), .B(G150), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n799), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n766), .A2(new_n515), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G77), .B2(new_n802), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n1008), .C1(new_n218), .C2(new_n778), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1036), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n749), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n263), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT50), .B1(new_n263), .B2(G50), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n485), .A4(new_n693), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n218), .A2(new_n286), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n742), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT113), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n485), .B2(new_n239), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(G107), .B2(new_n207), .C1(new_n693), .C2(new_n747), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n753), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n684), .A2(new_n686), .A3(new_n752), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1047), .A2(new_n738), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n991), .A2(new_n997), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT112), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n694), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n992), .A2(KEYINPUT115), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n733), .B2(new_n991), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT115), .B1(new_n992), .B2(new_n1061), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1058), .B(new_n1060), .C1(new_n1063), .C2(new_n1064), .ZN(G393));
  OAI21_X1  g0865(.A(new_n992), .B1(new_n987), .B2(new_n988), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n995), .A2(new_n1066), .A3(new_n1061), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n960), .A2(new_n752), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1001), .A2(new_n1013), .B1(new_n1015), .B2(new_n786), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT52), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n763), .B2(new_n778), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n781), .A2(new_n1029), .B1(new_n787), .B2(new_n784), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1072), .A2(new_n796), .A3(new_n281), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT117), .Z(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n782), .B2(new_n761), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1071), .B(new_n1075), .C1(new_n466), .C2(new_n766), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n281), .B1(new_n784), .B2(new_n837), .C1(new_n781), .C2(new_n218), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G87), .B2(new_n772), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT116), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n767), .A2(new_n286), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n832), .A2(G159), .B1(G150), .B2(new_n789), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(new_n1081), .B2(KEYINPUT51), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n263), .B2(new_n778), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n761), .A2(new_n202), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1081), .A2(KEYINPUT51), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1079), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n749), .B1(new_n1076), .B2(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n753), .B1(new_n246), .B2(new_n207), .C1(new_n249), .C2(new_n743), .ZN(new_n1088));
  AND4_X1   g0888(.A1(new_n738), .A2(new_n1068), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n989), .B2(new_n997), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1067), .A2(new_n1090), .ZN(G390));
  NAND4_X1  g0891(.A1(new_n942), .A2(new_n320), .A3(new_n641), .A4(new_n924), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT118), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n813), .A2(new_n814), .ZN(new_n1095));
  INV_X1    g0895(.A(G330), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n920), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n732), .A2(new_n825), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(new_n919), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1095), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n919), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n707), .A2(new_n350), .A3(new_n685), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n891), .B1(new_n897), .B2(new_n1096), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n814), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n642), .A2(KEYINPUT118), .A3(new_n942), .A4(new_n924), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1094), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1102), .A2(new_n814), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n936), .B1(new_n1108), .B2(new_n919), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1109), .A2(new_n884), .A3(new_n899), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n936), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1095), .A2(new_n919), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1111), .A2(new_n1112), .B1(new_n935), .B2(new_n937), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1110), .A2(new_n1113), .B1(new_n1096), .B2(new_n920), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n935), .A2(new_n937), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n936), .B2(new_n930), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n884), .A3(new_n899), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1116), .A2(new_n919), .A3(new_n1098), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT119), .B1(new_n1107), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1094), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT119), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n1114), .A4(new_n1118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1107), .A2(new_n1119), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1120), .A2(new_n1061), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1115), .A2(new_n750), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT54), .B(G143), .Z(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n281), .B1(new_n202), .B2(new_n771), .C1(new_n778), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n827), .A2(G137), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n802), .A2(new_n1040), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT53), .Z(new_n1132));
  NAND2_X1  g0932(.A1(new_n799), .A2(G125), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n789), .A2(G128), .B1(new_n766), .B2(G159), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1129), .B(new_n1135), .C1(G132), .C2(new_n832), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1080), .B1(G87), .B2(new_n802), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(new_n278), .C1(new_n1029), .C2(new_n1001), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n784), .A2(new_n763), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n761), .A2(new_n606), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n841), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n778), .B2(new_n246), .C1(new_n549), .C2(new_n786), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n749), .B1(new_n1136), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n848), .A2(new_n263), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1126), .A2(new_n738), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1119), .A2(new_n997), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT120), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1119), .A2(KEYINPUT120), .A3(new_n997), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1125), .A2(new_n1146), .A3(new_n1151), .ZN(G378));
  NAND2_X1  g0952(.A1(new_n1094), .A2(new_n1106), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n1119), .B2(new_n1105), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n317), .A2(new_n320), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n270), .A3(new_n853), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n853), .A2(new_n270), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n317), .A2(new_n320), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1158), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n922), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1166), .A2(new_n900), .A3(new_n921), .A4(G330), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n939), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n940), .A3(new_n1169), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1156), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n694), .B1(new_n1155), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1168), .A2(new_n940), .A3(new_n1169), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n940), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT123), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT123), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1171), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1154), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1174), .B1(new_n1180), .B2(KEYINPUT57), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1167), .A2(new_n750), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n202), .B1(new_n276), .B2(G41), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n789), .A2(G125), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n838), .B2(new_n767), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n779), .A2(G137), .ZN(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n786), .C1(new_n781), .C2(new_n1128), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1185), .B(new_n1188), .C1(G132), .C2(new_n827), .ZN(new_n1189));
  XOR2_X1   g0989(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1190));
  AOI21_X1  g0990(.A(G33), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n772), .A2(new_n800), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G41), .B1(new_n799), .B2(G124), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n281), .B1(new_n827), .B2(G97), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n606), .B2(new_n786), .C1(new_n549), .C2(new_n1001), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n784), .A2(new_n1029), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n771), .A2(new_n416), .B1(new_n781), .B2(new_n286), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1197), .A2(new_n1003), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1200), .B(new_n487), .C1(new_n323), .C2(new_n778), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1183), .B1(new_n1194), .B2(new_n1195), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n749), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n848), .A2(new_n202), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1182), .A2(new_n738), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n997), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1181), .A2(new_n1210), .ZN(G375));
  NAND3_X1  g1011(.A1(new_n1153), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(new_n977), .A3(new_n1121), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n891), .A2(new_n750), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n827), .A2(new_n466), .B1(G303), .B2(new_n799), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n286), .B2(new_n771), .C1(new_n606), .C2(new_n778), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n781), .A2(new_n246), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1042), .A2(new_n278), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1001), .A2(new_n763), .B1(new_n1029), .B2(new_n786), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n761), .A2(new_n1128), .B1(new_n838), .B2(new_n778), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G137), .B2(new_n832), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n281), .B1(new_n771), .B2(new_n416), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT124), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n789), .A2(G132), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n802), .A2(G159), .B1(new_n799), .B2(G128), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G50), .B2(new_n766), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n749), .B1(new_n1220), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n848), .A2(new_n218), .ZN(new_n1230));
  AND4_X1   g1030(.A1(new_n738), .A2(new_n1214), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1105), .B2(new_n997), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1213), .A2(new_n1232), .ZN(G381));
  NOR2_X1   g1033(.A1(G375), .A2(G378), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n998), .A3(new_n1024), .ZN(new_n1237));
  OR2_X1    g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1237), .A2(G384), .A3(G381), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1235), .B1(new_n1239), .B2(KEYINPUT125), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(KEYINPUT125), .B2(new_n1239), .ZN(G407));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G343), .C2(new_n1235), .ZN(G409));
  XNOR2_X1  g1042(.A(G393), .B(new_n811), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1236), .A2(new_n998), .A3(new_n1024), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1236), .B1(new_n998), .B2(new_n1024), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G387), .A2(G390), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1243), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1237), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1155), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT57), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1061), .B1(new_n1253), .B2(new_n1154), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G378), .B(new_n1210), .C1(new_n1251), .C2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1181), .A2(KEYINPUT126), .A3(G378), .A4(new_n1210), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1180), .A2(new_n977), .B1(new_n997), .B2(new_n1252), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G378), .B1(new_n1260), .B2(new_n1207), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(G213), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G343), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1061), .B(new_n1121), .C1(new_n1212), .C2(new_n1267), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1212), .A2(new_n1267), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1270), .B2(new_n1232), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G384), .B(new_n1232), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1263), .A2(new_n1266), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1265), .A2(G2897), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G2897), .B(new_n1265), .C1(new_n1271), .C2(new_n1273), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1261), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1277), .B(new_n1278), .C1(new_n1279), .C2(new_n1265), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT62), .B1(new_n1275), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1274), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1279), .A2(new_n1265), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT62), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1282), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1250), .B1(new_n1281), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT63), .B1(new_n1289), .B2(new_n1284), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1250), .A2(KEYINPUT61), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1275), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1287), .A2(new_n1294), .ZN(G405));
  NAND3_X1  g1095(.A1(new_n1250), .A2(KEYINPUT127), .A3(new_n1274), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1274), .A2(KEYINPUT127), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1246), .A2(new_n1249), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G378), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1257), .A2(new_n1258), .B1(new_n1300), .B2(G375), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1296), .A2(new_n1301), .A3(new_n1298), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(G402));
endmodule


