// Benchmark "locked_c1908" written by ABC on Sat Dec 16 10:46:22 2023

module locked_c1908 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110,
    G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146,
    G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478,
    G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104,
    G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140,
    G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472,
    G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123, new_n124, new_n125, new_n126, new_n127, new_n128, new_n129,
    new_n130, new_n131, new_n132, new_n133, new_n134, new_n135, new_n136,
    new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n431, new_n432,
    new_n433, new_n434, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n476, new_n477, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n501, new_n503, new_n504, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n511, new_n512, new_n514,
    new_n515, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696;
  INV_X1    g000(.A(G902), .ZN(new_n123));
  INV_X1    g001(.A(G217), .ZN(new_n124));
  XNOR2_X1  g002(.A(G125), .B(G140), .ZN(new_n125));
  NAND2_X1  g003(.A1(new_n125), .A2(KEYINPUT16), .ZN(new_n126));
  INV_X1    g004(.A(G140), .ZN(new_n127));
  NAND2_X1  g005(.A1(new_n127), .A2(G125), .ZN(new_n128));
  OR2_X1    g006(.A1(new_n128), .A2(KEYINPUT16), .ZN(new_n129));
  NAND2_X1  g007(.A1(new_n126), .A2(new_n129), .ZN(new_n130));
  INV_X1    g008(.A(G146), .ZN(new_n131));
  NAND2_X1  g009(.A1(new_n130), .A2(new_n131), .ZN(new_n132));
  NAND3_X1  g010(.A1(new_n126), .A2(G146), .A3(new_n129), .ZN(new_n133));
  NAND2_X1  g011(.A1(new_n132), .A2(new_n133), .ZN(new_n134));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n135));
  XNOR2_X1  g013(.A(G119), .B(G128), .ZN(new_n136));
  NAND2_X1  g014(.A1(new_n135), .A2(new_n136), .ZN(new_n137));
  INV_X1    g015(.A(G119), .ZN(new_n138));
  NOR3_X1   g016(.A1(new_n138), .A2(KEYINPUT23), .A3(G128), .ZN(new_n139));
  AOI21_X1  g017(.A(new_n139), .B1(new_n136), .B2(KEYINPUT23), .ZN(new_n140));
  NAND2_X1  g018(.A1(new_n140), .A2(G110), .ZN(new_n141));
  NAND3_X1  g019(.A1(new_n134), .A2(new_n137), .A3(new_n141), .ZN(new_n142));
  XOR2_X1   g020(.A(KEYINPUT22), .B(G137), .Z(new_n143));
  INV_X1    g021(.A(G953), .ZN(new_n144));
  NAND3_X1  g022(.A1(new_n144), .A2(G221), .A3(G234), .ZN(new_n145));
  XNOR2_X1  g023(.A(new_n143), .B(new_n145), .ZN(new_n146));
  NAND2_X1  g024(.A1(new_n125), .A2(new_n131), .ZN(new_n147));
  NOR2_X1   g025(.A1(new_n140), .A2(G110), .ZN(new_n148));
  NOR2_X1   g026(.A1(new_n135), .A2(new_n136), .ZN(new_n149));
  OAI211_X1 g027(.A(new_n133), .B(new_n147), .C1(new_n148), .C2(new_n149), .ZN(new_n150));
  AND3_X1   g028(.A1(new_n142), .A2(new_n146), .A3(new_n150), .ZN(new_n151));
  AOI21_X1  g029(.A(new_n146), .B1(new_n142), .B2(new_n150), .ZN(new_n152));
  OAI221_X1 g030(.A(new_n123), .B1(new_n124), .B2(G234), .C1(new_n151), .C2(new_n152), .ZN(new_n153));
  INV_X1    g031(.A(new_n153), .ZN(new_n154));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n155));
  NOR2_X1   g033(.A1(new_n151), .A2(new_n152), .ZN(new_n156));
  OAI21_X1  g034(.A(new_n155), .B1(new_n156), .B2(G902), .ZN(new_n157));
  OAI211_X1 g035(.A(KEYINPUT25), .B(new_n123), .C1(new_n151), .C2(new_n152), .ZN(new_n158));
  NAND2_X1  g036(.A1(new_n157), .A2(new_n158), .ZN(new_n159));
  AOI21_X1  g037(.A(new_n124), .B1(G234), .B2(new_n123), .ZN(new_n160));
  AOI21_X1  g038(.A(new_n154), .B1(new_n159), .B2(new_n160), .ZN(new_n161));
  INV_X1    g039(.A(new_n161), .ZN(new_n162));
  NAND2_X1  g040(.A1(new_n131), .A2(G143), .ZN(new_n163));
  INV_X1    g041(.A(G143), .ZN(new_n164));
  NAND2_X1  g042(.A1(new_n164), .A2(G146), .ZN(new_n165));
  NAND2_X1  g043(.A1(new_n163), .A2(new_n165), .ZN(new_n166));
  OR2_X1    g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n167));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n168));
  NAND3_X1  g046(.A1(new_n166), .A2(new_n167), .A3(new_n168), .ZN(new_n169));
  NAND4_X1  g047(.A1(new_n163), .A2(new_n165), .A3(KEYINPUT0), .A4(G128), .ZN(new_n170));
  INV_X1    g048(.A(G131), .ZN(new_n171));
  INV_X1    g049(.A(G137), .ZN(new_n172));
  NAND3_X1  g050(.A1(new_n172), .A2(KEYINPUT11), .A3(G134), .ZN(new_n173));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n174));
  INV_X1    g052(.A(G134), .ZN(new_n175));
  AOI21_X1  g053(.A(new_n174), .B1(new_n175), .B2(G137), .ZN(new_n176));
  NOR2_X1   g054(.A1(new_n175), .A2(G137), .ZN(new_n177));
  OAI211_X1 g055(.A(new_n171), .B(new_n173), .C1(new_n176), .C2(new_n177), .ZN(new_n178));
  INV_X1    g056(.A(new_n178), .ZN(new_n179));
  OAI21_X1  g057(.A(KEYINPUT11), .B1(new_n172), .B2(G134), .ZN(new_n180));
  NAND2_X1  g058(.A1(new_n172), .A2(G134), .ZN(new_n181));
  NAND2_X1  g059(.A1(new_n180), .A2(new_n181), .ZN(new_n182));
  AOI21_X1  g060(.A(new_n171), .B1(new_n182), .B2(new_n173), .ZN(new_n183));
  OAI211_X1 g061(.A(new_n169), .B(new_n170), .C1(new_n179), .C2(new_n183), .ZN(new_n184));
  NOR2_X1   g062(.A1(new_n172), .A2(G134), .ZN(new_n185));
  OAI21_X1  g063(.A(G131), .B1(new_n177), .B2(new_n185), .ZN(new_n186));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n187));
  AND4_X1   g065(.A1(new_n187), .A2(new_n163), .A3(new_n165), .A4(G128), .ZN(new_n188));
  OAI21_X1  g066(.A(KEYINPUT1), .B1(new_n164), .B2(G146), .ZN(new_n189));
  AOI22_X1  g067(.A1(new_n189), .A2(G128), .B1(new_n163), .B2(new_n165), .ZN(new_n190));
  OAI211_X1 g068(.A(new_n178), .B(new_n186), .C1(new_n188), .C2(new_n190), .ZN(new_n191));
  NAND2_X1  g069(.A1(new_n184), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g070(.A(G116), .B(G119), .ZN(new_n193));
  XNOR2_X1  g071(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  XOR2_X1   g072(.A(new_n193), .B(new_n194), .Z(new_n195));
  NAND2_X1  g073(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g074(.A(new_n193), .B(new_n194), .ZN(new_n197));
  NAND3_X1  g075(.A1(new_n184), .A2(new_n197), .A3(new_n191), .ZN(new_n198));
  AND2_X1   g076(.A1(new_n198), .A2(KEYINPUT28), .ZN(new_n199));
  NOR2_X1   g077(.A1(new_n198), .A2(KEYINPUT28), .ZN(new_n200));
  OAI21_X1  g078(.A(new_n196), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n202));
  NAND2_X1  g080(.A1(new_n202), .A2(G210), .ZN(new_n203));
  XNOR2_X1  g081(.A(new_n203), .B(KEYINPUT27), .ZN(new_n204));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n205));
  XNOR2_X1  g083(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g084(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g085(.A1(new_n201), .A2(new_n207), .ZN(new_n208));
  INV_X1    g086(.A(new_n198), .ZN(new_n209));
  NAND2_X1  g087(.A1(new_n169), .A2(new_n170), .ZN(new_n210));
  NAND2_X1  g088(.A1(new_n182), .A2(new_n173), .ZN(new_n211));
  NAND2_X1  g089(.A1(new_n211), .A2(G131), .ZN(new_n212));
  AOI21_X1  g090(.A(new_n210), .B1(new_n212), .B2(new_n178), .ZN(new_n213));
  NOR2_X1   g091(.A1(new_n188), .A2(new_n190), .ZN(new_n214));
  NAND2_X1  g092(.A1(new_n178), .A2(new_n186), .ZN(new_n215));
  NOR2_X1   g093(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g094(.A(KEYINPUT30), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n218));
  NAND3_X1  g096(.A1(new_n184), .A2(new_n218), .A3(new_n191), .ZN(new_n219));
  NAND2_X1  g097(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g098(.A(new_n209), .B1(new_n220), .B2(new_n195), .ZN(new_n221));
  AOI21_X1  g099(.A(KEYINPUT31), .B1(new_n221), .B2(new_n206), .ZN(new_n222));
  AOI21_X1  g100(.A(new_n197), .B1(new_n217), .B2(new_n219), .ZN(new_n223));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n224));
  NOR4_X1   g102(.A1(new_n223), .A2(new_n224), .A3(new_n209), .A4(new_n207), .ZN(new_n225));
  OAI21_X1  g103(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g104(.A(G472), .ZN(new_n227));
  NAND3_X1  g105(.A1(new_n226), .A2(new_n227), .A3(new_n123), .ZN(new_n228));
  NAND2_X1  g106(.A1(new_n228), .A2(KEYINPUT32), .ZN(new_n229));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n230));
  NAND4_X1  g108(.A1(new_n226), .A2(new_n230), .A3(new_n227), .A4(new_n123), .ZN(new_n231));
  NAND2_X1  g109(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g110(.A(KEYINPUT29), .B1(new_n201), .B2(new_n207), .ZN(new_n233));
  OAI21_X1  g111(.A(new_n207), .B1(new_n223), .B2(new_n209), .ZN(new_n234));
  XNOR2_X1  g112(.A(new_n198), .B(KEYINPUT28), .ZN(new_n235));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n236));
  NAND4_X1  g114(.A1(new_n235), .A2(new_n236), .A3(new_n206), .A4(new_n196), .ZN(new_n237));
  NAND3_X1  g115(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g116(.A(new_n227), .B1(new_n238), .B2(new_n123), .ZN(new_n239));
  INV_X1    g117(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g118(.A(new_n162), .B1(new_n232), .B2(new_n240), .ZN(new_n241));
  INV_X1    g119(.A(G469), .ZN(new_n242));
  INV_X1    g120(.A(G101), .ZN(new_n243));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n244));
  INV_X1    g122(.A(G107), .ZN(new_n245));
  NAND3_X1  g123(.A1(new_n244), .A2(new_n245), .A3(G104), .ZN(new_n246));
  INV_X1    g124(.A(G104), .ZN(new_n247));
  AOI21_X1  g125(.A(KEYINPUT3), .B1(new_n247), .B2(G107), .ZN(new_n248));
  NOR2_X1   g126(.A1(new_n247), .A2(G107), .ZN(new_n249));
  OAI211_X1 g127(.A(new_n243), .B(new_n246), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NOR2_X1   g128(.A1(new_n245), .A2(G104), .ZN(new_n251));
  OAI21_X1  g129(.A(G101), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g130(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g131(.A1(new_n214), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g132(.A(new_n250), .B(new_n252), .C1(new_n188), .C2(new_n190), .ZN(new_n255));
  NAND2_X1  g133(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g134(.A1(new_n179), .A2(new_n183), .ZN(new_n257));
  INV_X1    g135(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g136(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g137(.A1(new_n259), .A2(KEYINPUT12), .ZN(new_n260));
  OAI21_X1  g138(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n261));
  NAND2_X1  g139(.A1(new_n261), .A2(G101), .ZN(new_n262));
  NAND3_X1  g140(.A1(new_n262), .A2(KEYINPUT4), .A3(new_n250), .ZN(new_n263));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g142(.A1(new_n261), .A2(new_n264), .A3(G101), .ZN(new_n265));
  NAND4_X1  g143(.A1(new_n263), .A2(new_n169), .A3(new_n170), .A4(new_n265), .ZN(new_n266));
  AND2_X1   g144(.A1(new_n255), .A2(KEYINPUT10), .ZN(new_n267));
  NOR2_X1   g145(.A1(new_n255), .A2(KEYINPUT10), .ZN(new_n268));
  OAI211_X1 g146(.A(new_n266), .B(new_n257), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g147(.A(KEYINPUT12), .ZN(new_n270));
  NAND3_X1  g148(.A1(new_n256), .A2(new_n270), .A3(new_n258), .ZN(new_n271));
  NAND3_X1  g149(.A1(new_n260), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g150(.A(G110), .B(G140), .ZN(new_n273));
  AND2_X1   g151(.A1(new_n144), .A2(G227), .ZN(new_n274));
  XOR2_X1   g152(.A(new_n273), .B(new_n274), .Z(new_n275));
  INV_X1    g153(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g154(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g155(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n278));
  NAND2_X1  g156(.A1(new_n278), .A2(new_n258), .ZN(new_n279));
  AOI21_X1  g157(.A(new_n275), .B1(new_n279), .B2(new_n269), .ZN(new_n280));
  OAI211_X1 g158(.A(new_n242), .B(new_n123), .C1(new_n277), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g159(.A1(new_n272), .A2(new_n276), .ZN(new_n282));
  NAND3_X1  g160(.A1(new_n279), .A2(new_n269), .A3(new_n275), .ZN(new_n283));
  AOI21_X1  g161(.A(G902), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g162(.A(new_n281), .B1(new_n242), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g163(.A(KEYINPUT9), .B(G234), .ZN(new_n286));
  OAI21_X1  g164(.A(G221), .B1(new_n286), .B2(G902), .ZN(new_n287));
  NAND2_X1  g165(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g166(.A(new_n288), .ZN(new_n289));
  INV_X1    g167(.A(G475), .ZN(new_n290));
  INV_X1    g168(.A(G237), .ZN(new_n291));
  NAND3_X1  g169(.A1(new_n291), .A2(new_n144), .A3(G214), .ZN(new_n292));
  NAND2_X1  g170(.A1(new_n292), .A2(new_n164), .ZN(new_n293));
  NAND3_X1  g171(.A1(new_n202), .A2(G143), .A3(G214), .ZN(new_n294));
  NAND2_X1  g172(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g173(.A1(new_n295), .A2(G131), .ZN(new_n296));
  INV_X1    g174(.A(KEYINPUT17), .ZN(new_n297));
  NAND3_X1  g175(.A1(new_n293), .A2(new_n171), .A3(new_n294), .ZN(new_n298));
  NAND3_X1  g176(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g177(.A1(new_n295), .A2(KEYINPUT17), .A3(G131), .ZN(new_n300));
  NAND4_X1  g178(.A1(new_n299), .A2(new_n132), .A3(new_n300), .A4(new_n133), .ZN(new_n301));
  XNOR2_X1  g179(.A(G113), .B(G122), .ZN(new_n302));
  XNOR2_X1  g180(.A(new_n302), .B(new_n247), .ZN(new_n303));
  NAND3_X1  g181(.A1(new_n295), .A2(KEYINPUT18), .A3(G131), .ZN(new_n304));
  XNOR2_X1  g182(.A(new_n125), .B(new_n131), .ZN(new_n305));
  NAND2_X1  g183(.A1(KEYINPUT18), .A2(G131), .ZN(new_n306));
  NAND3_X1  g184(.A1(new_n293), .A2(new_n294), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g185(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g186(.A1(new_n301), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  INV_X1    g187(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g188(.A1(new_n296), .A2(new_n298), .ZN(new_n311));
  AND2_X1   g189(.A1(new_n125), .A2(KEYINPUT19), .ZN(new_n312));
  NOR2_X1   g190(.A1(new_n125), .A2(KEYINPUT19), .ZN(new_n313));
  NOR2_X1   g191(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g192(.A(new_n311), .B(new_n133), .C1(G146), .C2(new_n314), .ZN(new_n315));
  AOI21_X1  g193(.A(new_n303), .B1(new_n315), .B2(new_n308), .ZN(new_n316));
  OAI211_X1 g194(.A(new_n290), .B(new_n123), .C1(new_n310), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g195(.A1(new_n317), .A2(KEYINPUT20), .ZN(new_n318));
  NAND2_X1  g196(.A1(new_n315), .A2(new_n308), .ZN(new_n319));
  INV_X1    g197(.A(new_n303), .ZN(new_n320));
  NAND2_X1  g198(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g199(.A(G475), .B1(new_n321), .B2(new_n309), .ZN(new_n322));
  INV_X1    g200(.A(KEYINPUT20), .ZN(new_n323));
  NAND3_X1  g201(.A1(new_n322), .A2(new_n323), .A3(new_n123), .ZN(new_n324));
  NAND2_X1  g202(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g203(.A(new_n303), .B1(new_n301), .B2(new_n308), .ZN(new_n326));
  OAI21_X1  g204(.A(new_n123), .B1(new_n310), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g205(.A1(new_n327), .A2(G475), .ZN(new_n328));
  AND2_X1   g206(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g207(.A(G116), .B(G122), .Z(new_n330));
  NAND2_X1  g208(.A1(new_n330), .A2(G107), .ZN(new_n331));
  XNOR2_X1  g209(.A(G116), .B(G122), .ZN(new_n332));
  NAND2_X1  g210(.A1(new_n332), .A2(new_n245), .ZN(new_n333));
  NAND2_X1  g211(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g212(.A1(new_n164), .A2(G128), .ZN(new_n335));
  INV_X1    g213(.A(G128), .ZN(new_n336));
  NAND2_X1  g214(.A1(new_n336), .A2(G143), .ZN(new_n337));
  NAND3_X1  g215(.A1(new_n335), .A2(new_n337), .A3(new_n175), .ZN(new_n338));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n339));
  OAI21_X1  g217(.A(new_n337), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g218(.A(KEYINPUT13), .B1(new_n164), .B2(G128), .ZN(new_n341));
  OAI21_X1  g219(.A(G134), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g220(.A1(new_n334), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  INV_X1    g221(.A(G116), .ZN(new_n344));
  NAND3_X1  g222(.A1(new_n344), .A2(KEYINPUT14), .A3(G122), .ZN(new_n345));
  OAI211_X1 g223(.A(G107), .B(new_n345), .C1(new_n330), .C2(KEYINPUT14), .ZN(new_n346));
  NAND2_X1  g224(.A1(new_n335), .A2(new_n337), .ZN(new_n347));
  NAND2_X1  g225(.A1(new_n347), .A2(G134), .ZN(new_n348));
  NAND2_X1  g226(.A1(new_n348), .A2(new_n338), .ZN(new_n349));
  NAND3_X1  g227(.A1(new_n346), .A2(new_n349), .A3(new_n333), .ZN(new_n350));
  NOR3_X1   g228(.A1(new_n286), .A2(new_n124), .A3(G953), .ZN(new_n351));
  AND3_X1   g229(.A1(new_n343), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g230(.A(new_n351), .B1(new_n343), .B2(new_n350), .ZN(new_n353));
  NOR2_X1   g231(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g232(.A1(new_n354), .A2(G902), .ZN(new_n355));
  INV_X1    g233(.A(G478), .ZN(new_n356));
  OR3_X1    g234(.A1(new_n355), .A2(KEYINPUT15), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g235(.A(new_n355), .B1(KEYINPUT15), .B2(new_n356), .ZN(new_n358));
  NAND2_X1  g236(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g237(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g238(.A1(new_n329), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g239(.A(G214), .B1(G237), .B2(G902), .ZN(new_n362));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n363));
  XNOR2_X1  g241(.A(new_n363), .B(KEYINPUT8), .ZN(new_n364));
  INV_X1    g242(.A(new_n253), .ZN(new_n365));
  INV_X1    g243(.A(new_n194), .ZN(new_n366));
  NAND2_X1  g244(.A1(new_n366), .A2(new_n193), .ZN(new_n367));
  NAND3_X1  g245(.A1(new_n138), .A2(KEYINPUT5), .A3(G116), .ZN(new_n368));
  OAI21_X1  g246(.A(new_n368), .B1(G116), .B2(new_n138), .ZN(new_n369));
  AOI21_X1  g247(.A(KEYINPUT5), .B1(new_n138), .B2(G116), .ZN(new_n370));
  OAI21_X1  g248(.A(G113), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND3_X1   g249(.A1(new_n365), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  AOI22_X1  g250(.A1(new_n371), .A2(new_n367), .B1(new_n250), .B2(new_n252), .ZN(new_n373));
  OAI21_X1  g251(.A(new_n364), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g252(.A1(new_n195), .A2(new_n263), .A3(new_n265), .ZN(new_n375));
  NAND3_X1  g253(.A1(new_n365), .A2(new_n367), .A3(new_n371), .ZN(new_n376));
  NAND3_X1  g254(.A1(new_n375), .A2(new_n376), .A3(new_n363), .ZN(new_n377));
  INV_X1    g255(.A(G125), .ZN(new_n378));
  OAI21_X1  g256(.A(new_n378), .B1(new_n188), .B2(new_n190), .ZN(new_n379));
  NAND3_X1  g257(.A1(new_n169), .A2(G125), .A3(new_n170), .ZN(new_n380));
  NAND2_X1  g258(.A1(new_n144), .A2(G224), .ZN(new_n381));
  NAND2_X1  g259(.A1(new_n381), .A2(KEYINPUT7), .ZN(new_n382));
  NAND3_X1  g260(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g261(.A1(new_n379), .A2(new_n380), .ZN(new_n384));
  NAND3_X1  g262(.A1(new_n384), .A2(KEYINPUT7), .A3(new_n381), .ZN(new_n385));
  NAND4_X1  g263(.A1(new_n374), .A2(new_n377), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  AND2_X1   g264(.A1(new_n386), .A2(new_n123), .ZN(new_n387));
  NAND2_X1  g265(.A1(new_n375), .A2(new_n376), .ZN(new_n388));
  INV_X1    g266(.A(new_n363), .ZN(new_n389));
  NAND2_X1  g267(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g268(.A1(new_n390), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n391));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n392));
  NAND3_X1  g270(.A1(new_n388), .A2(new_n392), .A3(new_n389), .ZN(new_n393));
  XNOR2_X1  g271(.A(new_n384), .B(new_n381), .ZN(new_n394));
  NAND3_X1  g272(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n396));
  AND3_X1   g274(.A1(new_n387), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g275(.A(new_n396), .B1(new_n387), .B2(new_n395), .ZN(new_n398));
  OAI21_X1  g276(.A(new_n362), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g277(.A(G952), .ZN(new_n400));
  AOI211_X1 g278(.A(G953), .B(new_n400), .C1(G234), .C2(G237), .ZN(new_n401));
  XOR2_X1   g279(.A(KEYINPUT21), .B(G898), .Z(new_n402));
  NOR2_X1   g280(.A1(new_n402), .A2(new_n144), .ZN(new_n403));
  AOI21_X1  g281(.A(new_n123), .B1(G234), .B2(G237), .ZN(new_n404));
  AOI21_X1  g282(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR3_X1   g283(.A1(new_n361), .A2(new_n399), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g284(.A1(new_n241), .A2(new_n289), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g285(.A(new_n407), .B(G101), .ZN(G3));
  AOI21_X1  g286(.A(new_n206), .B1(new_n235), .B2(new_n196), .ZN(new_n409));
  AND3_X1   g287(.A1(new_n184), .A2(new_n218), .A3(new_n191), .ZN(new_n410));
  AOI21_X1  g288(.A(new_n218), .B1(new_n184), .B2(new_n191), .ZN(new_n411));
  OAI21_X1  g289(.A(new_n195), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g290(.A1(new_n412), .A2(new_n206), .A3(new_n198), .ZN(new_n413));
  NAND2_X1  g291(.A1(new_n413), .A2(new_n224), .ZN(new_n414));
  NAND3_X1  g292(.A1(new_n221), .A2(KEYINPUT31), .A3(new_n206), .ZN(new_n415));
  AOI21_X1  g293(.A(new_n409), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g294(.A(G472), .B1(new_n416), .B2(G902), .ZN(new_n417));
  NAND3_X1  g295(.A1(new_n417), .A2(new_n228), .A3(new_n161), .ZN(new_n418));
  NOR3_X1   g296(.A1(new_n418), .A2(new_n288), .A3(new_n399), .ZN(new_n419));
  OR3_X1    g297(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT33), .ZN(new_n420));
  OAI21_X1  g298(.A(KEYINPUT33), .B1(new_n352), .B2(new_n353), .ZN(new_n421));
  NAND2_X1  g299(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g300(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g301(.A(G478), .B1(new_n423), .B2(G902), .ZN(new_n424));
  NAND2_X1  g302(.A1(new_n355), .A2(new_n356), .ZN(new_n425));
  NAND2_X1  g303(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g304(.A1(new_n329), .A2(new_n426), .A3(new_n405), .ZN(new_n427));
  NAND2_X1  g305(.A1(new_n419), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g306(.A(KEYINPUT34), .B(G104), .Z(new_n429));
  XNOR2_X1  g307(.A(new_n428), .B(new_n429), .ZN(G6));
  NAND2_X1  g308(.A1(new_n329), .A2(new_n359), .ZN(new_n431));
  NOR2_X1   g309(.A1(new_n431), .A2(new_n405), .ZN(new_n432));
  NAND2_X1  g310(.A1(new_n419), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G107), .Z(new_n434));
  XNOR2_X1  g312(.A(new_n433), .B(new_n434), .ZN(G9));
  NAND2_X1  g313(.A1(new_n417), .A2(new_n228), .ZN(new_n436));
  NAND2_X1  g314(.A1(new_n159), .A2(new_n160), .ZN(new_n437));
  NAND2_X1  g315(.A1(new_n142), .A2(new_n150), .ZN(new_n438));
  NOR2_X1   g316(.A1(new_n146), .A2(KEYINPUT36), .ZN(new_n439));
  XNOR2_X1  g317(.A(new_n438), .B(new_n439), .ZN(new_n440));
  OAI211_X1 g318(.A(new_n440), .B(new_n123), .C1(new_n124), .C2(G234), .ZN(new_n441));
  NAND2_X1  g319(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g320(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g321(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g322(.A1(new_n406), .A2(new_n444), .A3(new_n289), .ZN(new_n445));
  XOR2_X1   g323(.A(KEYINPUT37), .B(G110), .Z(new_n446));
  XNOR2_X1  g324(.A(new_n445), .B(new_n446), .ZN(G12));
  AOI21_X1  g325(.A(new_n443), .B1(new_n232), .B2(new_n240), .ZN(new_n448));
  INV_X1    g326(.A(new_n399), .ZN(new_n449));
  NOR2_X1   g327(.A1(new_n144), .A2(G900), .ZN(new_n450));
  AND2_X1   g328(.A1(new_n404), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g329(.A(new_n329), .B(new_n359), .C1(new_n401), .C2(new_n451), .ZN(new_n452));
  INV_X1    g330(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g331(.A1(new_n448), .A2(new_n289), .A3(new_n449), .A4(new_n453), .ZN(new_n454));
  XNOR2_X1  g332(.A(new_n454), .B(G128), .ZN(G30));
  INV_X1    g333(.A(new_n362), .ZN(new_n456));
  NOR2_X1   g334(.A1(new_n451), .A2(new_n401), .ZN(new_n457));
  XOR2_X1   g335(.A(new_n457), .B(KEYINPUT39), .Z(new_n458));
  NAND2_X1  g336(.A1(new_n289), .A2(new_n458), .ZN(new_n459));
  INV_X1    g337(.A(KEYINPUT40), .ZN(new_n460));
  NAND2_X1  g338(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g339(.A1(new_n289), .A2(KEYINPUT40), .A3(new_n458), .ZN(new_n462));
  AOI21_X1  g340(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g341(.A1(new_n397), .A2(new_n398), .ZN(new_n464));
  XOR2_X1   g342(.A(new_n464), .B(KEYINPUT38), .Z(new_n465));
  AOI21_X1  g343(.A(new_n206), .B1(new_n196), .B2(new_n198), .ZN(new_n466));
  AOI21_X1  g344(.A(new_n466), .B1(new_n221), .B2(new_n206), .ZN(new_n467));
  OAI21_X1  g345(.A(G472), .B1(new_n467), .B2(G902), .ZN(new_n468));
  NAND2_X1  g346(.A1(new_n232), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g347(.A1(new_n325), .A2(new_n328), .ZN(new_n470));
  NAND2_X1  g348(.A1(new_n470), .A2(new_n359), .ZN(new_n471));
  INV_X1    g349(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g350(.A1(new_n463), .A2(new_n465), .A3(new_n469), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g351(.A1(new_n473), .A2(new_n442), .ZN(new_n474));
  XNOR2_X1  g352(.A(new_n474), .B(new_n164), .ZN(G45));
  NOR3_X1   g353(.A1(new_n329), .A2(new_n426), .A3(new_n457), .ZN(new_n476));
  NAND4_X1  g354(.A1(new_n448), .A2(new_n289), .A3(new_n449), .A4(new_n476), .ZN(new_n477));
  XNOR2_X1  g355(.A(new_n477), .B(G146), .ZN(G48));
  NAND2_X1  g356(.A1(new_n414), .A2(new_n415), .ZN(new_n479));
  AOI21_X1  g357(.A(G902), .B1(new_n479), .B2(new_n208), .ZN(new_n480));
  AOI21_X1  g358(.A(new_n230), .B1(new_n480), .B2(new_n227), .ZN(new_n481));
  INV_X1    g359(.A(new_n231), .ZN(new_n482));
  OAI21_X1  g360(.A(new_n240), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g361(.A(new_n123), .B1(new_n277), .B2(new_n280), .ZN(new_n484));
  NAND2_X1  g362(.A1(new_n484), .A2(G469), .ZN(new_n485));
  NAND3_X1  g363(.A1(new_n485), .A2(new_n287), .A3(new_n281), .ZN(new_n486));
  NOR2_X1   g364(.A1(new_n486), .A2(new_n399), .ZN(new_n487));
  NAND4_X1  g365(.A1(new_n483), .A2(new_n161), .A3(new_n427), .A4(new_n487), .ZN(new_n488));
  XNOR2_X1  g366(.A(KEYINPUT41), .B(G113), .ZN(new_n489));
  XNOR2_X1  g367(.A(new_n488), .B(new_n489), .ZN(G15));
  NAND4_X1  g368(.A1(new_n483), .A2(new_n161), .A3(new_n432), .A4(new_n487), .ZN(new_n491));
  XNOR2_X1  g369(.A(new_n491), .B(G116), .ZN(G18));
  NOR2_X1   g370(.A1(new_n361), .A2(new_n405), .ZN(new_n493));
  INV_X1    g371(.A(new_n486), .ZN(new_n494));
  NAND4_X1  g372(.A1(new_n448), .A2(new_n449), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  XNOR2_X1  g373(.A(new_n495), .B(G119), .ZN(G21));
  NOR2_X1   g374(.A1(new_n418), .A2(new_n405), .ZN(new_n497));
  NOR3_X1   g375(.A1(new_n471), .A2(new_n486), .A3(new_n399), .ZN(new_n498));
  NAND2_X1  g376(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g377(.A(new_n499), .B(G122), .ZN(G24));
  NAND3_X1  g378(.A1(new_n444), .A2(new_n476), .A3(new_n487), .ZN(new_n501));
  XNOR2_X1  g379(.A(new_n501), .B(G125), .ZN(G27));
  NAND4_X1  g380(.A1(new_n464), .A2(new_n285), .A3(new_n287), .A4(new_n362), .ZN(new_n503));
  INV_X1    g381(.A(new_n503), .ZN(new_n504));
  NAND4_X1  g382(.A1(new_n483), .A2(new_n161), .A3(new_n476), .A4(new_n504), .ZN(new_n505));
  INV_X1    g383(.A(KEYINPUT42), .ZN(new_n506));
  NAND2_X1  g384(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g385(.A1(new_n241), .A2(KEYINPUT42), .A3(new_n476), .A4(new_n504), .ZN(new_n508));
  NAND2_X1  g386(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g387(.A(new_n509), .B(G131), .ZN(G33));
  AOI21_X1  g388(.A(new_n239), .B1(new_n229), .B2(new_n231), .ZN(new_n511));
  NOR4_X1   g389(.A1(new_n511), .A2(new_n452), .A3(new_n503), .A4(new_n162), .ZN(new_n512));
  XNOR2_X1  g390(.A(new_n512), .B(new_n175), .ZN(G36));
  INV_X1    g391(.A(new_n426), .ZN(new_n514));
  NAND2_X1  g392(.A1(new_n514), .A2(new_n329), .ZN(new_n515));
  NAND2_X1  g393(.A1(new_n515), .A2(KEYINPUT43), .ZN(new_n516));
  OR3_X1    g394(.A1(new_n426), .A2(new_n470), .A3(KEYINPUT43), .ZN(new_n517));
  AND2_X1   g395(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g396(.A1(new_n518), .A2(new_n436), .A3(new_n442), .ZN(new_n519));
  INV_X1    g397(.A(KEYINPUT44), .ZN(new_n520));
  OR2_X1    g398(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g399(.A1(new_n464), .A2(new_n362), .ZN(new_n522));
  INV_X1    g400(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g401(.A1(new_n519), .A2(new_n520), .ZN(new_n524));
  NAND2_X1  g402(.A1(new_n282), .A2(new_n283), .ZN(new_n525));
  XNOR2_X1  g403(.A(new_n525), .B(KEYINPUT45), .ZN(new_n526));
  OAI21_X1  g404(.A(G469), .B1(new_n526), .B2(G902), .ZN(new_n527));
  NAND2_X1  g405(.A1(new_n527), .A2(KEYINPUT46), .ZN(new_n528));
  INV_X1    g406(.A(KEYINPUT46), .ZN(new_n529));
  OAI211_X1 g407(.A(new_n529), .B(G469), .C1(new_n526), .C2(G902), .ZN(new_n530));
  NAND3_X1  g408(.A1(new_n528), .A2(new_n281), .A3(new_n530), .ZN(new_n531));
  AND3_X1   g409(.A1(new_n531), .A2(new_n287), .A3(new_n458), .ZN(new_n532));
  NAND4_X1  g410(.A1(new_n521), .A2(new_n523), .A3(new_n524), .A4(new_n532), .ZN(new_n533));
  XNOR2_X1  g411(.A(new_n533), .B(G137), .ZN(G39));
  NAND2_X1  g412(.A1(new_n531), .A2(new_n287), .ZN(new_n535));
  INV_X1    g413(.A(KEYINPUT47), .ZN(new_n536));
  NAND2_X1  g414(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g415(.A1(new_n531), .A2(KEYINPUT47), .A3(new_n287), .ZN(new_n538));
  AOI21_X1  g416(.A(new_n522), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g417(.A1(new_n539), .A2(new_n162), .A3(new_n511), .A4(new_n476), .ZN(new_n540));
  XNOR2_X1  g418(.A(new_n540), .B(G140), .ZN(G42));
  AND3_X1   g419(.A1(new_n516), .A2(new_n401), .A3(new_n517), .ZN(new_n542));
  INV_X1    g420(.A(new_n418), .ZN(new_n543));
  AND2_X1   g421(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g422(.A1(new_n465), .A2(new_n362), .ZN(new_n545));
  NAND3_X1  g423(.A1(new_n544), .A2(new_n494), .A3(new_n545), .ZN(new_n546));
  INV_X1    g424(.A(KEYINPUT50), .ZN(new_n547));
  NAND2_X1  g425(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g426(.A1(new_n544), .A2(KEYINPUT50), .A3(new_n494), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g427(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g428(.A1(new_n469), .A2(new_n162), .ZN(new_n551));
  NOR2_X1   g429(.A1(new_n514), .A2(new_n470), .ZN(new_n552));
  NAND3_X1  g430(.A1(new_n551), .A2(new_n401), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g431(.A1(new_n542), .A2(new_n444), .ZN(new_n554));
  AOI21_X1  g432(.A(new_n486), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g433(.A(new_n485), .ZN(new_n556));
  INV_X1    g434(.A(new_n281), .ZN(new_n557));
  NOR2_X1   g435(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g436(.A(new_n558), .ZN(new_n559));
  OAI211_X1 g437(.A(new_n537), .B(new_n538), .C1(new_n287), .C2(new_n559), .ZN(new_n560));
  AOI21_X1  g438(.A(new_n555), .B1(new_n560), .B2(new_n544), .ZN(new_n561));
  OAI21_X1  g439(.A(new_n550), .B1(new_n561), .B2(new_n522), .ZN(new_n562));
  INV_X1    g440(.A(KEYINPUT51), .ZN(new_n563));
  NAND2_X1  g441(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g442(.A(new_n550), .B(KEYINPUT51), .C1(new_n561), .C2(new_n522), .ZN(new_n565));
  NOR2_X1   g443(.A1(new_n522), .A2(new_n486), .ZN(new_n566));
  NAND3_X1  g444(.A1(new_n542), .A2(new_n241), .A3(new_n566), .ZN(new_n567));
  INV_X1    g445(.A(KEYINPUT48), .ZN(new_n568));
  AND2_X1   g446(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g447(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NOR2_X1   g448(.A1(new_n329), .A2(new_n426), .ZN(new_n571));
  AND4_X1   g449(.A1(new_n401), .A2(new_n551), .A3(new_n571), .A4(new_n566), .ZN(new_n572));
  NOR3_X1   g450(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g451(.A(new_n558), .B(KEYINPUT49), .Z(new_n574));
  NOR4_X1   g452(.A1(new_n574), .A2(new_n162), .A3(new_n456), .A4(new_n465), .ZN(new_n575));
  NAND2_X1  g453(.A1(new_n575), .A2(new_n287), .ZN(new_n576));
  OR3_X1    g454(.A1(new_n576), .A2(new_n469), .A3(new_n515), .ZN(new_n577));
  NAND4_X1  g455(.A1(new_n564), .A2(new_n565), .A3(new_n573), .A4(new_n577), .ZN(new_n578));
  INV_X1    g456(.A(KEYINPUT54), .ZN(new_n579));
  NOR2_X1   g457(.A1(new_n288), .A2(new_n457), .ZN(new_n580));
  NOR3_X1   g458(.A1(new_n471), .A2(new_n442), .A3(new_n399), .ZN(new_n581));
  NAND3_X1  g459(.A1(new_n469), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g460(.A1(new_n454), .A2(new_n477), .A3(new_n501), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g461(.A1(new_n583), .A2(KEYINPUT52), .ZN(new_n584));
  NOR3_X1   g462(.A1(new_n511), .A2(new_n399), .A3(new_n443), .ZN(new_n585));
  OAI211_X1 g463(.A(new_n585), .B(new_n289), .C1(new_n453), .C2(new_n476), .ZN(new_n586));
  INV_X1    g464(.A(KEYINPUT52), .ZN(new_n587));
  NAND4_X1  g465(.A1(new_n586), .A2(new_n587), .A3(new_n501), .A4(new_n582), .ZN(new_n588));
  AND2_X1   g466(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g467(.A1(new_n419), .A2(new_n432), .B1(new_n497), .B2(new_n498), .ZN(new_n590));
  NAND3_X1  g468(.A1(new_n495), .A2(new_n407), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g469(.A1(new_n488), .A2(new_n491), .A3(new_n428), .A4(new_n445), .ZN(new_n592));
  OR2_X1    g470(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g471(.A(new_n512), .ZN(new_n594));
  NAND3_X1  g472(.A1(new_n444), .A2(new_n504), .A3(new_n476), .ZN(new_n595));
  INV_X1    g473(.A(new_n361), .ZN(new_n596));
  NAND4_X1  g474(.A1(new_n448), .A2(new_n596), .A3(new_n523), .A4(new_n580), .ZN(new_n597));
  NAND4_X1  g475(.A1(new_n509), .A2(new_n594), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NOR2_X1   g476(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g477(.A(KEYINPUT53), .B1(new_n589), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g478(.A1(new_n591), .A2(new_n592), .ZN(new_n601));
  AOI21_X1  g479(.A(new_n512), .B1(new_n507), .B2(new_n508), .ZN(new_n602));
  NAND4_X1  g480(.A1(new_n601), .A2(new_n595), .A3(new_n602), .A4(new_n597), .ZN(new_n603));
  NAND2_X1  g481(.A1(new_n584), .A2(new_n588), .ZN(new_n604));
  INV_X1    g482(.A(KEYINPUT53), .ZN(new_n605));
  NOR3_X1   g483(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g484(.A(new_n579), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g485(.A1(new_n589), .A2(new_n599), .A3(KEYINPUT53), .ZN(new_n608));
  OAI21_X1  g486(.A(new_n605), .B1(new_n603), .B2(new_n604), .ZN(new_n609));
  NAND3_X1  g487(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT54), .ZN(new_n610));
  AOI21_X1  g488(.A(new_n578), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  AOI211_X1 g489(.A(new_n400), .B(G953), .C1(new_n544), .C2(new_n487), .ZN(new_n612));
  NOR2_X1   g490(.A1(G952), .A2(G953), .ZN(new_n613));
  AOI22_X1  g491(.A1(new_n611), .A2(new_n612), .B1(new_n577), .B2(new_n613), .ZN(G75));
  NAND2_X1  g492(.A1(new_n391), .A2(new_n393), .ZN(new_n615));
  XOR2_X1   g493(.A(new_n615), .B(new_n394), .Z(new_n616));
  XNOR2_X1  g494(.A(new_n616), .B(KEYINPUT55), .ZN(new_n617));
  AOI21_X1  g495(.A(new_n123), .B1(new_n608), .B2(new_n609), .ZN(new_n618));
  INV_X1    g496(.A(new_n396), .ZN(new_n619));
  AOI211_X1 g497(.A(KEYINPUT56), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g498(.A(new_n617), .ZN(new_n621));
  NAND2_X1  g499(.A1(new_n608), .A2(new_n609), .ZN(new_n622));
  NAND3_X1  g500(.A1(new_n622), .A2(G902), .A3(new_n619), .ZN(new_n623));
  INV_X1    g501(.A(KEYINPUT56), .ZN(new_n624));
  AOI21_X1  g502(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g503(.A1(new_n144), .A2(G952), .ZN(new_n626));
  NOR3_X1   g504(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(G51));
  NAND2_X1  g505(.A1(G469), .A2(G902), .ZN(new_n628));
  XOR2_X1   g506(.A(new_n628), .B(KEYINPUT57), .Z(new_n629));
  NAND3_X1  g507(.A1(new_n607), .A2(new_n610), .A3(new_n629), .ZN(new_n630));
  INV_X1    g508(.A(new_n277), .ZN(new_n631));
  INV_X1    g509(.A(new_n280), .ZN(new_n632));
  NAND2_X1  g510(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g511(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g512(.A1(new_n622), .A2(G469), .A3(G902), .A4(new_n526), .ZN(new_n635));
  AOI21_X1  g513(.A(new_n626), .B1(new_n634), .B2(new_n635), .ZN(G54));
  AND2_X1   g514(.A1(KEYINPUT58), .A2(G475), .ZN(new_n637));
  NAND2_X1  g515(.A1(new_n618), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g516(.A1(new_n638), .A2(new_n309), .A3(new_n321), .ZN(new_n639));
  INV_X1    g517(.A(new_n626), .ZN(new_n640));
  OAI211_X1 g518(.A(new_n618), .B(new_n637), .C1(new_n310), .C2(new_n316), .ZN(new_n641));
  AND3_X1   g519(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(G60));
  NAND2_X1  g520(.A1(G478), .A2(G902), .ZN(new_n643));
  XNOR2_X1  g521(.A(new_n643), .B(KEYINPUT59), .ZN(new_n644));
  NAND3_X1  g522(.A1(new_n607), .A2(new_n610), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g523(.A1(new_n645), .A2(new_n423), .ZN(new_n646));
  NAND4_X1  g524(.A1(new_n607), .A2(new_n422), .A3(new_n610), .A4(new_n644), .ZN(new_n647));
  AND3_X1   g525(.A1(new_n646), .A2(new_n640), .A3(new_n647), .ZN(G63));
  INV_X1    g526(.A(KEYINPUT61), .ZN(new_n649));
  NAND2_X1  g527(.A1(G217), .A2(G902), .ZN(new_n650));
  XOR2_X1   g528(.A(new_n650), .B(KEYINPUT60), .Z(new_n651));
  INV_X1    g529(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g530(.A(new_n652), .B1(new_n608), .B2(new_n609), .ZN(new_n653));
  NAND2_X1  g531(.A1(new_n653), .A2(new_n440), .ZN(new_n654));
  INV_X1    g532(.A(new_n654), .ZN(new_n655));
  INV_X1    g533(.A(new_n156), .ZN(new_n656));
  OAI21_X1  g534(.A(new_n640), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g535(.A(new_n649), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g536(.A1(new_n653), .A2(new_n656), .ZN(new_n659));
  NAND4_X1  g537(.A1(new_n659), .A2(new_n654), .A3(KEYINPUT61), .A4(new_n640), .ZN(new_n660));
  NAND2_X1  g538(.A1(new_n658), .A2(new_n660), .ZN(G66));
  NAND2_X1  g539(.A1(new_n402), .A2(G224), .ZN(new_n662));
  NAND2_X1  g540(.A1(new_n662), .A2(G953), .ZN(new_n663));
  OAI21_X1  g541(.A(new_n663), .B1(new_n601), .B2(G953), .ZN(new_n664));
  OAI21_X1  g542(.A(new_n615), .B1(G898), .B2(new_n144), .ZN(new_n665));
  XNOR2_X1  g543(.A(new_n664), .B(new_n665), .ZN(G69));
  AOI21_X1  g544(.A(new_n144), .B1(G227), .B2(G900), .ZN(new_n667));
  AND2_X1   g545(.A1(new_n540), .A2(new_n533), .ZN(new_n668));
  INV_X1    g546(.A(new_n459), .ZN(new_n669));
  OAI21_X1  g547(.A(new_n431), .B1(new_n329), .B2(new_n426), .ZN(new_n670));
  NAND4_X1  g548(.A1(new_n241), .A2(new_n669), .A3(new_n523), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g549(.A1(new_n586), .A2(new_n501), .ZN(new_n672));
  OAI21_X1  g550(.A(KEYINPUT62), .B1(new_n474), .B2(new_n672), .ZN(new_n673));
  INV_X1    g551(.A(new_n672), .ZN(new_n674));
  INV_X1    g552(.A(KEYINPUT62), .ZN(new_n675));
  OAI211_X1 g553(.A(new_n674), .B(new_n675), .C1(new_n442), .C2(new_n473), .ZN(new_n676));
  NAND4_X1  g554(.A1(new_n668), .A2(new_n671), .A3(new_n673), .A4(new_n676), .ZN(new_n677));
  AOI21_X1  g555(.A(new_n667), .B1(new_n677), .B2(new_n144), .ZN(new_n678));
  XNOR2_X1  g556(.A(new_n220), .B(new_n314), .ZN(new_n679));
  NOR2_X1   g557(.A1(new_n679), .A2(new_n450), .ZN(new_n680));
  NAND4_X1  g558(.A1(new_n532), .A2(new_n241), .A3(new_n449), .A4(new_n472), .ZN(new_n681));
  AND2_X1   g559(.A1(new_n681), .A2(new_n602), .ZN(new_n682));
  NAND4_X1  g560(.A1(new_n540), .A2(new_n682), .A3(new_n533), .A4(new_n674), .ZN(new_n683));
  NAND2_X1  g561(.A1(new_n683), .A2(new_n144), .ZN(new_n684));
  NAND2_X1  g562(.A1(new_n684), .A2(new_n680), .ZN(new_n685));
  OAI22_X1  g563(.A1(new_n678), .A2(new_n680), .B1(new_n667), .B2(new_n685), .ZN(G72));
  NAND2_X1  g564(.A1(G472), .A2(G902), .ZN(new_n687));
  XNOR2_X1  g565(.A(new_n687), .B(KEYINPUT63), .ZN(new_n688));
  INV_X1    g566(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g567(.A(new_n689), .B1(new_n683), .B2(new_n593), .ZN(new_n690));
  NAND3_X1  g568(.A1(new_n690), .A2(new_n207), .A3(new_n221), .ZN(new_n691));
  NAND2_X1  g569(.A1(new_n234), .A2(new_n413), .ZN(new_n692));
  NAND3_X1  g570(.A1(new_n622), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g571(.A1(new_n691), .A2(new_n693), .A3(new_n640), .ZN(new_n694));
  OAI21_X1  g572(.A(new_n689), .B1(new_n677), .B2(new_n593), .ZN(new_n695));
  NOR2_X1   g573(.A1(new_n221), .A2(new_n207), .ZN(new_n696));
  AOI21_X1  g574(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(G57));
endmodule


