//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n203), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR3_X1   g008(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT93), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT94), .ZN(new_n214));
  XOR2_X1   g013(.A(G57gat), .B(G64gat), .Z(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(KEYINPUT94), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G71gat), .B(G78gat), .Z(new_n219));
  OR2_X1    g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n206), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(KEYINPUT97), .Z(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n222), .ZN(new_n225));
  NAND2_X1  g024(.A1(G231gat), .A2(G233gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(G127gat), .B(G155gat), .Z(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT20), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n227), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT96), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n230), .A2(new_n232), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n224), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n235), .ZN(new_n237));
  INV_X1    g036(.A(new_n224), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n238), .A3(new_n233), .ZN(new_n239));
  XOR2_X1   g038(.A(G183gat), .B(G211gat), .Z(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n236), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n236), .B2(new_n239), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(G134gat), .B(G162gat), .Z(new_n245));
  XNOR2_X1  g044(.A(G190gat), .B(G218gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT99), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT14), .ZN(new_n248));
  INV_X1    g047(.A(G29gat), .ZN(new_n249));
  INV_X1    g048(.A(G36gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n251), .A2(new_n252), .B1(G29gat), .B2(G36gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT85), .ZN(new_n254));
  XNOR2_X1  g053(.A(G43gat), .B(G50gat), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n253), .A2(new_n254), .B1(KEYINPUT15), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n253), .B1(KEYINPUT15), .B2(new_n255), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n257), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT86), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT17), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n259), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT86), .B1(new_n264), .B2(KEYINPUT17), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n260), .A2(new_n262), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269));
  INV_X1    g068(.A(G85gat), .ZN(new_n270));
  INV_X1    g069(.A(G92gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(KEYINPUT8), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT7), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n270), .B2(new_n271), .ZN(new_n274));
  NAND3_X1  g073(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G99gat), .B(G106gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT98), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OR3_X1    g079(.A1(new_n276), .A2(new_n279), .A3(new_n277), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n277), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n266), .A2(new_n268), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT41), .ZN(new_n285));
  NAND2_X1  g084(.A1(G232gat), .A2(G233gat), .ZN(new_n286));
  OAI22_X1  g085(.A1(new_n283), .A2(new_n264), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n247), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n267), .B1(new_n265), .B2(new_n263), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n289), .B2(new_n283), .ZN(new_n290));
  INV_X1    g089(.A(new_n247), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n285), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n288), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n288), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n245), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n288), .A2(new_n292), .ZN(new_n297));
  INV_X1    g096(.A(new_n293), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n288), .A2(new_n292), .A3(new_n293), .ZN(new_n300));
  INV_X1    g099(.A(new_n245), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n244), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G176gat), .B(G204gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n221), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n282), .A2(KEYINPUT100), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n311), .A2(new_n278), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n278), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n218), .B(new_n220), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT10), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n283), .A2(new_n221), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G230gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n310), .A2(new_n314), .A3(new_n320), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n308), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT103), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(KEYINPUT103), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n314), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n316), .ZN(new_n328));
  INV_X1    g127(.A(new_n317), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n319), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n322), .B(KEYINPUT101), .ZN(new_n332));
  INV_X1    g131(.A(new_n308), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT102), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n334), .A2(new_n335), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n325), .B(new_n326), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n266), .A2(new_n206), .A3(new_n268), .ZN(new_n340));
  NAND2_X1  g139(.A1(G229gat), .A2(G233gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n264), .A2(new_n206), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n340), .A2(KEYINPUT18), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(KEYINPUT88), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT88), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n264), .A2(new_n206), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n264), .A2(KEYINPUT89), .A3(new_n206), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT89), .B1(new_n264), .B2(new_n206), .ZN(new_n349));
  OAI22_X1  g148(.A1(new_n345), .A2(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT87), .B(KEYINPUT13), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(new_n341), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n344), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G113gat), .B(G141gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT11), .ZN(new_n357));
  INV_X1    g156(.A(G169gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G197gat), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NOR2_X1   g161(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n342), .B1(new_n289), .B2(new_n206), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n341), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT18), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n365), .A2(KEYINPUT91), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT91), .B1(new_n365), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n363), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n355), .A2(KEYINPUT90), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n344), .A2(new_n354), .A3(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n370), .A2(new_n372), .B1(new_n366), .B2(new_n365), .ZN(new_n373));
  INV_X1    g172(.A(new_n362), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n339), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n377));
  OR2_X1    g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(KEYINPUT76), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n381));
  AND2_X1   g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT2), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n386), .B2(new_n389), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n378), .A2(new_n379), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT77), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394));
  INV_X1    g193(.A(G155gat), .ZN(new_n395));
  INV_X1    g194(.A(G162gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(new_n397), .B2(KEYINPUT2), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT77), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n382), .A2(new_n383), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n387), .A2(new_n390), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G197gat), .B(G204gat), .ZN(new_n403));
  INV_X1    g202(.A(G211gat), .ZN(new_n404));
  INV_X1    g203(.A(G218gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(KEYINPUT22), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G211gat), .B(G218gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n402), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT2), .B1(new_n380), .B2(new_n384), .ZN(new_n416));
  INV_X1    g215(.A(new_n390), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n399), .B1(new_n398), .B2(new_n400), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT77), .ZN(new_n419));
  OAI221_X1 g218(.A(new_n413), .B1(new_n416), .B2(new_n417), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n410), .B1(new_n420), .B2(new_n411), .ZN(new_n421));
  OR3_X1    g220(.A1(new_n414), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n415), .B1(new_n414), .B2(new_n421), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(G22gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT31), .B(G50gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  MUX2_X1   g227(.A(G22gat), .B(new_n425), .S(new_n428), .Z(new_n429));
  AND3_X1   g228(.A1(new_n422), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n422), .B2(new_n423), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  XOR2_X1   g232(.A(G127gat), .B(G134gat), .Z(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT1), .ZN(new_n435));
  INV_X1    g234(.A(G120gat), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n436), .A2(G113gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(KEYINPUT67), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G120gat), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n440), .A3(G113gat), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n437), .B1(new_n441), .B2(KEYINPUT68), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT68), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT67), .B(G120gat), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(G113gat), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n435), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G113gat), .B(G120gat), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n447), .A2(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n434), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  OAI22_X1  g249(.A1(new_n419), .A2(new_n418), .B1(new_n416), .B2(new_n417), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n441), .A2(KEYINPUT68), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n444), .A2(new_n443), .A3(G113gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n437), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n455), .A2(new_n435), .B1(new_n448), .B2(new_n434), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n402), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n433), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n451), .A2(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n420), .A3(new_n450), .ZN(new_n463));
  XOR2_X1   g262(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n450), .B2(new_n451), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n456), .A2(new_n402), .A3(KEYINPUT4), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n463), .A2(new_n459), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G1gat), .B(G29gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT0), .ZN(new_n470));
  XNOR2_X1  g269(.A(G57gat), .B(G85gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  OR2_X1    g271(.A1(new_n457), .A2(new_n464), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT4), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n460), .A2(KEYINPUT5), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n473), .A2(new_n463), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n468), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n472), .B1(new_n468), .B2(new_n477), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n468), .A2(new_n477), .ZN(new_n483));
  INV_X1    g282(.A(new_n472), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G8gat), .B(G36gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(G64gat), .B(G92gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G226gat), .ZN(new_n490));
  INV_X1    g289(.A(G233gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G183gat), .A2(G190gat), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(KEYINPUT24), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(KEYINPUT24), .ZN(new_n495));
  OAI22_X1  g294(.A1(new_n494), .A2(new_n495), .B1(G183gat), .B2(G190gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(G169gat), .A2(G176gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT23), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G169gat), .B2(G176gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(G169gat), .A2(G176gat), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n502), .A3(KEYINPUT25), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n504));
  NOR2_X1   g303(.A1(G183gat), .A2(G190gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT64), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n493), .B(KEYINPUT24), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n503), .B1(new_n509), .B2(KEYINPUT25), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT26), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G176gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n358), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(KEYINPUT65), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(new_n497), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n511), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT66), .A3(new_n493), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G183gat), .ZN(new_n523));
  INV_X1    g322(.A(G190gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G183gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT27), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT27), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(G183gat), .ZN(new_n529));
  AND4_X1   g328(.A1(new_n522), .A2(new_n527), .A3(new_n529), .A4(new_n524), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT66), .B1(new_n520), .B2(new_n493), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n510), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n492), .B1(new_n534), .B2(new_n411), .ZN(new_n535));
  INV_X1    g334(.A(new_n492), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n493), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT66), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n521), .A3(new_n531), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n536), .B1(new_n540), .B2(new_n510), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n535), .A2(new_n409), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT73), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT29), .B1(new_n540), .B2(new_n510), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(new_n492), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n534), .A2(new_n411), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(KEYINPUT73), .A3(new_n536), .ZN(new_n547));
  INV_X1    g346(.A(new_n541), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n489), .B(new_n542), .C1(new_n549), .C2(new_n409), .ZN(new_n550));
  OAI22_X1  g349(.A1(new_n482), .A2(new_n486), .B1(KEYINPUT30), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(KEYINPUT30), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n409), .ZN(new_n554));
  INV_X1    g353(.A(new_n542), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n553), .B1(new_n556), .B2(new_n489), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n542), .B1(new_n549), .B2(new_n409), .ZN(new_n558));
  INV_X1    g357(.A(new_n489), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n558), .A2(KEYINPUT74), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n552), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n551), .B1(new_n561), .B2(KEYINPUT75), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT74), .B1(new_n558), .B2(new_n559), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n541), .B1(new_n535), .B2(KEYINPUT73), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n410), .B1(new_n564), .B2(new_n545), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n553), .B(new_n489), .C1(new_n565), .C2(new_n542), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n563), .A2(new_n566), .B1(KEYINPUT30), .B2(new_n550), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n432), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT71), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n450), .B(new_n510), .C1(new_n532), .C2(new_n533), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n450), .B1(new_n540), .B2(new_n510), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n534), .A2(new_n456), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(KEYINPUT70), .A3(new_n573), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n576), .A2(new_n578), .B1(G227gat), .B2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT34), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n571), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G227gat), .A2(G233gat), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n577), .A2(KEYINPUT70), .A3(new_n573), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT70), .B1(new_n577), .B2(new_n573), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n577), .A2(new_n573), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n580), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT72), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT72), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n587), .A2(new_n590), .A3(new_n580), .A4(new_n582), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n581), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n577), .A2(G227gat), .A3(G233gat), .A4(new_n573), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(KEYINPUT32), .ZN(new_n597));
  XOR2_X1   g396(.A(G15gat), .B(G43gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT69), .ZN(new_n599));
  XNOR2_X1  g398(.A(G71gat), .B(G99gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n594), .B(KEYINPUT32), .C1(new_n595), .C2(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n593), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n607), .A2(new_n586), .A3(new_n581), .A4(new_n592), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n608), .A3(KEYINPUT36), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT36), .B1(new_n606), .B2(new_n608), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n377), .B1(new_n570), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n432), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n483), .A2(new_n484), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(new_n479), .A3(new_n478), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n558), .A2(new_n559), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT30), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n616), .A2(new_n485), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n567), .B2(new_n568), .ZN(new_n620));
  AOI221_X4 g419(.A(KEYINPUT75), .B1(new_n550), .B2(KEYINPUT30), .C1(new_n563), .C2(new_n566), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n611), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n609), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n624), .A3(KEYINPUT80), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n452), .A2(new_n457), .A3(new_n459), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n626), .A2(KEYINPUT39), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n627), .A2(KEYINPUT82), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(KEYINPUT82), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n473), .A2(new_n463), .A3(new_n475), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n460), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(KEYINPUT39), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n472), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT40), .A4(new_n472), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n615), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n617), .A2(new_n618), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n567), .A2(KEYINPUT81), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT81), .B1(new_n567), .B2(new_n640), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n549), .A2(new_n410), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT37), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n535), .A2(new_n541), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n647), .B2(new_n409), .ZN(new_n648));
  AOI211_X1 g447(.A(KEYINPUT38), .B(new_n559), .C1(new_n645), .C2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT83), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n558), .B2(new_n646), .ZN(new_n651));
  NOR4_X1   g450(.A1(new_n565), .A2(KEYINPUT83), .A3(KEYINPUT37), .A4(new_n542), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n616), .A2(new_n485), .A3(new_n617), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n554), .A2(new_n646), .A3(new_n555), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT83), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n558), .A2(new_n650), .A3(new_n646), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n559), .B1(new_n556), .B2(KEYINPUT37), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT38), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n614), .B1(new_n656), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n644), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n613), .A2(new_n625), .A3(new_n665), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n552), .B(new_n640), .C1(new_n557), .C2(new_n560), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT81), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n606), .A2(new_n608), .A3(new_n432), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n482), .A2(new_n486), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(KEYINPUT35), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n669), .A2(new_n670), .A3(new_n641), .A4(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n606), .A2(new_n608), .A3(new_n432), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n620), .A2(new_n621), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT35), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n305), .B(new_n376), .C1(new_n666), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n671), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g479(.A1(new_n642), .A2(new_n643), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n683), .B2(G8gat), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n687), .B2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(G15gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n606), .ZN(new_n693));
  INV_X1    g492(.A(new_n608), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n678), .A2(new_n612), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n692), .ZN(G1326gat));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n614), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NAND2_X1  g500(.A1(new_n666), .A2(new_n677), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n244), .A2(new_n376), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n702), .A2(new_n303), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n249), .A3(new_n671), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n702), .B2(new_n303), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n638), .B1(new_n669), .B2(new_n641), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n660), .B2(new_n661), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n432), .B1(new_n712), .B2(new_n655), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n622), .B(new_n624), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n714), .A2(new_n677), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n714), .B2(new_n677), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n303), .A2(new_n708), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n703), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n722), .B(new_n703), .C1(new_n709), .C2(new_n719), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(new_n671), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n707), .B1(new_n724), .B2(new_n249), .ZN(G1328gat));
  NAND3_X1  g524(.A1(new_n704), .A2(new_n250), .A3(new_n682), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT46), .Z(new_n727));
  AND3_X1   g526(.A1(new_n721), .A2(new_n682), .A3(new_n723), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n250), .B2(new_n728), .ZN(G1329gat));
  OAI21_X1  g528(.A(G43gat), .B1(new_n720), .B2(new_n624), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  INV_X1    g530(.A(new_n695), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n704), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n612), .A3(new_n723), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n738), .A2(G43gat), .B1(new_n704), .B2(new_n733), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n736), .B(new_n737), .C1(KEYINPUT47), .C2(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n721), .A2(new_n614), .A3(new_n723), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n743), .A3(G50gat), .ZN(new_n744));
  INV_X1    g543(.A(G50gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n704), .A2(new_n745), .A3(new_n614), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n742), .B2(G50gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n741), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G50gat), .B1(new_n720), .B2(new_n432), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(KEYINPUT48), .A3(new_n746), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1331gat));
  NOR2_X1   g551(.A1(new_n716), .A2(new_n717), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n305), .A2(new_n375), .A3(new_n339), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n671), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n682), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n760), .B2(new_n759), .ZN(G1333gat));
  NAND3_X1  g562(.A1(new_n756), .A2(G71gat), .A3(new_n612), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n755), .A2(new_n732), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(G71gat), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g566(.A1(new_n755), .A2(new_n432), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT109), .B(G78gat), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n244), .A2(new_n375), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n304), .B1(new_n714), .B2(new_n677), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(KEYINPUT110), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(KEYINPUT111), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n774), .A3(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT111), .B1(new_n776), .B2(new_n777), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT112), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n781), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n783), .A2(new_n779), .A3(new_n784), .A4(new_n778), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(new_n270), .A3(new_n671), .A4(new_n338), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n709), .A2(new_n719), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n788), .A2(new_n339), .A3(new_n772), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(new_n671), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n270), .B2(new_n790), .ZN(G1336gat));
  AOI21_X1  g590(.A(new_n271), .B1(new_n789), .B2(new_n682), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(KEYINPUT52), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n780), .A2(new_n781), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n682), .A2(new_n271), .A3(new_n338), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n776), .B(KEYINPUT51), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT52), .B1(new_n798), .B2(new_n792), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(G1337gat));
  NOR3_X1   g599(.A1(new_n339), .A2(G99gat), .A3(new_n732), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n789), .A2(new_n612), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G99gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1338gat));
  INV_X1    g604(.A(G106gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n789), .B2(new_n614), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n338), .A2(new_n806), .A3(new_n614), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n797), .A2(new_n809), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT53), .B1(new_n811), .B2(new_n807), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1339gat));
  INV_X1    g612(.A(new_n671), .ZN(new_n814));
  INV_X1    g613(.A(new_n244), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n330), .B2(new_n319), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT113), .B1(new_n318), .B2(new_n320), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  NOR4_X1   g620(.A1(new_n315), .A2(new_n821), .A3(new_n319), .A4(new_n317), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n333), .B1(new_n321), .B2(new_n817), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n330), .B2(new_n319), .ZN(new_n826));
  INV_X1    g625(.A(new_n822), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n819), .B1(new_n828), .B2(new_n818), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n816), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n334), .B(new_n335), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n820), .A2(new_n822), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n331), .A2(KEYINPUT54), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT114), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n823), .A4(new_n824), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n830), .A2(new_n375), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n364), .A2(new_n341), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n350), .A2(new_n353), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n360), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n338), .A2(new_n369), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n303), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n830), .A2(new_n303), .A3(new_n835), .A4(new_n831), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n369), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n815), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n375), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n244), .A2(new_n304), .A3(new_n848), .A4(new_n339), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n814), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n670), .A3(new_n681), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n848), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(KEYINPUT116), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n848), .A2(G113gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n851), .B2(new_n339), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n338), .A2(new_n444), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT117), .Z(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n853), .B2(new_n858), .ZN(G1341gat));
  NOR2_X1   g658(.A1(new_n851), .A2(new_n815), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(G127gat), .Z(G1342gat));
  NAND4_X1  g660(.A1(new_n850), .A2(new_n670), .A3(new_n681), .A4(new_n303), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(G134gat), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(G134gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n847), .A2(new_n849), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n614), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n432), .B1(new_n847), .B2(new_n849), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n681), .A2(new_n671), .A3(new_n624), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n868), .B2(new_n614), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n872), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n878), .A3(new_n375), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G141gat), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n612), .A2(new_n432), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT119), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n682), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n850), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(G141gat), .A3(new_n848), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT58), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n885), .B1(new_n879), .B2(G141gat), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT120), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(G141gat), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n879), .A2(KEYINPUT122), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n875), .A2(new_n878), .A3(new_n895), .A4(new_n375), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g696(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n898));
  NAND2_X1  g697(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n889), .B(new_n892), .C1(new_n897), .C2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  INV_X1    g700(.A(new_n884), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n901), .B(G148gat), .C1(new_n902), .C2(new_n338), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n844), .B(KEYINPUT123), .ZN(new_n904));
  INV_X1    g703(.A(new_n845), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n843), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n849), .B1(new_n906), .B2(new_n244), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n614), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n869), .A2(new_n870), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n339), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n876), .A2(new_n901), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n875), .A2(new_n878), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n901), .B1(new_n914), .B2(new_n339), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n903), .B1(new_n916), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g716(.A(G155gat), .B1(new_n914), .B2(new_n815), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n395), .A3(new_n244), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1346gat));
  OAI21_X1  g719(.A(G162gat), .B1(new_n914), .B2(new_n304), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n396), .A3(new_n303), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1347gat));
  NAND2_X1  g722(.A1(new_n682), .A2(new_n670), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n814), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n926), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n868), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n358), .B1(new_n928), .B2(new_n848), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n681), .A2(new_n671), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n847), .B2(new_n849), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n670), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n375), .A2(G169gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT125), .ZN(G1348gat));
  OAI21_X1  g735(.A(new_n513), .B1(new_n928), .B2(new_n339), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n338), .A2(G176gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT126), .Z(G1349gat));
  INV_X1    g739(.A(new_n933), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n526), .B1(new_n941), .B2(new_n244), .ZN(new_n942));
  INV_X1    g741(.A(new_n928), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n244), .A2(new_n523), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n933), .B2(new_n304), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n943), .A2(new_n524), .A3(new_n303), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1351gat));
  NOR2_X1   g749(.A1(new_n931), .A2(new_n612), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n951), .B1(new_n908), .B2(new_n909), .ZN(new_n952));
  INV_X1    g751(.A(G197gat), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n952), .A2(new_n953), .A3(new_n848), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n932), .A2(new_n881), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n375), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n954), .A2(new_n957), .ZN(G1352gat));
  NAND2_X1  g757(.A1(new_n911), .A2(new_n951), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G204gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n955), .A2(G204gat), .A3(new_n339), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT62), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n956), .A2(new_n404), .A3(new_n244), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n244), .B(new_n951), .C1(new_n908), .C2(new_n909), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g768(.A(KEYINPUT127), .B(KEYINPUT63), .C1(new_n965), .C2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n952), .B2(new_n304), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n405), .A3(new_n303), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


