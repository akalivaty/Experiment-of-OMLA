//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G104), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G107), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n198), .A3(G104), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n198), .A2(G104), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT79), .A2(G101), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT79), .A2(G101), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n204), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n205), .A2(new_n207), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT79), .A2(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT79), .A2(G101), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n201), .A3(new_n216), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n214), .A2(new_n217), .A3(KEYINPUT80), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n197), .B(new_n203), .C1(new_n213), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT83), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT5), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n194), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G116), .B(G119), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(G113), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n220), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n194), .A2(new_n222), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT66), .B1(new_n191), .B2(new_n193), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT5), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n227), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(KEYINPUT83), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n219), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n205), .A2(new_n207), .A3(new_n201), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G101), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n213), .B2(new_n218), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n223), .A2(new_n225), .A3(new_n195), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n197), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n235), .A3(G101), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n189), .B1(new_n234), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n228), .A2(new_n233), .ZN(new_n244));
  INV_X1    g058(.A(new_n219), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n240), .A2(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n238), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n248), .A3(new_n188), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n249), .A3(KEYINPUT6), .ZN(new_n250));
  INV_X1    g064(.A(G125), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT64), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  AOI21_X1  g072(.A(G146), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n254), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n256), .A2(new_n258), .A3(G146), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n255), .A2(G146), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n252), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n251), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(G128), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n259), .B2(new_n261), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(new_n265), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n251), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G224), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n280), .B(new_n189), .C1(new_n234), .C2(new_n242), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n250), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n278), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n283), .A4(new_n275), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(KEYINPUT7), .ZN(new_n285));
  INV_X1    g099(.A(new_n275), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n267), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n244), .A2(new_n245), .B1(new_n247), .B2(new_n238), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(new_n188), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n188), .B(KEYINPUT8), .ZN(new_n291));
  INV_X1    g105(.A(new_n203), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n208), .A2(new_n212), .A3(new_n204), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT80), .B1(new_n214), .B2(new_n217), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n244), .B2(new_n197), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n227), .B1(KEYINPUT5), .B2(new_n224), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n219), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n291), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n290), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n282), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT84), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n282), .B2(new_n300), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n282), .A2(new_n300), .A3(new_n306), .A4(new_n301), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G475), .ZN(new_n309));
  XNOR2_X1  g123(.A(G113), .B(G122), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(new_n200), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  AND2_X1   g126(.A1(KEYINPUT68), .A2(G237), .ZN(new_n313));
  NOR2_X1   g127(.A1(KEYINPUT68), .A2(G237), .ZN(new_n314));
  OAI211_X1 g128(.A(G214), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT64), .B(G143), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n315), .A2(KEYINPUT85), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT85), .ZN(new_n318));
  AOI21_X1  g132(.A(G143), .B1(new_n257), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G131), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT17), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n315), .A2(KEYINPUT85), .A3(new_n316), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n323), .B(new_n324), .C1(new_n315), .C2(new_n319), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT75), .B1(new_n251), .B2(G140), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT74), .B(G140), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(new_n251), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n330), .A2(KEYINPUT74), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(KEYINPUT74), .ZN(new_n332));
  OAI211_X1 g146(.A(KEYINPUT75), .B(G125), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT16), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n251), .B2(G140), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n260), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n336), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G146), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT17), .B(G131), .C1(new_n317), .C2(new_n320), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n326), .A2(new_n337), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT18), .A2(G131), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n317), .B2(new_n320), .ZN(new_n343));
  INV_X1    g157(.A(new_n342), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n323), .B(new_n344), .C1(new_n315), .C2(new_n319), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n329), .A2(G146), .A3(new_n333), .ZN(new_n347));
  XNOR2_X1  g161(.A(G125), .B(G140), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n260), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n347), .A2(KEYINPUT86), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT86), .B1(new_n347), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n311), .B1(new_n341), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n311), .A3(new_n352), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G902), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n309), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(G475), .A2(G902), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n341), .A2(new_n311), .A3(new_n352), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n329), .A2(KEYINPUT19), .A3(new_n333), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT19), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT87), .B1(new_n348), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n329), .A2(new_n333), .A3(KEYINPUT87), .A4(KEYINPUT19), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n260), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n321), .A2(new_n325), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n339), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n311), .B1(new_n369), .B2(new_n352), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n359), .B1(new_n360), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n339), .ZN(new_n372));
  AOI21_X1  g186(.A(G146), .B1(new_n364), .B2(new_n365), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n352), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n311), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT88), .B1(new_n376), .B2(new_n355), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n371), .B1(new_n377), .B2(KEYINPUT20), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n355), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n379), .A2(KEYINPUT88), .A3(new_n380), .A4(new_n359), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n358), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G116), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n192), .A2(G122), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT89), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(G107), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n316), .A2(G128), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n272), .A2(G143), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G134), .ZN(new_n394));
  INV_X1    g208(.A(G134), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n395), .A3(new_n392), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n390), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n192), .A2(KEYINPUT14), .A3(G122), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n398), .A2(G107), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(KEYINPUT14), .B2(new_n386), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT91), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n399), .B(KEYINPUT91), .C1(KEYINPUT14), .C2(new_n386), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT90), .B(KEYINPUT13), .Z(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(G128), .A3(new_n316), .ZN(new_n407));
  OAI211_X1 g221(.A(G134), .B(new_n407), .C1(new_n393), .C2(new_n406), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n387), .A2(G107), .A3(new_n389), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(new_n396), .C1(new_n409), .C2(new_n390), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT71), .B(G217), .Z(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT9), .B(G234), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n412), .A2(G953), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n405), .A2(new_n410), .A3(new_n414), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT92), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n419), .A3(new_n415), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n357), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n423), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n418), .A2(new_n357), .A3(new_n420), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(G234), .A2(G237), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n428), .A2(G902), .A3(G953), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(G898), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n428), .A2(G952), .A3(new_n312), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT93), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n427), .A2(new_n436), .ZN(new_n437));
  AND4_X1   g251(.A1(new_n187), .A2(new_n308), .A3(new_n382), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n412), .B1(G234), .B2(new_n357), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n272), .A2(G119), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n190), .A2(G128), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT72), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT72), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT24), .B(G110), .Z(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT73), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT73), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n443), .A2(new_n449), .A3(new_n445), .A4(new_n446), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n272), .A2(KEYINPUT23), .A3(G119), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n190), .A2(G128), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n451), .B(new_n441), .C1(new_n452), .C2(KEYINPUT23), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n448), .A2(new_n450), .B1(G110), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n337), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n260), .B1(new_n334), .B2(new_n336), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT76), .ZN(new_n458));
  OR3_X1    g272(.A1(new_n453), .A2(new_n458), .A3(G110), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n458), .B1(new_n453), .B2(G110), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n443), .A2(new_n445), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n446), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n339), .A3(new_n349), .ZN(new_n463));
  INV_X1    g277(.A(G137), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT22), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT22), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G137), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT77), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT22), .B(G137), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT77), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT78), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n312), .A2(G221), .A3(G234), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT78), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n474), .B2(new_n477), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n457), .A2(new_n463), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n457), .B2(new_n463), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT25), .B1(new_n483), .B2(new_n357), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n457), .A2(new_n463), .ZN(new_n485));
  INV_X1    g299(.A(new_n480), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n457), .A2(new_n463), .A3(new_n480), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(KEYINPUT25), .A3(new_n357), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n439), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n483), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n439), .A2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n491), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT28), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT67), .ZN(new_n498));
  OR2_X1    g312(.A1(KEYINPUT65), .A2(G137), .ZN(new_n499));
  AND2_X1   g313(.A1(KEYINPUT11), .A2(G134), .ZN(new_n500));
  NAND2_X1  g314(.A1(KEYINPUT65), .A2(G137), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT11), .A2(G134), .ZN(new_n503));
  NOR2_X1   g317(.A1(KEYINPUT11), .A2(G134), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n503), .B1(new_n504), .B2(G137), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n502), .A2(new_n324), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n324), .B1(new_n502), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n262), .A2(new_n266), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n498), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n261), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n316), .B2(G146), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n264), .B1(new_n316), .B2(G146), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n512), .A2(new_n254), .B1(new_n513), .B2(new_n252), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n502), .A2(new_n505), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G131), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n502), .A2(new_n505), .A3(new_n324), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n518), .A3(KEYINPUT67), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n499), .A2(new_n395), .A3(new_n501), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n324), .B1(G134), .B2(G137), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n271), .A2(new_n274), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n510), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n240), .ZN(new_n528));
  INV_X1    g342(.A(new_n240), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n510), .A2(new_n519), .A3(new_n529), .A4(new_n526), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n497), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n525), .ZN(new_n532));
  OAI22_X1  g346(.A1(new_n532), .A2(new_n523), .B1(new_n508), .B2(new_n509), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n497), .B1(new_n533), .B2(new_n240), .ZN(new_n534));
  OR2_X1    g348(.A1(KEYINPUT68), .A2(G237), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT68), .A2(G237), .ZN(new_n536));
  AOI21_X1  g350(.A(G953), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G210), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n538), .A2(KEYINPUT27), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(KEYINPUT27), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT26), .B(G101), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n534), .A2(new_n546), .A3(KEYINPUT29), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n357), .B1(new_n531), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n508), .A2(new_n509), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n523), .B1(new_n274), .B2(new_n271), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n240), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n530), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT28), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n514), .A2(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT28), .B1(new_n554), .B2(new_n529), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n544), .A2(new_n545), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n240), .B1(new_n554), .B2(KEYINPUT30), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n524), .B2(new_n525), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n510), .A2(new_n561), .A3(new_n519), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n530), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT29), .B1(new_n563), .B2(new_n556), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n548), .B1(new_n558), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G472), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n496), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n556), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n558), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n528), .A2(new_n530), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT28), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n555), .A2(new_n556), .A3(new_n569), .ZN(new_n573));
  AOI21_X1  g387(.A(G902), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT70), .A3(G472), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n530), .B(new_n546), .C1(new_n559), .C2(new_n562), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT31), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n497), .B1(new_n530), .B2(new_n551), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n556), .B1(new_n580), .B2(new_n555), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n533), .A2(new_n560), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n510), .A2(new_n561), .A3(new_n519), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n240), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n585));
  NAND4_X1  g399(.A1(new_n584), .A2(new_n530), .A3(new_n546), .A4(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n579), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(G472), .A2(G902), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n587), .A2(KEYINPUT32), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT32), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n495), .B1(new_n577), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT82), .B(G469), .Z(new_n593));
  OAI21_X1  g407(.A(new_n203), .B1(new_n213), .B2(new_n218), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n263), .A2(new_n265), .A3(new_n273), .ZN(new_n595));
  INV_X1    g409(.A(new_n513), .ZN(new_n596));
  OAI21_X1  g410(.A(G128), .B1(new_n259), .B2(new_n269), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n295), .A2(new_n525), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n518), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT12), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n532), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n257), .A2(G143), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n255), .A2(KEYINPUT64), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n260), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n272), .B1(new_n606), .B2(KEYINPUT1), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n274), .B1(new_n607), .B2(new_n513), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n295), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n508), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT12), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n262), .A2(new_n241), .A3(new_n266), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n271), .B2(new_n274), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n238), .A2(new_n613), .B1(new_n295), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n614), .B1(new_n594), .B2(new_n598), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n508), .ZN(new_n618));
  XNOR2_X1  g432(.A(G110), .B(G140), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n312), .A2(G227), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n619), .B(new_n620), .Z(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n602), .A2(new_n612), .A3(new_n618), .A4(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n618), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n508), .B1(new_n616), .B2(new_n617), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(G902), .B(new_n593), .C1(new_n623), .C2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n618), .B1(new_n611), .B2(new_n610), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n601), .A2(KEYINPUT12), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT81), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT81), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n602), .A2(new_n612), .A3(new_n632), .A4(new_n618), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n621), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n624), .A2(new_n625), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n622), .ZN(new_n636));
  AOI21_X1  g450(.A(G902), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G469), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n628), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G221), .ZN(new_n640));
  INV_X1    g454(.A(new_n413), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n357), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n438), .A2(new_n592), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n215), .A2(new_n216), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G3));
  NAND2_X1  g461(.A1(new_n587), .A2(new_n357), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(KEYINPUT94), .A3(G472), .ZN(new_n649));
  NAND2_X1  g463(.A1(KEYINPUT94), .A2(G472), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n587), .A2(new_n357), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n495), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n282), .A2(new_n300), .A3(new_n301), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n187), .B(new_n435), .C1(new_n654), .C2(new_n304), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT33), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n418), .A2(new_n656), .A3(new_n420), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n416), .A2(KEYINPUT33), .A3(new_n417), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n422), .A2(G902), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n421), .A2(new_n422), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n655), .A2(new_n382), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n644), .A2(new_n653), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  AND2_X1   g480(.A1(new_n424), .A2(new_n426), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n357), .B1(new_n360), .B2(new_n353), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n371), .A2(new_n380), .B1(new_n668), .B2(G475), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n379), .A2(KEYINPUT20), .A3(new_n359), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n655), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n644), .A2(new_n653), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT35), .B(G107), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  NAND2_X1  g489(.A1(new_n485), .A2(KEYINPUT95), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n486), .A2(KEYINPUT36), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT95), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n457), .A2(new_n463), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n677), .B1(new_n676), .B2(new_n679), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n493), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n491), .A2(KEYINPUT96), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT96), .ZN(new_n685));
  INV_X1    g499(.A(new_n439), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n487), .A2(new_n357), .A3(new_n488), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT25), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n686), .B1(new_n689), .B2(new_n489), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n676), .A2(new_n679), .ZN(new_n691));
  INV_X1    g505(.A(new_n677), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n494), .B1(new_n693), .B2(new_n680), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n685), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n684), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n652), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n438), .A2(new_n697), .A3(new_n644), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n187), .B1(new_n654), .B2(new_n304), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT97), .B(G900), .Z(new_n704));
  AND2_X1   g518(.A1(new_n704), .A2(new_n429), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT98), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n433), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n671), .A2(new_n667), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT70), .B1(new_n575), .B2(G472), .ZN(new_n712));
  AOI211_X1 g526(.A(new_n496), .B(new_n566), .C1(new_n570), .C2(new_n574), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n590), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n587), .A2(KEYINPUT32), .A3(new_n588), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n703), .B(new_n711), .C1(new_n714), .C2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n639), .A2(new_n643), .A3(new_n695), .A4(new_n684), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n701), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n643), .A2(new_n639), .A3(new_n695), .A4(new_n684), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n702), .B1(new_n577), .B2(new_n591), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(KEYINPUT99), .A3(new_n722), .A4(new_n711), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  XNOR2_X1  g539(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n709), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n644), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(new_n728), .B(KEYINPUT103), .Z(new_n729));
  OR2_X1    g543(.A1(new_n729), .A2(KEYINPUT40), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n571), .A2(new_n556), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT100), .A3(new_n578), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n357), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT100), .B1(new_n731), .B2(new_n578), .ZN(new_n734));
  OAI21_X1  g548(.A(G472), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n715), .A2(new_n735), .A3(new_n716), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n690), .A2(new_n694), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n736), .A2(new_n187), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n378), .A2(new_n381), .ZN(new_n739));
  INV_X1    g553(.A(new_n358), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n308), .B(KEYINPUT38), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n738), .A2(new_n741), .A3(new_n427), .A4(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(KEYINPUT101), .Z(new_n744));
  NAND2_X1  g558(.A1(new_n729), .A2(KEYINPUT40), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n730), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(new_n316), .Z(G45));
  NOR3_X1   g561(.A1(new_n382), .A2(new_n662), .A3(new_n710), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n703), .C1(new_n714), .C2(new_n717), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n719), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n260), .ZN(G48));
  AOI21_X1  g565(.A(G902), .B1(new_n623), .B2(new_n626), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT104), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n638), .B1(new_n752), .B2(KEYINPUT104), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n642), .B(new_n627), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n592), .A2(new_n663), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT41), .B(G113), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G15));
  NAND3_X1  g572(.A1(new_n592), .A2(new_n672), .A3(new_n755), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  AND4_X1   g574(.A1(new_n382), .A2(new_n684), .A3(new_n695), .A4(new_n437), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n722), .A2(new_n761), .A3(new_n755), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  INV_X1    g577(.A(new_n588), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n579), .A2(new_n586), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n556), .B1(new_n531), .B2(new_n555), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n566), .B1(new_n587), .B2(new_n357), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n495), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n702), .A2(new_n382), .A3(new_n667), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n435), .A4(new_n755), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  NOR3_X1   g586(.A1(new_n737), .A2(new_n767), .A3(new_n768), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n755), .A2(new_n773), .A3(new_n748), .A4(new_n703), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  INV_X1    g589(.A(new_n187), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n282), .A2(new_n300), .ZN(new_n777));
  INV_X1    g591(.A(new_n301), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n303), .A3(new_n643), .A4(new_n307), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n634), .A2(KEYINPUT105), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n602), .A2(new_n618), .A3(new_n612), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n622), .B1(new_n782), .B2(KEYINPUT81), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n783), .A2(new_n633), .B1(new_n635), .B2(new_n622), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n781), .B(G469), .C1(new_n784), .C2(KEYINPUT105), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n638), .A2(new_n357), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n627), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n780), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n592), .A3(new_n748), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT42), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n788), .A2(new_n592), .A3(KEYINPUT42), .A4(new_n748), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(KEYINPUT106), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT106), .B1(new_n791), .B2(new_n792), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G131), .ZN(G33));
  NAND3_X1  g611(.A1(new_n788), .A2(new_n592), .A3(new_n711), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G134), .ZN(G36));
  OAI211_X1 g613(.A(KEYINPUT45), .B(new_n781), .C1(new_n784), .C2(KEYINPUT105), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n800), .B(G469), .C1(KEYINPUT45), .C2(new_n784), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n786), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n628), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n643), .B(new_n727), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT107), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n807), .A2(KEYINPUT43), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(KEYINPUT43), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n660), .A2(new_n661), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n382), .A2(new_n811), .ZN(new_n812));
  MUX2_X1   g626(.A(new_n810), .B(new_n809), .S(new_n812), .Z(new_n813));
  AOI21_X1  g627(.A(new_n737), .B1(new_n651), .B2(new_n649), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT44), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(KEYINPUT44), .A3(new_n814), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n779), .A2(new_n303), .A3(new_n307), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n806), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(new_n464), .ZN(G39));
  OAI21_X1  g635(.A(new_n643), .B1(new_n804), .B2(new_n805), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n643), .B(new_n823), .C1(new_n804), .C2(new_n805), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n714), .A2(new_n717), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n827), .A2(new_n495), .A3(new_n748), .A4(new_n818), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  NAND3_X1  g644(.A1(new_n813), .A2(new_n432), .A3(new_n769), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n753), .A2(new_n754), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n628), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n742), .A2(new_n642), .A3(new_n187), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT50), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n834), .A2(new_n780), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n813), .A2(new_n432), .A3(new_n773), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT112), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n736), .A2(new_n495), .A3(new_n433), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n838), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n382), .A3(new_n662), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n834), .A2(new_n643), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n825), .B2(new_n826), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n831), .A2(new_n817), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n846), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n832), .A2(new_n703), .A3(new_n755), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n843), .A2(new_n741), .A3(new_n811), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(G952), .A3(new_n312), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n813), .A2(new_n592), .A3(new_n432), .A4(new_n838), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT48), .Z(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n837), .A2(new_n852), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n845), .A2(KEYINPUT113), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n845), .A2(KEYINPUT113), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n848), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(KEYINPUT114), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n850), .B1(new_n865), .B2(KEYINPUT114), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT115), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n720), .A2(new_n723), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n785), .A2(new_n787), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n690), .A2(new_n694), .A3(new_n642), .A4(new_n710), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n770), .A2(new_n872), .A3(new_n873), .A4(new_n736), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n874), .B(new_n774), .C1(new_n749), .C2(new_n719), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n870), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n724), .A3(KEYINPUT52), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n756), .A2(new_n762), .A3(new_n759), .A4(new_n771), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n741), .A2(KEYINPUT110), .A3(new_n811), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT110), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n382), .B2(new_n662), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n382), .A2(new_n427), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n308), .A2(new_n187), .A3(new_n435), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n644), .A3(new_n653), .A4(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n887), .A2(new_n645), .A3(new_n698), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n667), .A2(new_n670), .A3(new_n669), .A4(new_n709), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n577), .B2(new_n591), .ZN(new_n890));
  INV_X1    g704(.A(new_n696), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n644), .A3(new_n891), .A4(new_n818), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n788), .A2(new_n748), .A3(new_n773), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n892), .A2(new_n798), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n880), .A2(new_n888), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n879), .A2(new_n796), .A3(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT53), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(KEYINPUT53), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(KEYINPUT54), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n877), .A2(new_n724), .A3(KEYINPUT52), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT52), .B1(new_n877), .B2(new_n724), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n762), .A2(new_n756), .A3(new_n759), .A4(new_n771), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n887), .A2(new_n698), .A3(new_n645), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n791), .A2(new_n792), .ZN(new_n906));
  AND4_X1   g720(.A1(KEYINPUT53), .A2(new_n892), .A3(new_n798), .A4(new_n893), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT111), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n906), .A2(new_n907), .A3(new_n880), .A4(new_n888), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT111), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n879), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n909), .A2(new_n912), .B1(new_n896), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n869), .A2(new_n899), .A3(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n860), .A2(new_n868), .A3(KEYINPUT115), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n917), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  OR4_X1    g733(.A1(new_n495), .A2(new_n812), .A3(new_n642), .A4(new_n776), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT109), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n742), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n834), .A2(KEYINPUT49), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n834), .A2(KEYINPUT49), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n736), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(new_n925), .C1(new_n921), .C2(new_n920), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n926), .ZN(G75));
  NOR2_X1   g741(.A1(new_n312), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n914), .A2(new_n357), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(G210), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n250), .A2(new_n281), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n279), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT55), .Z(new_n935));
  XOR2_X1   g749(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n936));
  OR2_X1    g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n929), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n931), .B2(KEYINPUT116), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(KEYINPUT116), .B2(new_n931), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(new_n935), .ZN(G51));
  INV_X1    g755(.A(new_n795), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n905), .A3(new_n793), .A4(new_n894), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n913), .B1(new_n902), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n879), .A2(new_n910), .A3(new_n911), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n911), .B1(new_n879), .B2(new_n910), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT54), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n916), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n786), .B(KEYINPUT57), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n951), .A2(KEYINPUT118), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n623), .A2(new_n626), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(KEYINPUT118), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n930), .A2(new_n802), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n928), .B1(new_n955), .B2(new_n956), .ZN(G54));
  NAND3_X1  g771(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n958));
  INV_X1    g772(.A(new_n379), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n958), .A2(KEYINPUT119), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT119), .B1(new_n958), .B2(new_n959), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n928), .B1(new_n958), .B2(new_n959), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT59), .Z(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n916), .B2(new_n899), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n657), .B2(new_n658), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n657), .A2(new_n658), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n965), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n928), .B(new_n967), .C1(new_n949), .C2(new_n969), .ZN(G63));
  INV_X1    g784(.A(KEYINPUT120), .ZN(new_n971));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT60), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n914), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n947), .A2(KEYINPUT120), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n976), .A3(new_n492), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n929), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n974), .A2(new_n976), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n681), .A2(new_n682), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT121), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT121), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n983), .B(new_n980), .C1(new_n974), .C2(new_n976), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n978), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT122), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n982), .B2(new_n984), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI221_X1 g803(.A(new_n978), .B1(new_n986), .B2(KEYINPUT61), .C1(new_n982), .C2(new_n984), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G66));
  OAI21_X1  g805(.A(G953), .B1(new_n430), .B2(new_n277), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n905), .B(KEYINPUT123), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n994), .B2(G953), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n933), .B1(G898), .B2(new_n312), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G69));
  INV_X1    g811(.A(new_n806), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n592), .A3(new_n770), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n796), .A2(new_n798), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n999), .A2(new_n1000), .A3(new_n829), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT125), .ZN(new_n1003));
  INV_X1    g817(.A(new_n774), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n750), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n724), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1003), .B1(new_n820), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1006), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n819), .A2(new_n815), .ZN(new_n1009));
  OAI211_X1 g823(.A(KEYINPUT125), .B(new_n1008), .C1(new_n1009), .C2(new_n806), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(G953), .B1(new_n1002), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n312), .A2(G900), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(KEYINPUT126), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n582), .A2(new_n583), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(new_n366), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT124), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n746), .A2(new_n1008), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n885), .A2(new_n592), .A3(new_n818), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n729), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n820), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1025), .A2(new_n829), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n312), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1023), .B1(new_n1031), .B2(new_n1020), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n312), .B1(G227), .B2(G900), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n1022), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1033), .B1(new_n1022), .B2(new_n1032), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1034), .A2(new_n1035), .ZN(G72));
  NAND2_X1  g850(.A1(new_n563), .A2(new_n546), .ZN(new_n1037));
  OR2_X1    g851(.A1(new_n1030), .A2(new_n993), .ZN(new_n1038));
  NAND2_X1  g852(.A1(G472), .A2(G902), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1039), .B(KEYINPUT63), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT127), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1037), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1002), .A2(new_n1011), .A3(new_n994), .ZN(new_n1043));
  AOI211_X1 g857(.A(new_n546), .B(new_n563), .C1(new_n1043), .C2(new_n1041), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n897), .A2(new_n898), .ZN(new_n1045));
  AOI211_X1 g859(.A(new_n1040), .B(new_n1045), .C1(new_n578), .C2(new_n568), .ZN(new_n1046));
  NOR4_X1   g860(.A1(new_n1042), .A2(new_n928), .A3(new_n1044), .A4(new_n1046), .ZN(G57));
endmodule


