//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  AND2_X1   g002(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT28), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n208), .B(new_n203), .C1(new_n205), .C2(new_n204), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n210), .A2(new_n211), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n222), .A2(new_n223), .A3(new_n216), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT64), .A4(KEYINPUT23), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n203), .ZN(new_n232));
  NAND3_X1  g031(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n224), .A2(new_n227), .A3(new_n228), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n211), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT24), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n211), .A2(new_n237), .A3(new_n229), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n231), .A2(new_n203), .A3(KEYINPUT66), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n239), .A2(new_n240), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n225), .A2(new_n222), .A3(new_n216), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n223), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n202), .B1(new_n236), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n240), .B1(new_n229), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n243), .A2(new_n242), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n245), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT25), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(KEYINPUT77), .A3(new_n220), .A4(new_n235), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n248), .B(KEYINPUT76), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n236), .A2(new_n246), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT29), .ZN(new_n259));
  INV_X1    g058(.A(G197gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT75), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(G204gat), .ZN(new_n262));
  INV_X1    g061(.A(G204gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT75), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n260), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT22), .ZN(new_n266));
  INV_X1    g065(.A(G211gat), .ZN(new_n267));
  INV_X1    g066(.A(G218gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(KEYINPUT75), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n261), .A2(G204gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(G197gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n265), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n276), .A2(new_n269), .A3(new_n265), .A4(new_n272), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n259), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n258), .A2(new_n257), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n247), .A2(new_n282), .A3(new_n255), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n283), .B2(new_n248), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n284), .B2(new_n279), .ZN(new_n285));
  XOR2_X1   g084(.A(G8gat), .B(G36gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(G64gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G92gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT79), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n285), .A2(new_n292), .A3(new_n288), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(KEYINPUT30), .A3(new_n288), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n288), .B(KEYINPUT78), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(new_n280), .C1(new_n284), .C2(new_n279), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n300));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301));
  INV_X1    g100(.A(G113gat), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT68), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G120gat), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n303), .A2(G113gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n300), .B(new_n301), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n301), .ZN(new_n310));
  XNOR2_X1  g109(.A(G113gat), .B(G120gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(KEYINPUT1), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT80), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G141gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(G148gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT80), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n326), .A2(new_n320), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT81), .B(G141gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n322), .B1(new_n330), .B2(new_n317), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n320), .B1(new_n326), .B2(KEYINPUT2), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n329), .B1(new_n328), .B2(new_n333), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT4), .B(new_n313), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n328), .A2(new_n333), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n309), .A2(new_n312), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n325), .A2(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n338), .B2(new_n340), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n336), .A2(new_n337), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n341), .B(new_n340), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n348), .A2(new_n337), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT5), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n338), .A2(new_n345), .A3(new_n340), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n337), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(KEYINPUT5), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n328), .A2(new_n342), .A3(new_n333), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n342), .B1(new_n328), .B2(new_n333), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n345), .B1(new_n357), .B2(new_n340), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n338), .A2(KEYINPUT82), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n329), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n340), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n352), .B(new_n354), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G1gat), .B(G29gat), .Z(new_n363));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n367), .B1(new_n350), .B2(new_n362), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI211_X1 g171(.A(new_n369), .B(new_n367), .C1(new_n350), .C2(new_n362), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n294), .B(new_n299), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n275), .B2(new_n277), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n342), .B1(new_n376), .B2(KEYINPUT84), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n378));
  AOI211_X1 g177(.A(new_n378), .B(KEYINPUT29), .C1(new_n275), .C2(new_n277), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n338), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n279), .B1(new_n355), .B2(KEYINPUT29), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n359), .A2(new_n360), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n341), .B2(new_n342), .ZN(new_n387));
  OAI22_X1  g186(.A1(new_n385), .A2(new_n386), .B1(new_n278), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n381), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G22gat), .ZN(new_n391));
  INV_X1    g190(.A(G22gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n384), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT31), .B(G50gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n391), .A2(KEYINPUT85), .A3(new_n393), .A4(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n400), .A2(new_n396), .B1(new_n391), .B2(new_n393), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n375), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n396), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n391), .A2(new_n393), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT86), .A3(new_n397), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n374), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n313), .B1(new_n236), .B2(new_n246), .ZN(new_n408));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n254), .A2(new_n340), .A3(new_n220), .A4(new_n235), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n413));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G15gat), .B(G43gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G71gat), .ZN(new_n418));
  INV_X1    g217(.A(G99gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT70), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n416), .A2(KEYINPUT70), .A3(new_n420), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n418), .B(G99gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT71), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(KEYINPUT71), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n413), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(KEYINPUT32), .A3(new_n412), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n408), .A2(new_n411), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n409), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT34), .B1(new_n410), .B2(KEYINPUT72), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n435), .A2(new_n423), .A3(new_n424), .A4(new_n430), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(KEYINPUT74), .A3(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n435), .A4(new_n430), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT36), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n437), .A2(new_n438), .ZN(new_n447));
  OAI22_X1  g246(.A1(new_n443), .A2(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n407), .A2(KEYINPUT87), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n367), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT39), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n352), .B1(new_n358), .B2(new_n361), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n353), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n348), .A2(new_n337), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n353), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n455), .A2(KEYINPUT89), .A3(KEYINPUT40), .A4(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n344), .A2(KEYINPUT4), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n385), .A2(new_n313), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n351), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(KEYINPUT39), .B(new_n454), .C1(new_n462), .C2(new_n337), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n457), .A3(new_n367), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n294), .A2(new_n299), .B1(new_n465), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n350), .A2(new_n362), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n450), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n372), .A2(new_n373), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n285), .A2(new_n292), .A3(new_n288), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n292), .B1(new_n285), .B2(new_n288), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n476), .B(new_n280), .C1(new_n284), .C2(new_n279), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n256), .A2(new_n259), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n278), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT90), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n481), .A3(new_n278), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n284), .B2(new_n278), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n477), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(new_n296), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n285), .A2(KEYINPUT37), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n488), .A2(new_n477), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT38), .B1(new_n489), .B2(new_n288), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n472), .A2(new_n475), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n398), .A2(new_n401), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n471), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT87), .B1(new_n407), .B2(new_n448), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n449), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n298), .B1(new_n475), .B2(new_n291), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n470), .A2(new_n369), .A3(new_n368), .ZN(new_n498));
  INV_X1    g297(.A(new_n373), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n497), .A2(new_n443), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n398), .B2(new_n401), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(KEYINPUT91), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n497), .A2(new_n443), .A3(new_n500), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(new_n503), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n447), .B1(new_n405), .B2(new_n397), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(new_n500), .A3(new_n497), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n505), .A2(new_n508), .B1(KEYINPUT35), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n496), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n513), .A2(G1gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT16), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n515), .B2(G1gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g320(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n514), .A2(new_n516), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n526), .A2(G71gat), .A3(G78gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n525), .A2(new_n531), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n532), .A2(new_n533), .A3(new_n526), .ZN(new_n534));
  XNOR2_X1  g333(.A(G71gat), .B(G78gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT21), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n524), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G183gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(G127gat), .B(G155gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT98), .B(G211gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n536), .A2(new_n537), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n548), .B(new_n549), .Z(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n546), .B2(new_n547), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT99), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT99), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(G85gat), .A3(G92gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT7), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT7), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G99gat), .B(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n561), .A2(new_n568), .A3(new_n565), .A4(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT100), .Z(new_n573));
  NAND2_X1  g372(.A1(G29gat), .A2(G36gat), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR3_X1   g375(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(G43gat), .B(G50gat), .ZN(new_n578));
  OAI221_X1 g377(.A(new_n574), .B1(new_n576), .B2(new_n577), .C1(new_n578), .C2(KEYINPUT15), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(KEYINPUT15), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT17), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n579), .A2(KEYINPUT15), .A3(new_n578), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n579), .B1(KEYINPUT15), .B2(new_n578), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n573), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G190gat), .B(G218gat), .Z(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n581), .ZN(new_n590));
  INV_X1    g389(.A(new_n572), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT101), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n587), .A2(new_n589), .A3(new_n592), .ZN(new_n599));
  INV_X1    g398(.A(new_n588), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n593), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT102), .B1(new_n554), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n553), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n551), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n603), .A2(new_n604), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT107), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n214), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n263), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT106), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n567), .A2(KEYINPUT104), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT104), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n561), .A2(new_n620), .A3(new_n565), .A4(new_n566), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n568), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n536), .B1(new_n623), .B2(KEYINPUT105), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n571), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT103), .B1(new_n536), .B2(new_n572), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n536), .A2(new_n572), .A3(KEYINPUT103), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n627), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n536), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n591), .A3(KEYINPUT10), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n618), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n626), .A2(new_n571), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n622), .B2(new_n625), .ZN(new_n638));
  INV_X1    g437(.A(new_n630), .ZN(new_n639));
  OAI22_X1  g438(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(new_n628), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n618), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n613), .B(new_n616), .C1(new_n636), .C2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n635), .B1(new_n640), .B2(KEYINPUT10), .ZN(new_n645));
  INV_X1    g444(.A(new_n618), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n641), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n616), .B1(new_n648), .B2(new_n613), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n582), .A2(new_n586), .A3(new_n524), .ZN(new_n651));
  NAND2_X1  g450(.A1(G229gat), .A2(G233gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n524), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n590), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n581), .B2(new_n524), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n652), .B(KEYINPUT94), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT13), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n590), .A2(new_n653), .A3(new_n658), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n651), .A2(KEYINPUT18), .A3(new_n652), .A4(new_n654), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n657), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT11), .B(G169gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G197gat), .ZN(new_n668));
  XOR2_X1   g467(.A(G113gat), .B(G141gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT12), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT92), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT96), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n657), .A2(new_n671), .A3(new_n664), .A4(new_n665), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n666), .A2(new_n676), .A3(new_n672), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  AND4_X1   g477(.A1(new_n512), .A2(new_n612), .A3(new_n650), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n472), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT108), .B(G1gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1324gat));
  NAND2_X1  g481(.A1(new_n294), .A2(new_n299), .ZN(new_n683));
  NAND2_X1  g482(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n515), .A2(new_n519), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n679), .A2(new_n683), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n519), .B1(new_n679), .B2(new_n683), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n688), .B2(new_n686), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT110), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n689), .A2(new_n691), .A3(new_n692), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1325gat));
  AOI21_X1  g496(.A(G15gat), .B1(new_n679), .B2(new_n443), .ZN(new_n698));
  INV_X1    g497(.A(new_n448), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n679), .A2(G15gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(G1326gat));
  NAND2_X1  g500(.A1(new_n402), .A2(new_n406), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n679), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  INV_X1    g505(.A(new_n650), .ZN(new_n707));
  INV_X1    g506(.A(new_n678), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n608), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n512), .A2(new_n605), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(G29gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n472), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n713), .A2(KEYINPUT45), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT45), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n605), .B1(new_n496), .B2(new_n511), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT91), .B1(new_n501), .B2(new_n504), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n507), .A2(new_n506), .A3(new_n503), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n407), .A2(new_n448), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n494), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT112), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n731), .A3(new_n605), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n720), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n730), .A2(new_n718), .A3(new_n731), .A4(new_n605), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n709), .ZN(new_n736));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736), .B2(new_n500), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n737), .ZN(G1328gat));
  INV_X1    g537(.A(new_n710), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(G36gat), .A3(new_n497), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n736), .B2(new_n497), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1329gat));
  INV_X1    g542(.A(G43gat), .ZN(new_n744));
  INV_X1    g543(.A(new_n443), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n735), .A2(G43gat), .A3(new_n709), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(new_n448), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n750), .B(new_n746), .C1(new_n747), .C2(new_n448), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1330gat));
  OAI21_X1  g551(.A(G50gat), .B1(new_n736), .B2(new_n493), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n710), .A2(KEYINPUT114), .ZN(new_n754));
  INV_X1    g553(.A(G50gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(new_n703), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n710), .A2(KEYINPUT114), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n753), .A2(KEYINPUT48), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n735), .A2(new_n703), .A3(new_n709), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n758), .B1(new_n761), .B2(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(KEYINPUT48), .B2(new_n762), .ZN(G1331gat));
  AND3_X1   g562(.A1(new_n730), .A2(new_n612), .A3(new_n708), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n707), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n472), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n497), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  NAND3_X1  g572(.A1(new_n766), .A2(G71gat), .A3(new_n699), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n443), .B(KEYINPUT115), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n776), .B2(G71gat), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n765), .A2(new_n702), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT116), .B(G78gat), .Z(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1335gat));
  NOR2_X1   g580(.A1(new_n608), .A2(new_n678), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n730), .A2(new_n605), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n783), .A2(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n650), .ZN(new_n787));
  AOI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n472), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n608), .A2(new_n650), .A3(new_n678), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n735), .A2(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n790), .A2(new_n563), .A3(new_n500), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n788), .A2(new_n791), .ZN(G1336gat));
  NAND3_X1  g591(.A1(new_n735), .A2(new_n683), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G92gat), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n497), .A2(G92gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n783), .A2(new_n799), .A3(KEYINPUT51), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT51), .B1(new_n783), .B2(new_n799), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n800), .A2(new_n801), .A3(new_n650), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n793), .A2(G92gat), .B1(new_n802), .B2(new_n795), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n797), .B2(new_n803), .ZN(G1337gat));
  OAI21_X1  g603(.A(KEYINPUT118), .B1(new_n790), .B2(new_n448), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n735), .A2(new_n806), .A3(new_n699), .A4(new_n789), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(G99gat), .A3(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n650), .A2(new_n745), .A3(G99gat), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT119), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n786), .B2(new_n810), .ZN(G1338gat));
  NAND4_X1  g610(.A1(new_n733), .A2(new_n492), .A3(new_n734), .A4(new_n789), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G106gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n493), .A2(G106gat), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n784), .A2(new_n707), .A3(new_n785), .A4(new_n815), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n733), .A2(new_n703), .A3(new_n734), .A4(new_n789), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G106gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n783), .A2(new_n799), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n783), .A2(new_n799), .A3(KEYINPUT51), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n822), .A2(new_n707), .A3(new_n823), .A4(new_n815), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n814), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT120), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n802), .A2(new_n815), .B1(G106gat), .B2(new_n818), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n814), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(G1339gat));
  NAND4_X1  g630(.A1(new_n606), .A2(new_n611), .A3(new_n650), .A4(new_n708), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n618), .B(new_n635), .C1(new_n640), .C2(KEYINPUT10), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n616), .B1(new_n647), .B2(KEYINPUT54), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n616), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n647), .A2(new_n641), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n636), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n834), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n662), .B1(new_n660), .B2(new_n663), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n652), .B1(new_n651), .B2(new_n654), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n670), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n675), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n609), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n837), .A2(new_n678), .A3(new_n843), .A4(new_n839), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n644), .B2(new_n649), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n605), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n554), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n832), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n500), .A2(new_n683), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n509), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n302), .A3(new_n678), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n443), .A3(new_n702), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n708), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1340gat));
  OAI21_X1  g661(.A(G120gat), .B1(new_n860), .B2(new_n650), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n650), .B1(new_n304), .B2(new_n306), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1341gat));
  AOI21_X1  g665(.A(G127gat), .B1(new_n858), .B2(new_n608), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n860), .A2(new_n554), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(G127gat), .B2(new_n868), .ZN(G1342gat));
  INV_X1    g668(.A(G134gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n858), .A2(new_n870), .A3(new_n605), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT56), .Z(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n860), .B2(new_n609), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(new_n330), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n448), .A2(new_n856), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n851), .A2(new_n852), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n609), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT121), .B(new_n605), .C1(new_n851), .C2(new_n852), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n850), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n608), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n832), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT57), .B(new_n703), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n855), .A2(new_n492), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n876), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n875), .B1(new_n889), .B2(new_n678), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n886), .A2(new_n876), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n315), .A3(new_n678), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT122), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  AOI211_X1 g694(.A(new_n708), .B(new_n876), .C1(new_n885), .C2(new_n888), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n895), .B(new_n892), .C1(new_n896), .C2(new_n875), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n894), .A2(KEYINPUT58), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT58), .B1(new_n894), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1344gat));
  NAND3_X1  g699(.A1(new_n891), .A2(new_n317), .A3(new_n707), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT123), .Z(new_n902));
  XNOR2_X1  g701(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n832), .B2(new_n854), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n886), .A2(KEYINPUT57), .B1(new_n904), .B2(new_n703), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n707), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n876), .A2(KEYINPUT125), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n876), .A2(KEYINPUT125), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT59), .B(new_n317), .C1(new_n889), .C2(new_n707), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n902), .B1(new_n910), .B2(new_n911), .ZN(G1345gat));
  AOI21_X1  g711(.A(G155gat), .B1(new_n891), .B2(new_n608), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n608), .A2(G155gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n889), .B2(new_n914), .ZN(G1346gat));
  AOI21_X1  g714(.A(G162gat), .B1(new_n891), .B2(new_n605), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n889), .A2(new_n605), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n472), .A2(new_n497), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n855), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n509), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n213), .A3(new_n678), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n702), .A3(new_n775), .ZN(new_n924));
  OAI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n708), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1348gat));
  AOI21_X1  g725(.A(G176gat), .B1(new_n922), .B2(new_n707), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n924), .A2(new_n214), .A3(new_n650), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  OAI21_X1  g728(.A(G183gat), .B1(new_n924), .B2(new_n554), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n608), .B1(new_n205), .B2(new_n204), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n921), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n922), .A2(new_n203), .A3(new_n605), .ZN(new_n934));
  OAI21_X1  g733(.A(G190gat), .B1(new_n924), .B2(new_n609), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT126), .ZN(G1351gat));
  NAND2_X1  g738(.A1(new_n448), .A2(new_n919), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n905), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n708), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n886), .A2(new_n940), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n260), .A3(new_n678), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1352gat));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n263), .A3(new_n707), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n263), .B1(new_n906), .B2(new_n941), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n948), .A2(new_n949), .ZN(G1353gat));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n951), .B1(new_n942), .B2(new_n554), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n905), .A2(KEYINPUT127), .A3(new_n608), .A4(new_n941), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(G211gat), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n944), .A2(new_n267), .A3(new_n608), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n942), .B2(new_n609), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n268), .A3(new_n605), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1355gat));
endmodule


