

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U549 ( .A1(n922), .A2(n702), .ZN(n712) );
  NAND2_X1 U550 ( .A1(n692), .A2(n691), .ZN(n737) );
  NOR2_X1 U551 ( .A1(G164), .A2(G1384), .ZN(n691) );
  XOR2_X1 U552 ( .A(KEYINPUT81), .B(n557), .Z(n514) );
  AND2_X1 U553 ( .A1(n752), .A2(n751), .ZN(n515) );
  NAND2_X1 U554 ( .A1(n761), .A2(n760), .ZN(n516) );
  AND2_X1 U555 ( .A1(n707), .A2(G1996), .ZN(n699) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U557 ( .A(n723), .B(n722), .ZN(n728) );
  NOR2_X1 U558 ( .A1(n753), .A2(n515), .ZN(n754) );
  INV_X1 U559 ( .A(n923), .ZN(n765) );
  INV_X1 U560 ( .A(KEYINPUT93), .ZN(n777) );
  XNOR2_X1 U561 ( .A(n778), .B(n777), .ZN(n779) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XNOR2_X1 U563 ( .A(n517), .B(KEYINPUT65), .ZN(n852) );
  NOR2_X1 U564 ( .A1(n650), .A2(G651), .ZN(n644) );
  NOR2_X1 U565 ( .A1(n527), .A2(n526), .ZN(G160) );
  NAND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NAND2_X1 U567 ( .A1(n852), .A2(G113), .ZN(n520) );
  INV_X1 U568 ( .A(G2105), .ZN(n523) );
  AND2_X1 U569 ( .A1(n523), .A2(G2104), .ZN(n857) );
  NAND2_X1 U570 ( .A1(G101), .A2(n857), .ZN(n518) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U572 ( .A1(n520), .A2(n519), .ZN(n527) );
  XOR2_X1 U573 ( .A(KEYINPUT66), .B(n521), .Z(n522) );
  XNOR2_X1 U574 ( .A(KEYINPUT17), .B(n522), .ZN(n849) );
  NAND2_X1 U575 ( .A1(G137), .A2(n849), .ZN(n525) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n523), .ZN(n851) );
  NAND2_X1 U577 ( .A1(n851), .A2(G125), .ZN(n524) );
  NAND2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  INV_X1 U580 ( .A(G651), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n650), .A2(n531), .ZN(n636) );
  NAND2_X1 U582 ( .A1(n636), .A2(G72), .ZN(n530) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n528) );
  XNOR2_X1 U584 ( .A(n528), .B(KEYINPUT64), .ZN(n637) );
  NAND2_X1 U585 ( .A1(G85), .A2(n637), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U587 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n532), .Z(n649) );
  NAND2_X1 U589 ( .A1(G60), .A2(n649), .ZN(n534) );
  NAND2_X1 U590 ( .A1(G47), .A2(n644), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n535) );
  OR2_X1 U592 ( .A1(n536), .A2(n535), .ZN(G290) );
  XOR2_X1 U593 ( .A(G2451), .B(G2454), .Z(n538) );
  XNOR2_X1 U594 ( .A(G2430), .B(KEYINPUT96), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U596 ( .A(n539), .B(G2446), .Z(n541) );
  XNOR2_X1 U597 ( .A(G1341), .B(G1348), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n541), .B(n540), .ZN(n545) );
  XOR2_X1 U599 ( .A(G2438), .B(G2427), .Z(n543) );
  XNOR2_X1 U600 ( .A(G2443), .B(G2435), .ZN(n542) );
  XNOR2_X1 U601 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U602 ( .A(n545), .B(n544), .Z(n546) );
  AND2_X1 U603 ( .A1(G14), .A2(n546), .ZN(G401) );
  NAND2_X1 U604 ( .A1(G64), .A2(n649), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G52), .A2(n644), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n636), .A2(G77), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G90), .A2(n637), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(n551), .ZN(n552) );
  XNOR2_X1 U611 ( .A(KEYINPUT67), .B(n552), .ZN(n553) );
  NOR2_X1 U612 ( .A1(n554), .A2(n553), .ZN(G171) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(G102), .A2(n857), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G138), .A2(n849), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n852), .A2(G114), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n851), .A2(G126), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n514), .A2(n558), .ZN(n559) );
  NOR2_X1 U620 ( .A1(n560), .A2(n559), .ZN(G164) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U623 ( .A(KEYINPUT70), .B(KEYINPUT6), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G63), .A2(n649), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G51), .A2(n644), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n564), .B(n563), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G89), .A2(n637), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G76), .A2(n636), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT69), .B(n568), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT5), .B(n569), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT7), .B(n572), .Z(G168) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U639 ( .A(G223), .ZN(n821) );
  NAND2_X1 U640 ( .A1(n821), .A2(G567), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U642 ( .A1(G56), .A2(n649), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n575), .Z(n581) );
  NAND2_X1 U644 ( .A1(G81), .A2(n637), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G68), .A2(n636), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n579), .Z(n580) );
  NOR2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n644), .A2(G43), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n922) );
  INV_X1 U652 ( .A(G860), .ZN(n602) );
  OR2_X1 U653 ( .A1(n922), .A2(n602), .ZN(G153) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G66), .A2(n649), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G92), .A2(n637), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G79), .A2(n636), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G54), .A2(n644), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n590), .Z(n909) );
  OR2_X1 U664 ( .A1(n909), .A2(G868), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G65), .A2(n649), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G53), .A2(n644), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n636), .A2(G78), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G91), .A2(n637), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n906) );
  INV_X1 U673 ( .A(n906), .ZN(G299) );
  XNOR2_X1 U674 ( .A(KEYINPUT71), .B(G868), .ZN(n599) );
  NOR2_X1 U675 ( .A1(G286), .A2(n599), .ZN(n601) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U677 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n603), .A2(n909), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n922), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n909), .A2(G868), .ZN(n605) );
  NOR2_X1 U683 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(G282) );
  XOR2_X1 U685 ( .A(KEYINPUT72), .B(KEYINPUT18), .Z(n609) );
  NAND2_X1 U686 ( .A1(G123), .A2(n851), .ZN(n608) );
  XNOR2_X1 U687 ( .A(n609), .B(n608), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G99), .A2(n857), .ZN(n611) );
  NAND2_X1 U689 ( .A1(G111), .A2(n852), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n612), .B(KEYINPUT73), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G135), .A2(n849), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n984) );
  XNOR2_X1 U695 ( .A(G2096), .B(n984), .ZN(n618) );
  INV_X1 U696 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G559), .A2(n909), .ZN(n619) );
  XNOR2_X1 U699 ( .A(n922), .B(n619), .ZN(n660) );
  NOR2_X1 U700 ( .A1(n660), .A2(G860), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n636), .A2(G80), .ZN(n621) );
  NAND2_X1 U702 ( .A1(G93), .A2(n637), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n649), .A2(G67), .ZN(n622) );
  XNOR2_X1 U705 ( .A(n622), .B(KEYINPUT74), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G55), .A2(n644), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U708 ( .A(KEYINPUT75), .B(n625), .Z(n626) );
  NOR2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n656) );
  XNOR2_X1 U710 ( .A(n628), .B(n656), .ZN(G145) );
  NAND2_X1 U711 ( .A1(G61), .A2(n649), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G86), .A2(n637), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n636), .A2(G73), .ZN(n631) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n631), .Z(n632) );
  NOR2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n644), .A2(G48), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U719 ( .A1(n636), .A2(G75), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G88), .A2(n637), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G62), .A2(n649), .ZN(n641) );
  NAND2_X1 U723 ( .A1(G50), .A2(n644), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U725 ( .A1(n643), .A2(n642), .ZN(G166) );
  INV_X1 U726 ( .A(G166), .ZN(G303) );
  NAND2_X1 U727 ( .A1(G49), .A2(n644), .ZN(n646) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U730 ( .A(KEYINPUT76), .B(n647), .ZN(n648) );
  NOR2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n650), .A2(G87), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(G288) );
  NOR2_X1 U734 ( .A1(G868), .A2(n656), .ZN(n653) );
  XNOR2_X1 U735 ( .A(n653), .B(KEYINPUT77), .ZN(n663) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(G305), .ZN(n654) );
  XNOR2_X1 U737 ( .A(n654), .B(G303), .ZN(n655) );
  XNOR2_X1 U738 ( .A(n656), .B(n655), .ZN(n658) );
  XNOR2_X1 U739 ( .A(G290), .B(n906), .ZN(n657) );
  XNOR2_X1 U740 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U741 ( .A(n659), .B(G288), .ZN(n871) );
  XOR2_X1 U742 ( .A(n871), .B(n660), .Z(n661) );
  NAND2_X1 U743 ( .A1(G868), .A2(n661), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U747 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n666), .B(KEYINPUT78), .ZN(n667) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U750 ( .A1(G2072), .A2(n668), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U752 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  NOR2_X1 U753 ( .A1(G219), .A2(G220), .ZN(n669) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U755 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U756 ( .A1(G96), .A2(n671), .ZN(n825) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n825), .ZN(n675) );
  NAND2_X1 U758 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U759 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G108), .A2(n673), .ZN(n826) );
  NAND2_X1 U761 ( .A1(G567), .A2(n826), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U763 ( .A(KEYINPUT79), .B(n676), .ZN(G319) );
  INV_X1 U764 ( .A(G319), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n677) );
  XNOR2_X1 U766 ( .A(KEYINPUT80), .B(n677), .ZN(n678) );
  NOR2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n824) );
  NAND2_X1 U768 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n690) );
  NOR2_X1 U770 ( .A1(n690), .A2(n691), .ZN(n816) );
  XNOR2_X1 U771 ( .A(G2067), .B(KEYINPUT37), .ZN(n814) );
  NAND2_X1 U772 ( .A1(G104), .A2(n857), .ZN(n682) );
  NAND2_X1 U773 ( .A1(G140), .A2(n849), .ZN(n681) );
  NAND2_X1 U774 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U775 ( .A(KEYINPUT34), .B(n683), .ZN(n688) );
  NAND2_X1 U776 ( .A1(G128), .A2(n851), .ZN(n685) );
  NAND2_X1 U777 ( .A1(G116), .A2(n852), .ZN(n684) );
  NAND2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U779 ( .A(KEYINPUT35), .B(n686), .Z(n687) );
  NOR2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U781 ( .A(KEYINPUT36), .B(n689), .ZN(n846) );
  NOR2_X1 U782 ( .A1(n814), .A2(n846), .ZN(n989) );
  NAND2_X1 U783 ( .A1(n816), .A2(n989), .ZN(n811) );
  INV_X1 U784 ( .A(n811), .ZN(n782) );
  INV_X1 U785 ( .A(n690), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n737), .A2(G8), .ZN(n693) );
  XNOR2_X2 U787 ( .A(n693), .B(KEYINPUT86), .ZN(n774) );
  NOR2_X1 U788 ( .A1(G1981), .A2(G305), .ZN(n694) );
  XOR2_X1 U789 ( .A(n694), .B(KEYINPUT24), .Z(n695) );
  NOR2_X1 U790 ( .A1(n774), .A2(n695), .ZN(n780) );
  INV_X1 U791 ( .A(n737), .ZN(n707) );
  NOR2_X1 U792 ( .A1(n707), .A2(G1348), .ZN(n697) );
  NOR2_X1 U793 ( .A1(G2067), .A2(n737), .ZN(n696) );
  NOR2_X1 U794 ( .A1(n697), .A2(n696), .ZN(n704) );
  XNOR2_X1 U795 ( .A(KEYINPUT26), .B(KEYINPUT89), .ZN(n698) );
  XNOR2_X1 U796 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n737), .A2(G1341), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n909), .A2(n712), .ZN(n703) );
  NAND2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U801 ( .A(n705), .B(KEYINPUT90), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n707), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U803 ( .A(n706), .B(KEYINPUT27), .ZN(n709) );
  INV_X1 U804 ( .A(G1956), .ZN(n934) );
  NOR2_X1 U805 ( .A1(n934), .A2(n707), .ZN(n708) );
  NOR2_X1 U806 ( .A1(n709), .A2(n708), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n717), .A2(n906), .ZN(n711) );
  XOR2_X1 U808 ( .A(KEYINPUT28), .B(KEYINPUT88), .Z(n710) );
  XNOR2_X1 U809 ( .A(n711), .B(n710), .ZN(n716) );
  OR2_X1 U810 ( .A1(n712), .A2(n909), .ZN(n713) );
  AND2_X1 U811 ( .A1(n716), .A2(n713), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n721) );
  INV_X1 U813 ( .A(n716), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n717), .A2(n906), .ZN(n718) );
  OR2_X1 U815 ( .A1(n719), .A2(n718), .ZN(n720) );
  AND2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n723) );
  XOR2_X1 U817 ( .A(G2078), .B(KEYINPUT25), .Z(n724) );
  XNOR2_X1 U818 ( .A(KEYINPUT87), .B(n724), .ZN(n969) );
  NOR2_X1 U819 ( .A1(n737), .A2(n969), .ZN(n726) );
  AND2_X1 U820 ( .A1(n737), .A2(G1961), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n732) );
  NAND2_X1 U822 ( .A1(G171), .A2(n732), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n728), .A2(n727), .ZN(n751) );
  NOR2_X1 U824 ( .A1(n774), .A2(G1966), .ZN(n753) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n737), .ZN(n750) );
  NOR2_X1 U826 ( .A1(n753), .A2(n750), .ZN(n729) );
  NAND2_X1 U827 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U828 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U829 ( .A1(G168), .A2(n731), .ZN(n734) );
  NOR2_X1 U830 ( .A1(G171), .A2(n732), .ZN(n733) );
  NOR2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n736) );
  XNOR2_X1 U832 ( .A(KEYINPUT91), .B(KEYINPUT31), .ZN(n735) );
  XNOR2_X1 U833 ( .A(n736), .B(n735), .ZN(n752) );
  INV_X1 U834 ( .A(G8), .ZN(n742) );
  NOR2_X1 U835 ( .A1(n774), .A2(G1971), .ZN(n739) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n737), .ZN(n738) );
  NOR2_X1 U837 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U838 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n744) );
  AND2_X1 U840 ( .A1(n752), .A2(n744), .ZN(n743) );
  NAND2_X1 U841 ( .A1(n751), .A2(n743), .ZN(n748) );
  INV_X1 U842 ( .A(n744), .ZN(n746) );
  AND2_X1 U843 ( .A1(G286), .A2(G8), .ZN(n745) );
  OR2_X1 U844 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U845 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U846 ( .A(n749), .B(KEYINPUT32), .ZN(n757) );
  NAND2_X1 U847 ( .A1(G8), .A2(n750), .ZN(n755) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n771) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U852 ( .A1(n763), .A2(n758), .ZN(n916) );
  NAND2_X1 U853 ( .A1(n771), .A2(n916), .ZN(n761) );
  INV_X1 U854 ( .A(n774), .ZN(n759) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n915) );
  AND2_X1 U856 ( .A1(n759), .A2(n915), .ZN(n760) );
  INV_X1 U857 ( .A(KEYINPUT33), .ZN(n762) );
  NAND2_X1 U858 ( .A1(n516), .A2(n762), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n763), .A2(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U860 ( .A1(n774), .A2(n764), .ZN(n766) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n923) );
  NOR2_X1 U862 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n776) );
  NOR2_X1 U864 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U865 ( .A1(G8), .A2(n769), .ZN(n770) );
  XNOR2_X1 U866 ( .A(n770), .B(KEYINPUT92), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U868 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n778) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n804) );
  NAND2_X1 U872 ( .A1(G95), .A2(n857), .ZN(n784) );
  NAND2_X1 U873 ( .A1(G131), .A2(n849), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U875 ( .A(KEYINPUT82), .B(n785), .Z(n789) );
  NAND2_X1 U876 ( .A1(G119), .A2(n851), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G107), .A2(n852), .ZN(n786) );
  AND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n864) );
  NAND2_X1 U880 ( .A1(G1991), .A2(n864), .ZN(n790) );
  XNOR2_X1 U881 ( .A(n790), .B(KEYINPUT83), .ZN(n801) );
  NAND2_X1 U882 ( .A1(n849), .A2(G141), .ZN(n791) );
  XNOR2_X1 U883 ( .A(n791), .B(KEYINPUT84), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G129), .A2(n851), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G117), .A2(n852), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n857), .A2(G105), .ZN(n794) );
  XOR2_X1 U888 ( .A(KEYINPUT38), .B(n794), .Z(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U891 ( .A(KEYINPUT85), .B(n799), .Z(n843) );
  AND2_X1 U892 ( .A1(G1996), .A2(n843), .ZN(n800) );
  NOR2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n991) );
  XOR2_X1 U894 ( .A(G1986), .B(G290), .Z(n907) );
  NAND2_X1 U895 ( .A1(n991), .A2(n907), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n802), .A2(n816), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n819) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n843), .ZN(n994) );
  INV_X1 U899 ( .A(n991), .ZN(n808) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n864), .A2(G1991), .ZN(n805) );
  XNOR2_X1 U902 ( .A(n805), .B(KEYINPUT94), .ZN(n983) );
  NOR2_X1 U903 ( .A1(n806), .A2(n983), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n994), .A2(n809), .ZN(n810) );
  XNOR2_X1 U906 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U908 ( .A(KEYINPUT95), .B(n813), .Z(n815) );
  NAND2_X1 U909 ( .A1(n814), .A2(n846), .ZN(n1006) );
  NAND2_X1 U910 ( .A1(n815), .A2(n1006), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U913 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U916 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(G188) );
  XNOR2_X1 U919 ( .A(G96), .B(KEYINPUT97), .ZN(G221) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G69), .ZN(G235) );
  NOR2_X1 U923 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  NAND2_X1 U925 ( .A1(G124), .A2(n851), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n827), .B(KEYINPUT44), .ZN(n834) );
  NAND2_X1 U927 ( .A1(G100), .A2(n857), .ZN(n829) );
  NAND2_X1 U928 ( .A1(G136), .A2(n849), .ZN(n828) );
  NAND2_X1 U929 ( .A1(n829), .A2(n828), .ZN(n832) );
  NAND2_X1 U930 ( .A1(G112), .A2(n852), .ZN(n830) );
  XNOR2_X1 U931 ( .A(KEYINPUT105), .B(n830), .ZN(n831) );
  NOR2_X1 U932 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U933 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U934 ( .A(KEYINPUT106), .B(n835), .Z(G162) );
  NAND2_X1 U935 ( .A1(G130), .A2(n851), .ZN(n837) );
  NAND2_X1 U936 ( .A1(G118), .A2(n852), .ZN(n836) );
  NAND2_X1 U937 ( .A1(n837), .A2(n836), .ZN(n842) );
  NAND2_X1 U938 ( .A1(G106), .A2(n857), .ZN(n839) );
  NAND2_X1 U939 ( .A1(G142), .A2(n849), .ZN(n838) );
  NAND2_X1 U940 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n840), .B(KEYINPUT45), .Z(n841) );
  NOR2_X1 U942 ( .A1(n842), .A2(n841), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U944 ( .A(G164), .B(n984), .Z(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n863) );
  NAND2_X1 U947 ( .A1(G139), .A2(n849), .ZN(n850) );
  XNOR2_X1 U948 ( .A(KEYINPUT107), .B(n850), .ZN(n861) );
  NAND2_X1 U949 ( .A1(G127), .A2(n851), .ZN(n854) );
  NAND2_X1 U950 ( .A1(G115), .A2(n852), .ZN(n853) );
  NAND2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n855), .B(KEYINPUT47), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n856), .B(KEYINPUT108), .ZN(n859) );
  NAND2_X1 U954 ( .A1(n857), .A2(G103), .ZN(n858) );
  NAND2_X1 U955 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U956 ( .A1(n861), .A2(n860), .ZN(n999) );
  XNOR2_X1 U957 ( .A(G162), .B(n999), .ZN(n862) );
  XNOR2_X1 U958 ( .A(n863), .B(n862), .ZN(n869) );
  XNOR2_X1 U959 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n866) );
  XNOR2_X1 U960 ( .A(n864), .B(KEYINPUT109), .ZN(n865) );
  XNOR2_X1 U961 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U962 ( .A(G160), .B(n867), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n869), .B(n868), .ZN(n870) );
  NOR2_X1 U964 ( .A1(G37), .A2(n870), .ZN(G395) );
  XOR2_X1 U965 ( .A(n871), .B(G286), .Z(n873) );
  XNOR2_X1 U966 ( .A(G171), .B(n909), .ZN(n872) );
  XNOR2_X1 U967 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U968 ( .A(n874), .B(n922), .Z(n875) );
  NOR2_X1 U969 ( .A1(G37), .A2(n875), .ZN(G397) );
  XOR2_X1 U970 ( .A(KEYINPUT101), .B(KEYINPUT104), .Z(n877) );
  XNOR2_X1 U971 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n876) );
  XNOR2_X1 U972 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U973 ( .A(n878), .B(KEYINPUT41), .Z(n880) );
  XNOR2_X1 U974 ( .A(G1971), .B(G1976), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n880), .B(n879), .ZN(n888) );
  XOR2_X1 U976 ( .A(G1956), .B(G1966), .Z(n882) );
  XNOR2_X1 U977 ( .A(G1986), .B(G1981), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(n886) );
  XOR2_X1 U979 ( .A(G2474), .B(G1961), .Z(n884) );
  XNOR2_X1 U980 ( .A(G1996), .B(G1991), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n886), .B(n885), .Z(n887) );
  XNOR2_X1 U983 ( .A(n888), .B(n887), .ZN(G229) );
  XOR2_X1 U984 ( .A(G2678), .B(KEYINPUT99), .Z(n890) );
  XNOR2_X1 U985 ( .A(KEYINPUT98), .B(G2096), .ZN(n889) );
  XNOR2_X1 U986 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U987 ( .A(n891), .B(KEYINPUT42), .Z(n893) );
  XNOR2_X1 U988 ( .A(G2078), .B(G2072), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U990 ( .A(G2100), .B(G2090), .Z(n895) );
  XNOR2_X1 U991 ( .A(G2067), .B(G2084), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U993 ( .A(n897), .B(n896), .Z(n899) );
  XNOR2_X1 U994 ( .A(KEYINPUT43), .B(KEYINPUT100), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(G227) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n900), .B(KEYINPUT110), .ZN(n901) );
  NAND2_X1 U998 ( .A1(G319), .A2(n901), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G401), .A2(n902), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n903) );
  XOR2_X1 U1001 ( .A(KEYINPUT49), .B(n903), .Z(n904) );
  NAND2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1005 ( .A(G16), .B(KEYINPUT56), .ZN(n932) );
  XNOR2_X1 U1006 ( .A(n906), .B(G1956), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(G171), .B(G1961), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n912) );
  XOR2_X1 U1009 ( .A(G1348), .B(n909), .Z(n910) );
  XNOR2_X1 U1010 ( .A(KEYINPUT120), .B(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n921) );
  AND2_X1 U1013 ( .A1(G303), .A2(G1971), .ZN(n918) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(KEYINPUT121), .B(n919), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n930) );
  XNOR2_X1 U1018 ( .A(n922), .B(G1341), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n924) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(KEYINPUT57), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT119), .B(n926), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n1016) );
  XOR2_X1 U1026 ( .A(G16), .B(KEYINPUT122), .Z(n960) );
  XNOR2_X1 U1027 ( .A(KEYINPUT127), .B(G1966), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(n933), .B(G21), .ZN(n950) );
  XNOR2_X1 U1029 ( .A(G1961), .B(G5), .ZN(n948) );
  XNOR2_X1 U1030 ( .A(n934), .B(G20), .ZN(n944) );
  XOR2_X1 U1031 ( .A(G1341), .B(G19), .Z(n939) );
  XOR2_X1 U1032 ( .A(KEYINPUT125), .B(G4), .Z(n936) );
  XNOR2_X1 U1033 ( .A(G1348), .B(KEYINPUT59), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(n936), .B(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT124), .B(n937), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n942) );
  XOR2_X1 U1037 ( .A(KEYINPUT123), .B(G1981), .Z(n940) );
  XNOR2_X1 U1038 ( .A(G6), .B(n940), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT126), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT60), .B(n946), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n957) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G22), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G23), .B(G1976), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n954) );
  XOR2_X1 U1048 ( .A(G1986), .B(G24), .Z(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT58), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(n958), .B(KEYINPUT61), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n961), .ZN(n1014) );
  XNOR2_X1 U1055 ( .A(G1996), .B(G32), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G33), .B(G2072), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n968) );
  XOR2_X1 U1058 ( .A(G1991), .B(G25), .Z(n964) );
  NAND2_X1 U1059 ( .A1(n964), .A2(G28), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G26), .B(G2067), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1063 ( .A(G27), .B(n969), .Z(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1065 ( .A(KEYINPUT53), .B(n972), .Z(n976) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(G34), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G2084), .B(n974), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G35), .B(G2090), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(KEYINPUT116), .B(n977), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(KEYINPUT118), .B(n980), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(G29), .A2(n981), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT55), .ZN(n1012) );
  XOR2_X1 U1076 ( .A(KEYINPUT115), .B(KEYINPUT52), .Z(n1009) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1078 ( .A(KEYINPUT111), .B(n985), .Z(n987) );
  XNOR2_X1 U1079 ( .A(G160), .B(G2084), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(KEYINPUT112), .B(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT113), .ZN(n998) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n995) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT51), .B(n996), .Z(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1005) );
  XOR2_X1 U1089 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(KEYINPUT114), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1009), .B(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(G29), .A2(n1010), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1017), .Z(G311) );
  INV_X1 U1102 ( .A(G311), .ZN(G150) );
endmodule

