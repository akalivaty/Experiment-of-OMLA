//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT83), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G122), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT2), .A2(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT68), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT2), .A3(G113), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n192), .A2(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G119), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G101), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n201), .A2(new_n204), .A3(new_n208), .A4(new_n205), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n211), .A3(G101), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n200), .A2(G107), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n203), .A2(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G116), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n219), .B(G113), .C1(KEYINPUT5), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n197), .A2(new_n198), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI211_X1 g038(.A(KEYINPUT6), .B(new_n190), .C1(new_n213), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  OR2_X1    g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G146), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G143), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n226), .B(new_n227), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n228), .B2(G146), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(KEYINPUT64), .A3(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(G146), .ZN(new_n236));
  INV_X1    g050(.A(new_n226), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n234), .A2(new_n235), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G125), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT82), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n238), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(G125), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n230), .A2(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n246), .A2(G128), .B1(new_n245), .B2(new_n236), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n234), .A2(new_n235), .A3(new_n250), .A4(new_n236), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n241), .B(new_n244), .C1(new_n254), .C2(G125), .ZN(new_n255));
  INV_X1    g069(.A(G224), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n235), .A2(new_n236), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n234), .A4(new_n250), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n247), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n240), .ZN(new_n264));
  INV_X1    g078(.A(new_n257), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n241), .A4(new_n244), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n197), .A2(new_n198), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n192), .A2(new_n194), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n195), .A2(new_n196), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n268), .A2(new_n269), .A3(new_n198), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n212), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n210), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n224), .B(new_n190), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT81), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n213), .A2(new_n275), .A3(new_n224), .A4(new_n190), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n190), .B1(new_n213), .B2(new_n224), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI221_X4 g094(.A(new_n225), .B1(new_n258), .B2(new_n266), .C1(new_n277), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n277), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n265), .A2(KEYINPUT7), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n255), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n284), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n264), .A2(new_n241), .A3(new_n244), .A4(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n190), .B(KEYINPUT8), .ZN(new_n288));
  INV_X1    g102(.A(new_n224), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n218), .B1(new_n223), .B2(new_n222), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n282), .B1(new_n283), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n189), .B1(new_n281), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n292), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n296), .B2(new_n277), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n277), .A2(new_n280), .ZN(new_n298));
  INV_X1    g112(.A(new_n225), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n258), .A2(new_n266), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n301), .A3(new_n188), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n294), .A2(new_n295), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(G110), .B(G140), .ZN(new_n304));
  INV_X1    g118(.A(G227), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G953), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n304), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n254), .A2(KEYINPUT69), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n263), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n217), .A2(new_n311), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G137), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT11), .B1(new_n314), .B2(G134), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(G134), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OR2_X1    g131(.A1(KEYINPUT65), .A2(G137), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT65), .A2(G137), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT11), .A2(G134), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n317), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n210), .A2(new_n239), .A3(new_n212), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n261), .A2(new_n262), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n259), .A2(new_n234), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n246), .A2(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n217), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n327), .B1(new_n332), .B2(KEYINPUT10), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n313), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n326), .ZN(new_n335));
  INV_X1    g149(.A(new_n327), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n328), .A2(new_n331), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n218), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n338), .B2(new_n311), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n307), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n328), .A2(new_n248), .A3(new_n217), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n326), .B1(new_n343), .B2(new_n332), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT12), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT12), .B(new_n326), .C1(new_n343), .C2(new_n332), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n339), .A2(new_n335), .A3(new_n340), .ZN(new_n349));
  INV_X1    g163(.A(new_n307), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n342), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G469), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n282), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n326), .B1(new_n313), .B2(new_n333), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n349), .A3(new_n350), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n313), .A2(new_n333), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n357), .A2(new_n335), .B1(new_n346), .B2(new_n347), .ZN(new_n358));
  OAI211_X1 g172(.A(G469), .B(new_n356), .C1(new_n358), .C2(new_n350), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n353), .A2(new_n282), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n354), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT9), .B(G234), .ZN(new_n363));
  OAI21_X1  g177(.A(G221), .B1(new_n363), .B2(G902), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n364), .B(KEYINPUT80), .Z(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n303), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT16), .ZN(new_n369));
  INV_X1    g183(.A(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n240), .A2(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n371), .B1(new_n374), .B2(new_n369), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n230), .ZN(new_n376));
  NOR2_X1   g190(.A1(G237), .A2(G953), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(G143), .A3(G214), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(G143), .B1(new_n377), .B2(G214), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT17), .B(G131), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(G146), .B(new_n371), .C1(new_n374), .C2(new_n369), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  INV_X1    g200(.A(G953), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n228), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n378), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT85), .B1(new_n390), .B2(G131), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(G131), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n389), .A2(new_n394), .A3(new_n324), .A4(new_n378), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n376), .A2(new_n381), .A3(KEYINPUT87), .A4(new_n382), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n385), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n379), .A2(new_n380), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT18), .A2(G131), .ZN(new_n400));
  XNOR2_X1  g214(.A(G125), .B(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n230), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n374), .A2(G146), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n399), .A2(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n405));
  INV_X1    g219(.A(new_n400), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(new_n390), .B2(new_n406), .ZN(new_n407));
  AOI211_X1 g221(.A(KEYINPUT84), .B(new_n400), .C1(new_n389), .C2(new_n378), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(G113), .B(G122), .Z(new_n410));
  XOR2_X1   g224(.A(KEYINPUT86), .B(G104), .Z(new_n411));
  XOR2_X1   g225(.A(new_n410), .B(new_n411), .Z(new_n412));
  NAND3_X1  g226(.A1(new_n398), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n391), .A2(new_n393), .A3(new_n395), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n382), .A2(KEYINPUT78), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n401), .A2(KEYINPUT16), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT78), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(G146), .A4(new_n371), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n374), .B(KEYINPUT19), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n415), .B(new_n418), .C1(new_n419), .C2(G146), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n409), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n412), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(G475), .A2(G902), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n368), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n425), .ZN(new_n427));
  AOI211_X1 g241(.A(KEYINPUT20), .B(new_n427), .C1(new_n413), .C2(new_n423), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n398), .A2(new_n409), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n422), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n430), .B2(new_n413), .ZN(new_n431));
  INV_X1    g245(.A(G475), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n426), .A2(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n282), .B(new_n387), .C1(G234), .C2(G237), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G898), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n387), .A2(G952), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(G234), .B2(G237), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT95), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n433), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G128), .B(G143), .ZN(new_n444));
  INV_X1    g258(.A(G134), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G122), .ZN(new_n447));
  OR3_X1    g261(.A1(new_n447), .A2(KEYINPUT14), .A3(G116), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n447), .B2(G116), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n451));
  INV_X1    g265(.A(G116), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n451), .B1(new_n452), .B2(G122), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n447), .A2(KEYINPUT88), .A3(G116), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G107), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n453), .A2(new_n454), .B1(new_n452), .B2(G122), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n457), .A2(KEYINPUT90), .A3(new_n203), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT90), .B1(new_n457), .B2(new_n203), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n446), .B(new_n456), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G217), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n363), .A2(new_n461), .A3(G953), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT91), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n444), .A2(KEYINPUT89), .A3(new_n445), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n249), .A2(G143), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT13), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n445), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n228), .A2(G128), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n249), .A2(G143), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n445), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n465), .A2(new_n468), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n457), .A2(new_n203), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n457), .A2(new_n203), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n464), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n460), .A2(new_n463), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n463), .B1(new_n460), .B2(new_n476), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT93), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n480), .A2(new_n481), .A3(new_n282), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n460), .A2(new_n476), .ZN(new_n486));
  INV_X1    g300(.A(new_n463), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n488), .A2(new_n282), .A3(new_n484), .A4(new_n477), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT93), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n282), .A3(new_n477), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT92), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n488), .A2(new_n494), .A3(new_n282), .A4(new_n477), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n483), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n497), .B1(new_n491), .B2(new_n496), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n443), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n367), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n317), .A2(new_n321), .A3(new_n324), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n324), .B1(new_n317), .B2(new_n321), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n238), .B(new_n232), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n309), .B1(new_n328), .B2(new_n248), .ZN(new_n507));
  AOI211_X1 g321(.A(KEYINPUT69), .B(new_n247), .C1(new_n261), .C2(new_n262), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(G134), .B1(new_n318), .B2(new_n319), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n445), .B2(G137), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n314), .A2(KEYINPUT66), .A3(G134), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n325), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n506), .B1(new_n509), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n199), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT28), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n308), .A2(new_n310), .A3(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n505), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n199), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n519), .A3(new_n505), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n520), .B1(new_n525), .B2(KEYINPUT28), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(G101), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n377), .A2(G210), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n534), .A3(new_n532), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n538), .A2(KEYINPUT29), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n526), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n254), .A2(new_n517), .B1(new_n326), .B2(new_n239), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n519), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n505), .B1(new_n263), .B2(new_n516), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(KEYINPUT72), .A3(new_n199), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n524), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT28), .ZN(new_n547));
  INV_X1    g361(.A(new_n520), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n538), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n521), .A2(KEYINPUT30), .A3(new_n505), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n519), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n524), .ZN(new_n554));
  INV_X1    g368(.A(new_n538), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT29), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n540), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G472), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n547), .A2(new_n548), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n199), .B1(new_n542), .B2(KEYINPUT30), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n518), .B2(KEYINPUT30), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n524), .A2(new_n538), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n553), .A2(KEYINPUT31), .A3(new_n524), .A4(new_n538), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n561), .A2(new_n555), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(G472), .A2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n560), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n560), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT73), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n566), .A2(new_n567), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT28), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n544), .A2(KEYINPUT72), .A3(new_n199), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT72), .B1(new_n544), .B2(new_n199), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n579), .B2(new_n524), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n555), .B1(new_n580), .B2(new_n520), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n572), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n559), .A2(new_n571), .A3(new_n574), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n461), .B1(G234), .B2(new_n282), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n387), .A2(G221), .A3(G234), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n415), .A2(new_n418), .A3(new_n402), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT74), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n220), .B2(G128), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n249), .A2(KEYINPUT74), .A3(G119), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n249), .B2(G119), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n220), .A2(KEYINPUT75), .A3(G128), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT24), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(G110), .ZN(new_n602));
  INV_X1    g416(.A(G110), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT24), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT76), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(KEYINPUT24), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n601), .A2(G110), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT76), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n596), .A2(new_n600), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT23), .B1(new_n249), .B2(G119), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n249), .A2(G119), .ZN(new_n612));
  AND2_X1   g426(.A1(KEYINPUT23), .A2(G119), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n611), .A2(new_n612), .B1(new_n249), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n603), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT77), .B1(new_n610), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n600), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n608), .B1(new_n606), .B2(new_n607), .ZN(new_n620));
  OAI22_X1  g434(.A1(new_n618), .A2(new_n595), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT77), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n615), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n591), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n605), .A2(new_n609), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n600), .A2(new_n593), .A3(new_n594), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n376), .A2(new_n382), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n614), .A2(new_n603), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n624), .A2(KEYINPUT79), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT79), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n415), .A2(new_n418), .A3(new_n402), .ZN(new_n633));
  AOI221_X4 g447(.A(KEYINPUT77), .B1(new_n614), .B2(new_n603), .C1(new_n625), .C2(new_n626), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n622), .B1(new_n621), .B2(new_n615), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n590), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n590), .B1(new_n636), .B2(new_n637), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT25), .B1(new_n642), .B2(new_n282), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT79), .B1(new_n624), .B2(new_n630), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n636), .A2(new_n632), .A3(new_n637), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n589), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(KEYINPUT25), .B(new_n282), .C1(new_n646), .C2(new_n640), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n586), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n586), .A2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n502), .A2(new_n585), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G101), .ZN(G3));
  NAND4_X1  g469(.A1(new_n362), .A2(new_n649), .A3(new_n651), .A4(new_n366), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n575), .B2(new_n581), .ZN(new_n658));
  INV_X1    g472(.A(G472), .ZN(new_n659));
  OAI22_X1  g473(.A1(new_n658), .A2(new_n659), .B1(new_n568), .B2(new_n570), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n294), .A2(new_n302), .A3(new_n295), .A4(new_n441), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT33), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n463), .B2(KEYINPUT96), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n488), .A2(new_n477), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n665), .B1(new_n488), .B2(new_n477), .ZN(new_n667));
  OAI211_X1 g481(.A(G478), .B(new_n282), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n493), .A2(new_n482), .A3(new_n495), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n433), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT97), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT97), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n663), .B2(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n662), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT34), .B(G104), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G6));
  NOR2_X1   g493(.A1(new_n431), .A2(new_n432), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n424), .A2(new_n368), .A3(new_n425), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT98), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n681), .B1(new_n426), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n424), .A2(KEYINPUT98), .A3(new_n368), .A4(new_n425), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n491), .A2(new_n496), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT94), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n685), .A2(new_n687), .A3(new_n498), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n663), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n657), .A2(new_n661), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  OAI22_X1  g506(.A1(new_n631), .A2(new_n638), .B1(KEYINPUT36), .B2(new_n590), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n644), .A2(new_n645), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n650), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT25), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n646), .A2(new_n640), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n699), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n647), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n698), .B1(new_n702), .B2(new_n586), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n367), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n660), .A2(new_n501), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT37), .B(G110), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G12));
  INV_X1    g522(.A(G900), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT99), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(KEYINPUT99), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n434), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n439), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n685), .A2(new_n687), .A3(new_n498), .A4(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n704), .A2(new_n585), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  NAND2_X1  g531(.A1(new_n649), .A2(new_n697), .ZN(new_n718));
  INV_X1    g532(.A(new_n295), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n687), .A2(new_n498), .A3(new_n433), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n713), .B(KEYINPUT39), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n362), .A2(new_n366), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n294), .A2(new_n302), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT38), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n282), .B1(new_n525), .B2(new_n538), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n555), .B1(new_n553), .B2(new_n524), .ZN(new_n729));
  OAI21_X1  g543(.A(G472), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n571), .A2(new_n574), .A3(new_n584), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n721), .A2(new_n724), .A3(new_n727), .A4(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n228), .ZN(G45));
  AND3_X1   g549(.A1(new_n433), .A2(new_n670), .A3(new_n713), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n704), .A2(new_n585), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G146), .ZN(G48));
  INV_X1    g552(.A(new_n676), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n583), .B1(new_n582), .B2(new_n572), .ZN(new_n740));
  AOI211_X1 g554(.A(KEYINPUT73), .B(new_n573), .C1(new_n575), .C2(new_n581), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT32), .B1(new_n582), .B2(new_n569), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n659), .B1(new_n540), .B2(new_n557), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n652), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT100), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n352), .A2(new_n282), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(G469), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n354), .ZN(new_n750));
  INV_X1    g564(.A(new_n364), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n739), .A2(new_n746), .A3(new_n747), .A4(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n585), .A2(new_n653), .A3(new_n752), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT100), .B1(new_n754), .B2(new_n676), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT41), .B(G113), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G15));
  NAND4_X1  g572(.A1(new_n585), .A2(new_n653), .A3(new_n689), .A4(new_n752), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  NAND3_X1  g574(.A1(new_n294), .A2(new_n302), .A3(new_n295), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n750), .A2(new_n751), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n703), .A2(new_n501), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n585), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G119), .ZN(G21));
  INV_X1    g579(.A(new_n658), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n575), .B1(new_n538), .B2(new_n526), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n766), .A2(G472), .B1(new_n569), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n353), .B1(new_n352), .B2(new_n282), .ZN(new_n769));
  AOI211_X1 g583(.A(G469), .B(G902), .C1(new_n342), .C2(new_n351), .ZN(new_n770));
  NOR4_X1   g584(.A1(new_n769), .A2(new_n770), .A3(new_n751), .A4(new_n442), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n720), .A2(new_n761), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n768), .A2(new_n771), .A3(new_n653), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  OAI21_X1  g588(.A(G472), .B1(new_n568), .B2(G902), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n767), .A2(new_n569), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n718), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n769), .A2(new_n770), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n303), .A3(new_n736), .A4(new_n364), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n240), .ZN(G27));
  OAI21_X1  g595(.A(new_n745), .B1(new_n568), .B2(new_n573), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n751), .B(new_n719), .C1(new_n294), .C2(new_n302), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT101), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n359), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n348), .A2(new_n349), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n307), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT101), .A3(G469), .A4(new_n356), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(new_n354), .A3(new_n361), .A4(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n783), .A2(new_n736), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n782), .A2(KEYINPUT42), .A3(new_n790), .A4(new_n653), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n585), .A3(KEYINPUT102), .A4(new_n653), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT102), .B1(new_n746), .B2(new_n790), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G131), .ZN(G33));
  AND3_X1   g611(.A1(new_n715), .A2(new_n783), .A3(new_n789), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n746), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  AOI21_X1  g614(.A(new_n433), .B1(new_n669), .B2(new_n668), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT43), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT105), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n661), .A3(new_n703), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT44), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n294), .A2(new_n302), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n719), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(KEYINPUT44), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n787), .A2(new_n356), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT45), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(G469), .A3(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(new_n361), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n814), .A2(KEYINPUT103), .A3(KEYINPUT46), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT103), .B1(new_n814), .B2(KEYINPUT46), .ZN(new_n816));
  OAI221_X1 g630(.A(new_n354), .B1(KEYINPUT46), .B2(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n364), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n722), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT104), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n818), .A2(KEYINPUT104), .A3(new_n722), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n809), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n314), .ZN(G39));
  INV_X1    g638(.A(new_n807), .ZN(new_n825));
  INV_X1    g639(.A(new_n736), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n585), .A2(new_n825), .A3(new_n653), .A4(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n818), .A2(KEYINPUT47), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n818), .A2(KEYINPUT47), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G140), .ZN(G42));
  NOR3_X1   g645(.A1(new_n652), .A2(new_n365), .A3(new_n719), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT106), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n778), .B(KEYINPUT49), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n834), .A2(new_n726), .A3(new_n801), .ZN(new_n835));
  INV_X1    g649(.A(new_n731), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT107), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n687), .A2(new_n498), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n582), .A2(new_n569), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n775), .A2(new_n840), .A3(new_n841), .A4(new_n443), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n367), .A3(new_n703), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n491), .A2(new_n496), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n433), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n303), .A2(new_n441), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n656), .A2(new_n846), .A3(new_n660), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n839), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n845), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n663), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n657), .A2(new_n661), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n706), .A2(new_n851), .A3(KEYINPUT107), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n657), .A2(new_n661), .A3(new_n672), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n848), .A2(new_n852), .A3(new_n654), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n759), .A2(new_n764), .A3(new_n773), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n753), .B2(new_n755), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n362), .A2(new_n366), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n725), .A2(new_n295), .A3(new_n844), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n685), .A2(new_n713), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n585), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n790), .A2(new_n768), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n864), .A2(new_n718), .B1(new_n746), .B2(new_n798), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n855), .A2(new_n796), .A3(new_n857), .A4(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n687), .A2(new_n498), .A3(new_n433), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n751), .B1(new_n439), .B2(new_n712), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n295), .A2(new_n294), .A3(new_n302), .A4(new_n868), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n703), .A2(new_n867), .A3(new_n869), .A4(new_n789), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n731), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n777), .A2(new_n779), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n716), .A2(new_n737), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT52), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n826), .B1(new_n742), .B2(new_n745), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n875), .A2(new_n704), .B1(new_n870), .B2(new_n731), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n714), .B1(new_n742), .B2(new_n745), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n780), .B1(new_n877), .B2(new_n704), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n866), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n857), .A2(KEYINPUT53), .A3(new_n796), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n874), .A2(new_n880), .A3(KEYINPUT108), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT108), .B1(new_n874), .B2(new_n880), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT110), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT109), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n585), .A2(new_n861), .B1(new_n790), .B2(new_n768), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n799), .B1(new_n891), .B2(new_n703), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n854), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT107), .B1(new_n706), .B2(new_n851), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n654), .A2(new_n853), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n865), .A3(KEYINPUT109), .A4(new_n852), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n888), .A2(new_n889), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n857), .A2(new_n796), .A3(KEYINPUT53), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT108), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n873), .A2(KEYINPUT52), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n879), .B1(new_n876), .B2(new_n878), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n874), .A2(new_n880), .A3(KEYINPUT108), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n893), .A2(new_n897), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT110), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n838), .B(new_n884), .C1(new_n899), .C2(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT111), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(KEYINPUT111), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n882), .A2(KEYINPUT53), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n904), .A2(new_n905), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n866), .A2(KEYINPUT53), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n910), .B(new_n911), .C1(new_n838), .C2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n782), .A2(new_n653), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n783), .A2(new_n438), .A3(new_n778), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n802), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n653), .A2(new_n802), .A3(new_n438), .A4(new_n768), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n303), .A3(new_n752), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n836), .A2(new_n653), .A3(new_n919), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n433), .A3(new_n670), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n437), .B(KEYINPUT112), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n923), .A2(new_n925), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT114), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n924), .A2(new_n719), .A3(new_n726), .A4(new_n752), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT50), .Z(new_n932));
  NOR2_X1   g746(.A1(new_n433), .A2(new_n670), .ZN(new_n933));
  INV_X1    g747(.A(new_n777), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n926), .A2(new_n933), .B1(new_n934), .B2(new_n920), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n828), .A2(new_n829), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n366), .B2(new_n750), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n924), .A2(new_n807), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n930), .B1(new_n940), .B2(KEYINPUT51), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n917), .B(new_n941), .C1(KEYINPUT51), .C2(new_n940), .ZN(new_n942));
  NOR2_X1   g756(.A1(G952), .A2(G953), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT115), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n837), .B1(new_n942), .B2(new_n944), .ZN(G75));
  NOR2_X1   g759(.A1(new_n387), .A2(G952), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n298), .A2(new_n299), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n300), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n884), .B1(new_n899), .B2(new_n908), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(new_n282), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n188), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT56), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g770(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n957));
  AND2_X1   g771(.A1(new_n950), .A2(new_n957), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n946), .B(new_n956), .C1(new_n954), .C2(new_n958), .ZN(G51));
  NAND2_X1  g773(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(KEYINPUT118), .A3(new_n909), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT118), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n951), .A2(new_n962), .A3(KEYINPUT54), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n360), .B(KEYINPUT57), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT119), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n961), .A2(KEYINPUT119), .A3(new_n963), .A4(new_n964), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n352), .A3(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n952), .A2(new_n282), .A3(new_n813), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT120), .ZN(new_n973));
  INV_X1    g787(.A(new_n946), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n352), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n965), .B2(new_n966), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n970), .B1(new_n977), .B2(new_n968), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT120), .B1(new_n978), .B2(new_n946), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n975), .A2(new_n979), .ZN(G54));
  NAND3_X1  g794(.A1(new_n953), .A2(KEYINPUT58), .A3(G475), .ZN(new_n981));
  INV_X1    g795(.A(new_n424), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT121), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n946), .B1(new_n981), .B2(new_n982), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(G60));
  OR2_X1    g802(.A1(new_n666), .A2(new_n667), .ZN(new_n989));
  NAND2_X1  g803(.A1(G478), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT59), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n989), .B1(new_n917), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n961), .A2(new_n963), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n989), .A2(new_n991), .ZN(new_n994));
  AOI211_X1 g808(.A(new_n946), .B(new_n992), .C1(new_n993), .C2(new_n994), .ZN(G63));
  XNOR2_X1  g809(.A(new_n700), .B(KEYINPUT123), .ZN(new_n996));
  NAND2_X1  g810(.A1(G217), .A2(G902), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT60), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n952), .B2(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n999), .A2(new_n974), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n952), .A2(new_n998), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n696), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1000), .A2(KEYINPUT61), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(KEYINPUT122), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT122), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1001), .A2(new_n1005), .A3(new_n696), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1004), .A2(new_n1000), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT124), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT61), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1008), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1003), .B1(new_n1010), .B2(new_n1011), .ZN(G66));
  OAI21_X1  g826(.A(G953), .B1(new_n435), .B2(new_n256), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT125), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n855), .A2(new_n857), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1014), .B1(new_n1015), .B2(new_n387), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n947), .B1(G898), .B2(new_n387), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1016), .B(new_n1017), .Z(G69));
  AOI211_X1 g832(.A(new_n723), .B(new_n825), .C1(new_n671), .C2(new_n849), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n746), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n878), .A2(new_n737), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(new_n734), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT62), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n830), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n1024), .A2(new_n823), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n550), .B1(KEYINPUT30), .B2(new_n542), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(new_n419), .Z(new_n1027));
  NAND3_X1  g841(.A1(new_n1025), .A2(new_n387), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(G953), .B1(new_n305), .B2(new_n709), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AND4_X1   g845(.A1(new_n737), .A2(new_n796), .A3(new_n799), .A4(new_n878), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n830), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n918), .A2(new_n772), .ZN(new_n1034));
  AOI22_X1  g848(.A1(new_n821), .A2(new_n822), .B1(new_n809), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(KEYINPUT126), .ZN(new_n1036));
  OR3_X1    g850(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1036), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1037), .A2(new_n387), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1039), .B1(new_n709), .B2(new_n387), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1027), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1031), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1042), .B(new_n1043), .ZN(G72));
  NAND4_X1  g858(.A1(new_n1037), .A2(new_n857), .A3(new_n855), .A4(new_n1038), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  AOI211_X1 g861(.A(new_n538), .B(new_n554), .C1(new_n1045), .C2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1047), .B1(new_n1025), .B2(new_n1015), .ZN(new_n1049));
  AND2_X1   g863(.A1(new_n1049), .A2(new_n729), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1047), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n564), .A2(new_n565), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1052), .B1(new_n555), .B2(new_n554), .ZN(new_n1053));
  NOR3_X1   g867(.A1(new_n916), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  NOR4_X1   g868(.A1(new_n1048), .A2(new_n946), .A3(new_n1050), .A4(new_n1054), .ZN(G57));
endmodule


