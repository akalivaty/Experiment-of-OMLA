

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n771), .A2(n521), .ZN(n772) );
  NAND2_X4 U555 ( .A1(n784), .A2(n685), .ZN(n733) );
  AND2_X1 U556 ( .A1(n696), .A2(n520), .ZN(n697) );
  OR2_X1 U557 ( .A1(n728), .A2(n717), .ZN(n719) );
  OR2_X1 U558 ( .A1(n727), .A2(n716), .ZN(n717) );
  INV_X1 U559 ( .A(KEYINPUT95), .ZN(n706) );
  NOR2_X1 U560 ( .A1(n705), .A2(n704), .ZN(n707) );
  NOR2_X1 U561 ( .A1(n733), .A2(n1000), .ZN(n693) );
  XNOR2_X1 U562 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n718) );
  NOR2_X2 U563 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X1 U564 ( .A(n767), .B(KEYINPUT101), .ZN(n771) );
  XNOR2_X1 U565 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X2 U566 ( .A(KEYINPUT17), .B(n523), .Z(n879) );
  AND2_X1 U567 ( .A1(n695), .A2(n694), .ZN(n520) );
  OR2_X1 U568 ( .A1(n770), .A2(n769), .ZN(n521) );
  NOR2_X1 U569 ( .A1(n770), .A2(n756), .ZN(n522) );
  INV_X1 U570 ( .A(n927), .ZN(n695) );
  INV_X1 U571 ( .A(KEYINPUT71), .ZN(n591) );
  XNOR2_X1 U572 ( .A(n591), .B(KEYINPUT15), .ZN(n592) );
  XNOR2_X1 U573 ( .A(n593), .B(n592), .ZN(n700) );
  NOR2_X2 U574 ( .A1(G2104), .A2(n528), .ZN(n875) );
  NAND2_X1 U575 ( .A1(n879), .A2(G138), .ZN(n525) );
  INV_X1 U576 ( .A(G2105), .ZN(n528) );
  AND2_X1 U577 ( .A1(n528), .A2(G2104), .ZN(n880) );
  NAND2_X1 U578 ( .A1(G102), .A2(n880), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n525), .A2(n524), .ZN(n527) );
  INV_X1 U580 ( .A(KEYINPUT85), .ZN(n526) );
  XNOR2_X1 U581 ( .A(n527), .B(n526), .ZN(n533) );
  NAND2_X1 U582 ( .A1(G126), .A2(n875), .ZN(n530) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U584 ( .A1(G114), .A2(n876), .ZN(n529) );
  NAND2_X1 U585 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U586 ( .A(KEYINPUT84), .B(n531), .ZN(n532) );
  NOR2_X1 U587 ( .A1(n533), .A2(n532), .ZN(G164) );
  XNOR2_X1 U588 ( .A(G651), .B(KEYINPUT65), .ZN(n538) );
  NOR2_X1 U589 ( .A1(G543), .A2(n538), .ZN(n534) );
  XOR2_X2 U590 ( .A(KEYINPUT1), .B(n534), .Z(n636) );
  NAND2_X1 U591 ( .A1(G65), .A2(n636), .ZN(n537) );
  XOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  NOR2_X1 U593 ( .A1(G651), .A2(n632), .ZN(n535) );
  XNOR2_X1 U594 ( .A(KEYINPUT64), .B(n535), .ZN(n586) );
  NAND2_X1 U595 ( .A1(G53), .A2(n586), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n542) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n637) );
  NAND2_X1 U598 ( .A1(G91), .A2(n637), .ZN(n540) );
  NOR2_X1 U599 ( .A1(n632), .A2(n538), .ZN(n641) );
  NAND2_X1 U600 ( .A1(G78), .A2(n641), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  OR2_X1 U602 ( .A1(n542), .A2(n541), .ZN(G299) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  INV_X1 U605 ( .A(G120), .ZN(G236) );
  INV_X1 U606 ( .A(G69), .ZN(G235) );
  INV_X1 U607 ( .A(G108), .ZN(G238) );
  NAND2_X1 U608 ( .A1(G88), .A2(n637), .ZN(n544) );
  NAND2_X1 U609 ( .A1(G75), .A2(n641), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U611 ( .A1(G62), .A2(n636), .ZN(n546) );
  NAND2_X1 U612 ( .A1(G50), .A2(n586), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(G166) );
  NAND2_X1 U615 ( .A1(G63), .A2(n636), .ZN(n550) );
  NAND2_X1 U616 ( .A1(G51), .A2(n586), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT6), .B(n551), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n637), .A2(G89), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U621 ( .A1(G76), .A2(n641), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(KEYINPUT5), .B(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(KEYINPUT73), .B(n556), .ZN(n557) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT75), .B(KEYINPUT7), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(KEYINPUT74), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G168) );
  XOR2_X1 U629 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U632 ( .A(KEYINPUT69), .B(KEYINPUT11), .Z(n564) );
  INV_X1 U633 ( .A(G223), .ZN(n829) );
  NAND2_X1 U634 ( .A1(G567), .A2(n829), .ZN(n563) );
  XNOR2_X1 U635 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U636 ( .A(KEYINPUT68), .B(n565), .Z(G234) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n567) );
  NAND2_X1 U638 ( .A1(G56), .A2(n636), .ZN(n566) );
  XNOR2_X1 U639 ( .A(n567), .B(n566), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n637), .A2(G81), .ZN(n568) );
  XNOR2_X1 U641 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U642 ( .A1(G68), .A2(n641), .ZN(n569) );
  NAND2_X1 U643 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n571), .Z(n572) );
  NOR2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G43), .A2(n586), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n927) );
  INV_X1 U648 ( .A(G860), .ZN(n599) );
  OR2_X1 U649 ( .A1(n927), .A2(n599), .ZN(G153) );
  NAND2_X1 U650 ( .A1(n637), .A2(G90), .ZN(n576) );
  XNOR2_X1 U651 ( .A(n576), .B(KEYINPUT66), .ZN(n578) );
  NAND2_X1 U652 ( .A1(G77), .A2(n641), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U654 ( .A(KEYINPUT9), .B(n579), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n586), .A2(G52), .ZN(n581) );
  NAND2_X1 U656 ( .A1(G64), .A2(n636), .ZN(n580) );
  AND2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G66), .A2(n636), .ZN(n585) );
  NAND2_X1 U660 ( .A1(G92), .A2(n637), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G79), .A2(n641), .ZN(n588) );
  NAND2_X1 U663 ( .A1(G54), .A2(n586), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n593) );
  NOR2_X1 U666 ( .A1(G868), .A2(n700), .ZN(n595) );
  INV_X1 U667 ( .A(G868), .ZN(n659) );
  NOR2_X1 U668 ( .A1(n659), .A2(G301), .ZN(n594) );
  NOR2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U670 ( .A(KEYINPUT72), .B(n596), .ZN(G284) );
  NAND2_X1 U671 ( .A1(G868), .A2(G286), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G299), .A2(n659), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n599), .A2(G559), .ZN(n600) );
  INV_X1 U675 ( .A(n700), .ZN(n920) );
  NAND2_X1 U676 ( .A1(n600), .A2(n920), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n927), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n920), .A2(G868), .ZN(n602) );
  NOR2_X1 U680 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G123), .A2(n875), .ZN(n605) );
  XNOR2_X1 U683 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n880), .A2(G99), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G135), .A2(n879), .ZN(n609) );
  NAND2_X1 U687 ( .A1(G111), .A2(n876), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n949) );
  XNOR2_X1 U690 ( .A(G2096), .B(n949), .ZN(n613) );
  INV_X1 U691 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U693 ( .A1(G559), .A2(n920), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n614), .B(n927), .ZN(n655) );
  NOR2_X1 U695 ( .A1(n655), .A2(G860), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G67), .A2(n636), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G93), .A2(n637), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G80), .A2(n641), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G55), .A2(n586), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n658) );
  XOR2_X1 U703 ( .A(n621), .B(n658), .Z(G145) );
  AND2_X1 U704 ( .A1(n636), .A2(G60), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G85), .A2(n637), .ZN(n623) );
  NAND2_X1 U706 ( .A1(G47), .A2(n586), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n641), .A2(G72), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(G290) );
  NAND2_X1 U711 ( .A1(G651), .A2(G74), .ZN(n629) );
  NAND2_X1 U712 ( .A1(G49), .A2(n586), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U714 ( .A1(n636), .A2(n630), .ZN(n631) );
  XNOR2_X1 U715 ( .A(KEYINPUT76), .B(n631), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n632), .A2(G87), .ZN(n633) );
  XOR2_X1 U717 ( .A(KEYINPUT77), .B(n633), .Z(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G48), .A2(n586), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G61), .A2(n636), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G86), .A2(n637), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U723 ( .A(KEYINPUT78), .B(n640), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n641), .A2(G73), .ZN(n642) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n647), .Z(G305) );
  XNOR2_X1 U729 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n649) );
  XNOR2_X1 U730 ( .A(G290), .B(KEYINPUT19), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n649), .B(n648), .ZN(n652) );
  XNOR2_X1 U732 ( .A(G166), .B(G299), .ZN(n650) );
  XNOR2_X1 U733 ( .A(n650), .B(G288), .ZN(n651) );
  XNOR2_X1 U734 ( .A(n652), .B(n651), .ZN(n654) );
  XOR2_X1 U735 ( .A(G305), .B(n658), .Z(n653) );
  XNOR2_X1 U736 ( .A(n654), .B(n653), .ZN(n899) );
  XNOR2_X1 U737 ( .A(KEYINPUT82), .B(n655), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n899), .B(n656), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U748 ( .A(KEYINPUT67), .B(G82), .ZN(G220) );
  NOR2_X1 U749 ( .A1(G235), .A2(G236), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n666), .B(KEYINPUT83), .ZN(n667) );
  NOR2_X1 U751 ( .A1(G238), .A2(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(G57), .A2(n668), .ZN(n833) );
  NAND2_X1 U753 ( .A1(n833), .A2(G567), .ZN(n673) );
  NOR2_X1 U754 ( .A1(G219), .A2(G220), .ZN(n669) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U756 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U757 ( .A1(G96), .A2(n671), .ZN(n834) );
  NAND2_X1 U758 ( .A1(n834), .A2(G2106), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n673), .A2(n672), .ZN(n835) );
  NAND2_X1 U760 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U761 ( .A1(n835), .A2(n674), .ZN(n832) );
  NAND2_X1 U762 ( .A1(n832), .A2(G36), .ZN(G176) );
  NAND2_X1 U763 ( .A1(n879), .A2(G137), .ZN(n677) );
  NAND2_X1 U764 ( .A1(G101), .A2(n880), .ZN(n675) );
  XOR2_X1 U765 ( .A(KEYINPUT23), .B(n675), .Z(n676) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(n684) );
  NAND2_X1 U767 ( .A1(G125), .A2(n875), .ZN(n679) );
  NAND2_X1 U768 ( .A1(G113), .A2(n876), .ZN(n678) );
  NAND2_X1 U769 ( .A1(n679), .A2(n678), .ZN(n682) );
  NOR2_X1 U770 ( .A1(n684), .A2(n682), .ZN(G160) );
  INV_X1 U771 ( .A(G166), .ZN(G303) );
  NOR2_X1 U772 ( .A1(G2090), .A2(G303), .ZN(n680) );
  NAND2_X1 U773 ( .A1(G8), .A2(n680), .ZN(n748) );
  NOR2_X2 U774 ( .A1(G164), .A2(G1384), .ZN(n784) );
  INV_X1 U775 ( .A(G40), .ZN(n681) );
  OR2_X1 U776 ( .A1(n682), .A2(n681), .ZN(n683) );
  OR2_X1 U777 ( .A1(n684), .A2(n683), .ZN(n785) );
  INV_X1 U778 ( .A(n785), .ZN(n685) );
  INV_X1 U779 ( .A(G2072), .ZN(n958) );
  NOR2_X1 U780 ( .A1(n733), .A2(n958), .ZN(n687) );
  XNOR2_X1 U781 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n686) );
  XNOR2_X1 U782 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n733), .A2(G1956), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n703) );
  NAND2_X1 U785 ( .A1(G299), .A2(n703), .ZN(n690) );
  XOR2_X1 U786 ( .A(KEYINPUT28), .B(n690), .Z(n709) );
  NAND2_X1 U787 ( .A1(G1348), .A2(n733), .ZN(n692) );
  INV_X1 U788 ( .A(n733), .ZN(n711) );
  NAND2_X1 U789 ( .A1(G2067), .A2(n711), .ZN(n691) );
  NAND2_X1 U790 ( .A1(n692), .A2(n691), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n698) );
  INV_X1 U792 ( .A(G1996), .ZN(n1000) );
  XOR2_X1 U793 ( .A(n693), .B(KEYINPUT26), .Z(n696) );
  NAND2_X1 U794 ( .A1(n733), .A2(G1341), .ZN(n694) );
  NOR2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n702) );
  AND2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n703), .A2(G299), .ZN(n704) );
  XNOR2_X1 U799 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U801 ( .A(n710), .B(KEYINPUT29), .ZN(n715) );
  NAND2_X1 U802 ( .A1(G1961), .A2(n733), .ZN(n713) );
  XOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .Z(n1001) );
  NAND2_X1 U804 ( .A1(n711), .A2(n1001), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n721) );
  OR2_X1 U806 ( .A1(n721), .A2(G301), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n738) );
  NAND2_X1 U808 ( .A1(G8), .A2(n733), .ZN(n770) );
  NOR2_X1 U809 ( .A1(G1966), .A2(n770), .ZN(n728) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n733), .ZN(n727) );
  INV_X1 U811 ( .A(G8), .ZN(n716) );
  NOR2_X1 U812 ( .A1(G168), .A2(n720), .ZN(n724) );
  NAND2_X1 U813 ( .A1(G301), .A2(n721), .ZN(n722) );
  XNOR2_X1 U814 ( .A(n722), .B(KEYINPUT97), .ZN(n723) );
  NOR2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U816 ( .A(n725), .B(KEYINPUT98), .Z(n726) );
  XNOR2_X1 U817 ( .A(KEYINPUT31), .B(n726), .ZN(n739) );
  AND2_X1 U818 ( .A1(n738), .A2(n739), .ZN(n731) );
  AND2_X1 U819 ( .A1(G8), .A2(n727), .ZN(n729) );
  OR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  OR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n747) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n770), .ZN(n732) );
  XNOR2_X1 U823 ( .A(KEYINPUT99), .B(n732), .ZN(n736) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U825 ( .A1(G166), .A2(n734), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  OR2_X1 U827 ( .A1(n716), .A2(n737), .ZN(n741) );
  AND2_X1 U828 ( .A1(n738), .A2(n741), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n744) );
  INV_X1 U830 ( .A(n741), .ZN(n742) );
  OR2_X1 U831 ( .A1(n742), .A2(G286), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT32), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n755) );
  NAND2_X1 U835 ( .A1(n748), .A2(n755), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n749), .A2(n770), .ZN(n766) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U838 ( .A1(G288), .A2(G1976), .ZN(n750) );
  XNOR2_X1 U839 ( .A(n750), .B(KEYINPUT100), .ZN(n759) );
  NOR2_X1 U840 ( .A1(n751), .A2(n759), .ZN(n753) );
  INV_X1 U841 ( .A(KEYINPUT33), .ZN(n752) );
  AND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n764) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n930) );
  INV_X1 U845 ( .A(n930), .ZN(n756) );
  OR2_X1 U846 ( .A1(KEYINPUT33), .A2(n522), .ZN(n758) );
  XNOR2_X1 U847 ( .A(G1981), .B(G305), .ZN(n933) );
  INV_X1 U848 ( .A(n933), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n762) );
  INV_X1 U850 ( .A(n759), .ZN(n936) );
  NOR2_X1 U851 ( .A1(n770), .A2(n936), .ZN(n760) );
  AND2_X1 U852 ( .A1(KEYINPUT33), .A2(n760), .ZN(n761) );
  NOR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XOR2_X1 U857 ( .A(n768), .B(KEYINPUT24), .Z(n769) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT102), .ZN(n788) );
  XNOR2_X1 U859 ( .A(KEYINPUT37), .B(G2067), .ZN(n821) );
  NAND2_X1 U860 ( .A1(n880), .A2(G104), .ZN(n773) );
  XOR2_X1 U861 ( .A(KEYINPUT87), .B(n773), .Z(n775) );
  NAND2_X1 U862 ( .A1(n879), .A2(G140), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U864 ( .A(KEYINPUT34), .B(n776), .ZN(n782) );
  NAND2_X1 U865 ( .A1(G128), .A2(n875), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G116), .A2(n876), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U868 ( .A(KEYINPUT88), .B(n779), .Z(n780) );
  XNOR2_X1 U869 ( .A(KEYINPUT35), .B(n780), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n783), .ZN(n896) );
  NOR2_X1 U872 ( .A1(n821), .A2(n896), .ZN(n967) );
  NOR2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n786), .B(KEYINPUT86), .ZN(n824) );
  NAND2_X1 U875 ( .A1(n967), .A2(n824), .ZN(n819) );
  INV_X1 U876 ( .A(n819), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n810) );
  INV_X1 U878 ( .A(n824), .ZN(n808) );
  NAND2_X1 U879 ( .A1(G131), .A2(n879), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G119), .A2(n875), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G95), .A2(n880), .ZN(n791) );
  XNOR2_X1 U883 ( .A(KEYINPUT89), .B(n791), .ZN(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n876), .A2(G107), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n872) );
  XNOR2_X1 U887 ( .A(KEYINPUT90), .B(G1991), .ZN(n1010) );
  NAND2_X1 U888 ( .A1(n872), .A2(n1010), .ZN(n806) );
  NAND2_X1 U889 ( .A1(n880), .A2(G105), .ZN(n797) );
  XNOR2_X1 U890 ( .A(KEYINPUT38), .B(KEYINPUT92), .ZN(n796) );
  XNOR2_X1 U891 ( .A(n797), .B(n796), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G141), .A2(n879), .ZN(n799) );
  NAND2_X1 U893 ( .A1(G129), .A2(n875), .ZN(n798) );
  NAND2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U895 ( .A1(G117), .A2(n876), .ZN(n800) );
  XNOR2_X1 U896 ( .A(KEYINPUT91), .B(n800), .ZN(n801) );
  NOR2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n873) );
  NAND2_X1 U899 ( .A1(G1996), .A2(n873), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U901 ( .A(KEYINPUT93), .B(n807), .ZN(n956) );
  NOR2_X1 U902 ( .A1(n808), .A2(n956), .ZN(n816) );
  INV_X1 U903 ( .A(n816), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U905 ( .A(n811), .B(KEYINPUT103), .ZN(n813) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n924) );
  NAND2_X1 U907 ( .A1(n924), .A2(n824), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n827) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n873), .ZN(n947) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U911 ( .A1(n1010), .A2(n872), .ZN(n950) );
  NOR2_X1 U912 ( .A1(n814), .A2(n950), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U914 ( .A1(n947), .A2(n817), .ZN(n818) );
  XNOR2_X1 U915 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n821), .A2(n896), .ZN(n964) );
  NAND2_X1 U918 ( .A1(n822), .A2(n964), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n825), .B(KEYINPUT104), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U923 ( .A(G301), .ZN(G171) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U926 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n835), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2474), .B(G1971), .Z(n837) );
  XNOR2_X1 U935 ( .A(G1986), .B(G1956), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U937 ( .A(n838), .B(KEYINPUT107), .Z(n840) );
  XNOR2_X1 U938 ( .A(G1991), .B(G1996), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(G1976), .B(G1961), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1981), .B(G1966), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G229) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2090), .B(G2678), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n849), .B(KEYINPUT106), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(G2100), .Z(n853) );
  XNOR2_X1 U953 ( .A(G2084), .B(G2078), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U956 ( .A1(G124), .A2(n875), .ZN(n856) );
  XOR2_X1 U957 ( .A(KEYINPUT109), .B(n856), .Z(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G100), .A2(n880), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G136), .A2(n879), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G112), .A2(n876), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G139), .A2(n879), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G103), .A2(n880), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G127), .A2(n875), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G115), .A2(n876), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U971 ( .A(KEYINPUT110), .B(n868), .Z(n869) );
  XNOR2_X1 U972 ( .A(KEYINPUT47), .B(n869), .ZN(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n957) );
  XNOR2_X1 U974 ( .A(n957), .B(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n887) );
  NAND2_X1 U976 ( .A1(G130), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G142), .A2(n879), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G106), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(n887), .B(n886), .Z(n889) );
  XNOR2_X1 U985 ( .A(G164), .B(G160), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n893) );
  XOR2_X1 U987 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n891) );
  XNOR2_X1 U988 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U991 ( .A(G162), .B(n949), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U994 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n899), .B(G301), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n900), .B(n927), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n920), .B(n901), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n902), .B(G286), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U1000 ( .A(KEYINPUT105), .B(G2427), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G2435), .B(G2438), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n912) );
  XOR2_X1 U1003 ( .A(G2443), .B(G2430), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G2454), .B(G2446), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1006 ( .A(n908), .B(G2451), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G57), .ZN(G237) );
  INV_X1 U1019 ( .A(n919), .ZN(G401) );
  XOR2_X1 U1020 ( .A(KEYINPUT56), .B(G16), .Z(n945) );
  XNOR2_X1 U1021 ( .A(n920), .B(G1348), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(n921), .B(KEYINPUT117), .ZN(n943) );
  XNOR2_X1 U1023 ( .A(G171), .B(G1961), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G1956), .B(KEYINPUT118), .ZN(n922) );
  XNOR2_X1 U1025 ( .A(n922), .B(G299), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(G1341), .B(n927), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n938) );
  XOR2_X1 U1031 ( .A(G168), .B(G1966), .Z(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT57), .B(n934), .Z(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(G1971), .B(KEYINPUT119), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(n939), .B(G303), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n1029) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT51), .B(n948), .Z(n952) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n954) );
  XOR2_X1 U1046 ( .A(G160), .B(G2084), .Z(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n963) );
  XOR2_X1 U1049 ( .A(G164), .B(G2078), .Z(n960) );
  XNOR2_X1 U1050 ( .A(n958), .B(n957), .ZN(n959) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1052 ( .A(KEYINPUT50), .B(n961), .Z(n962) );
  NOR2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n965) );
  NAND2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1055 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1056 ( .A(KEYINPUT52), .B(n968), .Z(n969) );
  NOR2_X1 U1057 ( .A1(KEYINPUT55), .A2(n969), .ZN(n970) );
  XNOR2_X1 U1058 ( .A(KEYINPUT113), .B(n970), .ZN(n971) );
  NAND2_X1 U1059 ( .A1(n971), .A2(G29), .ZN(n1027) );
  XOR2_X1 U1060 ( .A(G1976), .B(G23), .Z(n974) );
  XNOR2_X1 U1061 ( .A(G1986), .B(KEYINPUT125), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(n972), .B(G24), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1064 ( .A(G22), .B(G1971), .ZN(n975) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1066 ( .A(KEYINPUT58), .B(n977), .Z(n996) );
  XNOR2_X1 U1067 ( .A(KEYINPUT123), .B(G1966), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n978), .B(G21), .ZN(n991) );
  XOR2_X1 U1069 ( .A(KEYINPUT121), .B(G4), .Z(n980) );
  XNOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n980), .B(n979), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G20), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G19), .B(G1341), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(KEYINPUT120), .B(G1981), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(G6), .B(n985), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n988), .B(KEYINPUT60), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT122), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(G5), .B(G1961), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1084 ( .A(KEYINPUT124), .B(n994), .Z(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1086 ( .A(n997), .B(KEYINPUT61), .Z(n998) );
  XNOR2_X1 U1087 ( .A(KEYINPUT126), .B(n998), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(G16), .A2(n999), .ZN(n1025) );
  XOR2_X1 U1089 ( .A(G29), .B(KEYINPUT116), .Z(n1022) );
  XNOR2_X1 U1090 ( .A(G32), .B(n1000), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G2067), .B(G26), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G27), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G33), .B(G2072), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT114), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(G28), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G25), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1013), .B(KEYINPUT115), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1014), .B(KEYINPUT53), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(G2084), .B(G34), .Z(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT54), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(G35), .B(G2090), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(n1020), .B(KEYINPUT55), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(G11), .A2(n1023), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1030), .Z(n1031) );
  XNOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1031), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

