//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n455), .A2(G567), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n466), .A2(new_n468), .A3(G137), .A4(new_n464), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n464), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n478), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n485), .B2(G124), .ZN(G162));
  NAND4_X1  g061(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n464), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n477), .A2(new_n489), .A3(G138), .A4(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT70), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(G62), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n506), .A2(G88), .A3(new_n507), .A4(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n512), .A2(G50), .A3(G543), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G166));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n506), .A2(new_n507), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n503), .A2(new_n505), .B1(KEYINPUT5), .B2(new_n502), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G63), .ZN(new_n528));
  NAND2_X1  g103(.A1(G76), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n521), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n524), .A2(new_n512), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n512), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT7), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n540), .B1(new_n529), .B2(new_n521), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n520), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n527), .A2(G63), .B1(KEYINPUT7), .B2(new_n530), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n544), .B(KEYINPUT74), .C1(new_n521), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n534), .A2(G90), .B1(G52), .B2(new_n538), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n521), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n534), .A2(G81), .B1(G43), .B2(new_n538), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n521), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT75), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n522), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n567), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n524), .A2(G91), .A3(new_n512), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n571), .A2(new_n574), .ZN(G299));
  OR2_X1    g150(.A1(new_n550), .A2(KEYINPUT78), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n550), .A2(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G301));
  AND2_X1   g153(.A1(new_n543), .A2(new_n546), .ZN(G286));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n518), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g156(.A(KEYINPUT79), .B(new_n511), .C1(new_n516), .C2(new_n517), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G303));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n533), .A2(new_n584), .B1(new_n585), .B2(new_n537), .ZN(new_n586));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n523), .A2(new_n587), .A3(new_n526), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n586), .B1(G651), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  NAND3_X1  g165(.A1(new_n524), .A2(G86), .A3(new_n512), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT81), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n524), .A2(new_n593), .A3(G86), .A4(new_n512), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n506), .A2(G61), .A3(new_n507), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n599), .A2(new_n600), .A3(G651), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT80), .B1(new_n602), .B2(new_n521), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n596), .A2(new_n601), .A3(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n534), .A2(G85), .B1(G47), .B2(new_n538), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n521), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(G290));
  AND3_X1   g186(.A1(new_n524), .A2(G92), .A3(new_n512), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n522), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n538), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G301), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G284));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G321));
  NAND2_X1  g198(.A1(G299), .A2(new_n619), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G168), .B2(new_n619), .ZN(G297));
  OAI21_X1  g200(.A(new_n624), .B1(G168), .B2(new_n619), .ZN(G280));
  INV_X1    g201(.A(new_n618), .ZN(new_n627));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n554), .A2(new_n619), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT83), .Z(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n632), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n485), .A2(G123), .ZN(new_n635));
  INV_X1    g210(.A(new_n478), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G135), .ZN(new_n637));
  NOR3_X1   g212(.A1(new_n464), .A2(KEYINPUT84), .A3(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(KEYINPUT84), .B1(new_n464), .B2(G111), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(G2104), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n635), .B(new_n637), .C1(new_n638), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n477), .A2(new_n473), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT14), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2443), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  INV_X1    g239(.A(G14), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n659), .B2(new_n660), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(KEYINPUT17), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n677), .C1(new_n678), .C2(new_n674), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n677), .A2(KEYINPUT18), .A3(new_n673), .ZN(new_n680));
  OAI21_X1  g255(.A(KEYINPUT18), .B1(new_n677), .B2(new_n673), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT86), .ZN(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(new_n690), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n691), .B1(KEYINPUT20), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n688), .A2(new_n692), .A3(new_n690), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n694), .B(new_n695), .C1(KEYINPUT20), .C2(new_n693), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT87), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1981), .B(G1986), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OR3_X1    g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n701), .B2(new_n702), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(G229));
  NOR2_X1   g282(.A1(G16), .A2(G23), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n589), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT33), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT90), .B(G16), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G22), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n518), .B2(new_n712), .ZN(new_n715));
  INV_X1    g290(.A(G1971), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G6), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(G16), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G305), .B2(G16), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT32), .B(G1981), .Z(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(new_n715), .B2(new_n716), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n718), .B(new_n723), .C1(new_n721), .C2(new_n722), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT34), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT34), .ZN(new_n726));
  MUX2_X1   g301(.A(G24), .B(G290), .S(new_n712), .Z(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G1986), .ZN(new_n728));
  NOR2_X1   g303(.A1(G25), .A2(G29), .ZN(new_n729));
  INV_X1    g304(.A(G131), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n464), .A2(G107), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n478), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n485), .B2(G119), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT88), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n729), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT35), .B(G1991), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT89), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G1986), .B2(new_n727), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n725), .A2(new_n726), .A3(new_n728), .A4(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT36), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(KEYINPUT36), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT92), .Z(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT30), .B(G28), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  OR2_X1    g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  NAND2_X1  g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n751), .A2(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n642), .B2(new_n752), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G33), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n473), .A2(G103), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT25), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(KEYINPUT25), .ZN(new_n760));
  INV_X1    g335(.A(G139), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n759), .B(new_n760), .C1(new_n761), .C2(new_n478), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n477), .A2(G127), .ZN(new_n763));
  NAND2_X1  g338(.A1(G115), .A2(G2104), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n464), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n757), .B1(new_n766), .B2(G29), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G2072), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT95), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n756), .B(new_n769), .C1(G2072), .C2(new_n767), .ZN(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(KEYINPUT24), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(KEYINPUT24), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n752), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G160), .B2(new_n752), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2084), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(G171), .A2(G16), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G5), .B2(G16), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n770), .B(new_n777), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n713), .A2(G20), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT23), .Z(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G299), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1956), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n780), .A2(new_n778), .ZN(new_n786));
  NOR2_X1   g361(.A1(G27), .A2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G164), .B2(G29), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n785), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G4), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n618), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1348), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n752), .A2(G35), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G162), .B2(new_n752), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2090), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n781), .A2(new_n791), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n752), .A2(G26), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G116), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G2105), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n636), .A2(G140), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT94), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n807), .B2(new_n806), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n485), .A2(G128), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n802), .B1(new_n811), .B2(new_n752), .ZN(new_n812));
  MUX2_X1   g387(.A(new_n802), .B(new_n812), .S(KEYINPUT28), .Z(new_n813));
  INV_X1    g388(.A(G2067), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n473), .A2(G105), .ZN(new_n816));
  NAND3_X1  g391(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT26), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n816), .B(new_n818), .C1(new_n636), .C2(G141), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n485), .A2(KEYINPUT97), .A3(G129), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT97), .B1(new_n485), .B2(G129), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT98), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G29), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G29), .B2(G32), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT27), .B(G1996), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n815), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n801), .A2(new_n831), .ZN(new_n832));
  MUX2_X1   g407(.A(G21), .B(G286), .S(G16), .Z(new_n833));
  INV_X1    g408(.A(G1966), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n713), .A2(G19), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n555), .B2(new_n713), .ZN(new_n837));
  MUX2_X1   g412(.A(new_n836), .B(new_n837), .S(KEYINPUT93), .Z(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G1341), .Z(new_n839));
  NAND4_X1  g414(.A1(new_n750), .A2(new_n832), .A3(new_n835), .A4(new_n839), .ZN(G150));
  INV_X1    g415(.A(G150), .ZN(G311));
  AOI22_X1  g416(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n521), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT99), .B(G55), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n534), .A2(G93), .B1(new_n538), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(G860), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT100), .B1(new_n843), .B2(new_n846), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(new_n845), .C1(new_n842), .C2(new_n521), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n851), .A2(new_n555), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n555), .B1(new_n851), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n851), .A2(new_n853), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n554), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n851), .A2(new_n555), .A3(new_n853), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n627), .A2(G559), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n858), .A2(new_n863), .A3(G559), .A4(new_n627), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT39), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT39), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n850), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n849), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n875), .A2(new_n871), .A3(KEYINPUT102), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n848), .B1(new_n874), .B2(new_n876), .ZN(G145));
  XOR2_X1   g452(.A(new_n734), .B(new_n645), .Z(new_n878));
  INV_X1    g453(.A(G142), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n464), .A2(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  OAI22_X1  g456(.A1(new_n478), .A2(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n485), .A2(G130), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(KEYINPUT105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(KEYINPUT105), .B2(new_n883), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n878), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n826), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n823), .B2(new_n825), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n811), .B(new_n496), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n823), .A2(new_n825), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(KEYINPUT103), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n896), .B2(new_n890), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n766), .B(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n893), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n893), .A2(new_n897), .B1(new_n898), .B2(new_n766), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n887), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n893), .A2(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n766), .A2(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n893), .A2(new_n897), .A3(new_n899), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(new_n886), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n642), .B(G160), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G162), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT107), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(KEYINPUT106), .B(G37), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n902), .B(new_n907), .C1(new_n915), .C2(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(new_n918), .ZN(G395));
  XNOR2_X1  g494(.A(G305), .B(G288), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n609), .A2(new_n518), .A3(new_n610), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n518), .B1(new_n609), .B2(new_n610), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G290), .A2(G166), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n922), .A3(new_n920), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n928), .A2(KEYINPUT109), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n929), .A2(KEYINPUT109), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(KEYINPUT109), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n631), .B(KEYINPUT83), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n856), .B(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(G299), .B(new_n618), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT41), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n937), .B2(new_n936), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n934), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n936), .A2(new_n937), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n943), .A2(new_n930), .A3(new_n933), .A4(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n941), .B1(new_n934), .B2(new_n940), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n619), .B1(new_n843), .B2(new_n846), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(G295));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n948), .ZN(G331));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n543), .A2(new_n546), .A3(new_n550), .ZN(new_n952));
  NAND3_X1  g527(.A1(G168), .A2(new_n576), .A3(new_n577), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n862), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n952), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n856), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n954), .A2(new_n938), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n937), .B1(new_n954), .B2(new_n956), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n938), .A3(new_n956), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n954), .A2(new_n956), .ZN(new_n961));
  OAI211_X1 g536(.A(KEYINPUT111), .B(new_n960), .C1(new_n961), .C2(new_n937), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n923), .A2(new_n924), .A3(new_n921), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n920), .B1(new_n926), .B2(new_n922), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n925), .A2(new_n927), .A3(KEYINPUT112), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n962), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n957), .A2(new_n958), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n970), .B2(new_n928), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT43), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n968), .B1(new_n957), .B2(new_n958), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n928), .B(new_n960), .C1(new_n961), .C2(new_n937), .ZN(new_n974));
  AND4_X1   g549(.A1(KEYINPUT43), .A2(new_n973), .A3(new_n914), .A4(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT44), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n969), .B2(new_n971), .ZN(new_n979));
  AND4_X1   g554(.A1(new_n978), .A2(new_n973), .A3(new_n914), .A4(new_n974), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n976), .A2(new_n981), .ZN(G397));
  INV_X1    g557(.A(KEYINPUT127), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n491), .B2(new_n495), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n469), .A2(new_n470), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G2105), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n472), .A2(new_n474), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(G40), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT113), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  NAND3_X1  g568(.A1(G160), .A2(new_n993), .A3(G40), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n987), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n811), .A2(new_n814), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n809), .A2(new_n810), .A3(G2067), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n826), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n999), .B2(new_n826), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n734), .B(new_n738), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(G290), .B(G1986), .Z(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n995), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n497), .A2(new_n1008), .A3(new_n499), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n986), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n992), .A2(new_n994), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1971), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G2090), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n497), .A2(new_n1014), .A3(new_n1008), .A4(new_n499), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n992), .A2(new_n994), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n985), .A2(new_n1017), .ZN(new_n1018));
  AND4_X1   g593(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(G8), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1022), .B(new_n1023), .C1(new_n581), .C2(new_n582), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n596), .A2(new_n1027), .A3(new_n601), .A4(new_n603), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n591), .A2(new_n595), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n603), .A2(new_n601), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G1981), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1028), .A2(new_n1031), .A3(KEYINPUT49), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1023), .B1(new_n1016), .B2(new_n984), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1032), .A2(KEYINPUT117), .A3(new_n1033), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n993), .B1(G160), .B2(G40), .ZN(new_n1042));
  INV_X1    g617(.A(G40), .ZN(new_n1043));
  NOR4_X1   g618(.A1(new_n471), .A2(new_n475), .A3(KEYINPUT113), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n984), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n588), .A2(G651), .ZN(new_n1046));
  INV_X1    g621(.A(new_n586), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(G1976), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1048), .A3(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n589), .A2(G1976), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(KEYINPUT52), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(KEYINPUT52), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1026), .A2(new_n1041), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n543), .A2(new_n546), .A3(G8), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1017), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n496), .A2(new_n1008), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(KEYINPUT50), .B2(new_n1009), .ZN(new_n1062));
  INV_X1    g637(.A(G2084), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n1008), .A4(new_n499), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(new_n1016), .A3(new_n987), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1062), .A2(new_n1063), .B1(new_n834), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT51), .B(new_n1058), .C1(new_n1066), .C2(new_n1023), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n834), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n992), .A2(new_n994), .B1(new_n984), .B2(new_n1059), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1068), .B(G8), .C1(new_n1073), .C2(G286), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(G8), .A3(G286), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1067), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n491), .A2(new_n498), .A3(new_n495), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n498), .B1(new_n491), .B2(new_n495), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1079), .A2(new_n1080), .A3(G1384), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1071), .B(new_n1013), .C1(new_n1081), .C2(new_n1014), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(G8), .B1(new_n1083), .B2(new_n1012), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1078), .B1(new_n1084), .B2(new_n1025), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n716), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1023), .B1(new_n1087), .B2(new_n1082), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n513), .A2(new_n515), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT71), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT79), .B1(new_n1092), .B2(new_n511), .ZN(new_n1093));
  INV_X1    g668(.A(new_n582), .ZN(new_n1094));
  OAI21_X1  g669(.A(G8), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1022), .ZN(new_n1096));
  NAND3_X1  g671(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1088), .A2(KEYINPUT115), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1085), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1064), .A2(new_n987), .A3(new_n789), .A4(new_n1016), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1103), .B2(new_n1102), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1010), .A2(new_n789), .A3(new_n1011), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1071), .B1(new_n1081), .B2(new_n1014), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1106), .A2(new_n1101), .B1(new_n1107), .B2(new_n778), .ZN(new_n1108));
  AOI21_X1  g683(.A(G301), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1057), .A2(new_n1077), .A3(new_n1100), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1067), .A2(new_n1076), .A3(new_n1074), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1111), .A2(KEYINPUT62), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G288), .A2(G1976), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1041), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1028), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1038), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1066), .A2(new_n1023), .A3(G286), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1084), .A2(new_n1025), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1041), .A4(new_n1056), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT63), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT63), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1085), .A2(new_n1099), .B1(new_n1122), .B2(new_n1118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1041), .A2(new_n1056), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1117), .B(new_n1121), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1113), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n987), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n991), .A2(KEYINPUT124), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n1130));
  NAND3_X1  g705(.A1(G160), .A2(new_n1130), .A3(G40), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1129), .A2(new_n1131), .A3(KEYINPUT53), .A4(new_n789), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1128), .A2(KEYINPUT125), .A3(new_n1132), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1108), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(G171), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1105), .A2(G301), .A3(new_n1108), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT54), .ZN(new_n1140));
  AND4_X1   g715(.A1(new_n1140), .A2(new_n1057), .A3(new_n1111), .A4(new_n1100), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1010), .A2(new_n1011), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n1145));
  INV_X1    g720(.A(G1956), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1145), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1143), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(G299), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n571), .A2(new_n574), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT120), .B1(new_n1157), .B2(new_n1154), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(KEYINPUT57), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(KEYINPUT121), .B(new_n1143), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1152), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1160), .B(new_n1143), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n814), .B(new_n984), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1107), .B2(new_n795), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(new_n618), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n618), .B1(new_n1167), .B2(KEYINPUT60), .ZN(new_n1170));
  AOI21_X1  g745(.A(G1348), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n1172));
  NOR4_X1   g747(.A1(new_n1171), .A2(new_n1172), .A3(new_n627), .A4(new_n1166), .ZN(new_n1173));
  OAI22_X1  g748(.A1(new_n1170), .A2(new_n1173), .B1(KEYINPUT60), .B2(new_n1167), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1164), .A2(KEYINPUT61), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT122), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1010), .A2(new_n999), .A3(new_n1011), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT58), .B(G1341), .Z(new_n1179));
  NAND2_X1  g754(.A1(new_n1045), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1177), .B1(new_n1181), .B2(new_n555), .ZN(new_n1182));
  XOR2_X1   g757(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1183));
  AOI211_X1 g758(.A(new_n1183), .B(new_n554), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1174), .A2(new_n1175), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1150), .A2(new_n1161), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT61), .B1(new_n1187), .B2(new_n1164), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1163), .B(new_n1169), .C1(new_n1186), .C2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT54), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1137), .A2(new_n621), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1190), .B1(new_n1191), .B2(new_n1109), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1141), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1007), .B1(new_n1126), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n738), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1001), .A2(new_n1195), .A3(new_n735), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n995), .B1(new_n1196), .B2(new_n997), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n995), .A2(new_n999), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT46), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n895), .A2(new_n996), .A3(new_n997), .ZN(new_n1200));
  INV_X1    g775(.A(new_n995), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT47), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1003), .A2(new_n995), .ZN(new_n1204));
  NOR3_X1   g779(.A1(G290), .A2(G1986), .A3(new_n1201), .ZN(new_n1205));
  XNOR2_X1  g780(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1197), .A2(new_n1203), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n983), .B1(new_n1194), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1026), .A2(new_n1056), .A3(new_n1041), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1211), .B1(new_n1085), .B2(new_n1099), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1212), .A2(new_n1192), .A3(new_n1140), .A4(new_n1111), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1143), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1215), .A2(KEYINPUT118), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1214), .B1(new_n1216), .B2(new_n1147), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1161), .B1(new_n1217), .B2(KEYINPUT121), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1162), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1169), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AND3_X1   g795(.A1(new_n1174), .A2(new_n1175), .A3(new_n1185), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1187), .A2(new_n1164), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1220), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1213), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1122), .A2(new_n1118), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1100), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1228), .A2(new_n1041), .A3(new_n1056), .ZN(new_n1229));
  AOI22_X1  g804(.A1(new_n1038), .A2(new_n1116), .B1(new_n1120), .B2(KEYINPUT63), .ZN(new_n1230));
  OAI211_X1 g805(.A(new_n1229), .B(new_n1230), .C1(new_n1112), .C2(new_n1110), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1006), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g807(.A(new_n1209), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1232), .A2(KEYINPUT127), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1210), .A2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g810(.A1(G227), .A2(new_n462), .ZN(new_n1237));
  AND4_X1   g811(.A1(new_n667), .A2(new_n705), .A3(new_n706), .A4(new_n1237), .ZN(new_n1238));
  OAI211_X1 g812(.A(new_n917), .B(new_n1238), .C1(new_n979), .C2(new_n980), .ZN(G225));
  INV_X1    g813(.A(G225), .ZN(G308));
endmodule


