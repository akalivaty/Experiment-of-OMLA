//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT66), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n203), .A2(new_n205), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n214), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n226), .A2(new_n227), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n210), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n221), .B1(KEYINPUT1), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n219), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n247), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n215), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G87), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(KEYINPUT22), .A3(G20), .ZN(new_n266));
  OR2_X1    g0066(.A1(KEYINPUT76), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT76), .A2(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(KEYINPUT3), .A3(new_n268), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n269), .A2(new_n216), .A3(G87), .A4(new_n257), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n264), .A2(new_n266), .B1(new_n270), .B2(KEYINPUT22), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT23), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(new_n216), .B2(G107), .ZN(new_n273));
  INV_X1    g0073(.A(G107), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(KEYINPUT23), .A3(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT76), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT76), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G116), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n276), .B1(new_n282), .B2(G20), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n271), .A2(new_n283), .A3(KEYINPUT24), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT24), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n264), .A2(new_n266), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n270), .A2(KEYINPUT22), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n281), .A2(new_n216), .B1(new_n273), .B2(new_n275), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n255), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(G1), .A2(G13), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G250), .A2(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G257), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(G1698), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(new_n269), .A3(new_n257), .ZN(new_n298));
  OAI21_X1  g0098(.A(G294), .B1(new_n277), .B2(new_n278), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT5), .B(G41), .ZN(new_n301));
  INV_X1    g0101(.A(G1), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G45), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n294), .ZN(new_n306));
  INV_X1    g0106(.A(G264), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n301), .A2(new_n294), .A3(new_n304), .A4(G274), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n311), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n300), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(new_n314), .B2(G200), .ZN(new_n315));
  INV_X1    g0115(.A(new_n255), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n302), .A2(G13), .A3(G20), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n317), .C1(G1), .C2(new_n258), .ZN(new_n318));
  INV_X1    g0118(.A(new_n317), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n274), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT25), .B1(new_n319), .B2(new_n274), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n318), .A2(new_n274), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n291), .A2(new_n315), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT89), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT24), .B1(new_n271), .B2(new_n283), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n288), .A2(new_n285), .A3(new_n289), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n323), .B1(new_n329), .B2(new_n255), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT89), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n315), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n264), .A2(G222), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n264), .A2(G223), .A3(G1698), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n335), .B(new_n336), .C1(new_n224), .C2(new_n264), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n294), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G41), .ZN(new_n342));
  INV_X1    g0142(.A(G45), .ZN(new_n343));
  AOI21_X1  g0143(.A(G1), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT68), .B1(new_n344), .B2(G274), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n302), .B(G274), .C1(G41), .C2(G45), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT68), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G226), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n342), .A2(new_n343), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n302), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n294), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n341), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(G179), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n255), .B1(new_n302), .B2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G50), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT8), .A2(G58), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(KEYINPUT71), .A2(G58), .ZN(new_n363));
  NOR2_X1   g0163(.A1(KEYINPUT71), .A2(G58), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT8), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n258), .A2(G20), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G150), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G20), .A2(G33), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n367), .A2(new_n369), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n207), .B2(G20), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n360), .B1(G50), .B2(new_n317), .C1(new_n374), .C2(new_n316), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n355), .B1(new_n339), .B2(new_n340), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(G169), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n358), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n375), .B(KEYINPUT9), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n357), .A2(G200), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(G190), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT10), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT10), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n379), .A2(new_n380), .A3(new_n384), .A4(new_n381), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n378), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G226), .A2(G1698), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n237), .B2(G1698), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n264), .A2(new_n388), .B1(G33), .B2(G97), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n389), .A2(new_n294), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n302), .A2(new_n352), .B1(new_n292), .B2(new_n293), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n349), .B1(G238), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n389), .B2(new_n294), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G200), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n319), .A2(new_n202), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT12), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n359), .A2(G68), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n369), .A2(new_n224), .B1(new_n216), .B2(G68), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n372), .A2(new_n219), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n255), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g0204(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n405));
  OAI211_X1 g0205(.A(new_n400), .B(new_n401), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n404), .A2(new_n405), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n398), .B(new_n408), .C1(new_n310), .C2(new_n397), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n394), .A2(new_n396), .A3(G179), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT74), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n391), .B1(new_n390), .B2(new_n393), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n395), .A2(KEYINPUT13), .ZN(new_n415));
  OAI21_X1  g0215(.A(G169), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n411), .A2(KEYINPUT74), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n397), .A2(G169), .A3(new_n417), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n409), .B1(new_n421), .B2(new_n408), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n417), .B1(new_n397), .B2(G169), .ZN(new_n424));
  INV_X1    g0224(.A(G169), .ZN(new_n425));
  AOI211_X1 g0225(.A(new_n425), .B(new_n418), .C1(new_n394), .C2(new_n396), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n412), .B(new_n410), .C1(new_n424), .C2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n408), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT75), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n409), .ZN(new_n431));
  INV_X1    g0231(.A(new_n367), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n359), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n367), .A2(new_n319), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(KEYINPUT71), .A2(G58), .ZN(new_n436));
  NAND2_X1  g0236(.A1(KEYINPUT71), .A2(G58), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n202), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(G20), .B1(new_n438), .B2(new_n218), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n371), .A2(G159), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(G20), .B1(new_n269), .B2(new_n257), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT7), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n202), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n257), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n279), .B2(KEYINPUT3), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT7), .B1(new_n446), .B2(G20), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n441), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n316), .B1(new_n448), .B2(KEYINPUT16), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT16), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n262), .A2(new_n216), .A3(new_n263), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n443), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n259), .A2(KEYINPUT77), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT77), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(new_n258), .A3(KEYINPUT3), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n453), .B(new_n455), .C1(new_n279), .C2(KEYINPUT3), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n443), .A2(G20), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n202), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n450), .B1(new_n459), .B2(new_n441), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n435), .B1(new_n449), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n344), .A2(KEYINPUT68), .A3(G274), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n346), .A2(new_n347), .ZN(new_n463));
  AOI22_X1  g0263(.A1(G232), .A2(new_n392), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n258), .A2(new_n265), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G223), .A2(G1698), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n351), .B2(G1698), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n446), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(KEYINPUT79), .B(new_n464), .C1(new_n468), .C2(new_n294), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT79), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n269), .A3(new_n257), .ZN(new_n471));
  INV_X1    g0271(.A(new_n465), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n294), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n345), .A2(new_n348), .B1(new_n354), .B2(new_n237), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n425), .ZN(new_n477));
  INV_X1    g0277(.A(G179), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n478), .B(new_n464), .C1(new_n468), .C2(new_n294), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT78), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n471), .A2(new_n472), .ZN(new_n482));
  INV_X1    g0282(.A(new_n294), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(KEYINPUT78), .A3(new_n478), .A4(new_n464), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n477), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT18), .B1(new_n461), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT17), .ZN(new_n489));
  INV_X1    g0289(.A(new_n435), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT69), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT69), .B1(new_n257), .B2(new_n259), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT7), .B1(new_n493), .B2(new_n216), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n456), .A2(new_n457), .ZN(new_n495));
  OAI21_X1  g0295(.A(G68), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n205), .B(new_n203), .C1(new_n365), .C2(new_n202), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G20), .B1(G159), .B2(new_n371), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT16), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n277), .A2(new_n278), .A3(new_n256), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n443), .B(new_n216), .C1(new_n500), .C2(new_n445), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G68), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n442), .A2(new_n443), .ZN(new_n503));
  OAI211_X1 g0303(.A(KEYINPUT16), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n255), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n490), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G200), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n473), .A2(new_n474), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n476), .A2(new_n507), .B1(new_n310), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n489), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT18), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n425), .A2(new_n476), .B1(new_n481), .B2(new_n485), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT79), .B1(new_n484), .B2(new_n464), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n473), .A2(new_n474), .A3(new_n470), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n507), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n508), .A2(new_n310), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n461), .A2(new_n518), .A3(KEYINPUT17), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n488), .A2(new_n510), .A3(new_n513), .A4(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n294), .B1(new_n493), .B2(new_n274), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G232), .A2(G1698), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n223), .B2(G1698), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n493), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n349), .B1(G244), .B2(new_n392), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n359), .A2(G77), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n319), .A2(new_n224), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g0330(.A(KEYINPUT8), .B(G58), .Z(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n371), .B1(G20), .B2(G77), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT15), .B(G87), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT72), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n537), .B2(new_n369), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n530), .B1(new_n538), .B2(new_n255), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n527), .B(new_n539), .C1(new_n310), .C2(new_n526), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n526), .B2(new_n425), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n524), .A2(new_n478), .A3(new_n525), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n520), .A2(new_n544), .ZN(new_n545));
  AND4_X1   g0345(.A1(new_n386), .A2(new_n423), .A3(new_n431), .A4(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G257), .A2(G1698), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n307), .B2(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n446), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G303), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n264), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n483), .ZN(new_n552));
  INV_X1    g0352(.A(G270), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n311), .B1(new_n306), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(KEYINPUT87), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n493), .A2(G303), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n294), .B1(new_n558), .B2(new_n549), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n559), .B2(new_n554), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n317), .A2(G116), .ZN(new_n561));
  INV_X1    g0361(.A(new_n318), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(G116), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G283), .ZN(new_n564));
  INV_X1    g0364(.A(G97), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n216), .C1(G33), .C2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n566), .B(new_n255), .C1(new_n216), .C2(G116), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT20), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n567), .B(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n425), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n556), .A2(new_n560), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n559), .A2(new_n478), .A3(new_n554), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n563), .A2(new_n569), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n556), .A2(new_n560), .A3(KEYINPUT21), .A4(new_n570), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n556), .A2(new_n560), .A3(G200), .ZN(new_n579));
  INV_X1    g0379(.A(new_n575), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(KEYINPUT88), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n556), .A2(new_n560), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G190), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(new_n580), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT88), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n578), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(G250), .B(G1698), .C1(new_n491), .C2(new_n492), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n225), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n334), .B(new_n591), .C1(new_n491), .C2(new_n492), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n589), .A2(new_n592), .A3(new_n564), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n225), .A2(G1698), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n446), .A2(KEYINPUT82), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n269), .A2(new_n257), .A3(new_n594), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT82), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n598), .A3(new_n590), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n294), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n311), .B1(new_n306), .B2(new_n296), .ZN(new_n601));
  OAI21_X1  g0401(.A(G200), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n595), .A2(new_n590), .A3(new_n598), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n589), .A2(new_n592), .A3(new_n564), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n483), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n601), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(G190), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n274), .B1(new_n452), .B2(new_n458), .ZN(new_n608));
  XNOR2_X1  g0408(.A(G97), .B(G107), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT6), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n610), .A2(new_n565), .A3(G107), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n613), .A2(new_n216), .B1(new_n224), .B2(new_n372), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n255), .B1(new_n608), .B2(new_n614), .ZN(new_n615));
  OR3_X1    g0415(.A1(new_n317), .A2(KEYINPUT80), .A3(G97), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT80), .B1(new_n317), .B2(G97), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n318), .C2(new_n565), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT81), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n602), .A2(new_n607), .A3(new_n615), .A4(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n425), .B1(new_n600), .B2(new_n601), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n615), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n605), .A2(new_n478), .A3(new_n606), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n291), .A2(new_n324), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n314), .A2(G169), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n478), .B2(new_n314), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n294), .A2(G250), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT83), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n303), .B(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n632), .A2(new_n634), .B1(G274), .B2(new_n304), .ZN(new_n635));
  NOR2_X1   g0435(.A1(G238), .A2(G1698), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n225), .B2(G1698), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n281), .B1(new_n446), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n635), .B(new_n478), .C1(new_n638), .C2(new_n294), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n635), .B1(new_n638), .B2(new_n294), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n425), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n446), .A2(new_n216), .A3(G68), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT19), .B1(new_n368), .B2(G97), .ZN(new_n645));
  NAND2_X1  g0445(.A1(G33), .A2(G97), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT19), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n216), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n265), .A2(new_n565), .A3(new_n274), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(new_n255), .B1(new_n319), .B2(new_n537), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT85), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n537), .B2(new_n318), .ZN(new_n654));
  INV_X1    g0454(.A(new_n537), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n562), .A3(KEYINPUT85), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n641), .A2(new_n643), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n304), .A2(G274), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n303), .B(KEYINPUT83), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n631), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n446), .A2(new_n637), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n282), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n663), .B2(new_n483), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G190), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT86), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(KEYINPUT86), .A3(G190), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n642), .A2(G200), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n655), .A2(new_n317), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n316), .B1(new_n644), .B2(new_n650), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n318), .A2(new_n265), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n667), .A2(new_n668), .A3(new_n669), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n658), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n626), .A2(new_n630), .A3(new_n675), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n333), .A2(new_n546), .A3(new_n588), .A4(new_n676), .ZN(G372));
  AND2_X1   g0477(.A1(new_n488), .A2(new_n513), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n510), .A2(new_n519), .ZN(new_n679));
  INV_X1    g0479(.A(new_n543), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n427), .A2(new_n428), .B1(new_n680), .B2(new_n409), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT91), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n409), .A2(new_n680), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n429), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n678), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n383), .A2(new_n385), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n378), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n330), .A2(new_n331), .A3(new_n315), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n331), .B1(new_n330), .B2(new_n315), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n657), .A2(new_n643), .A3(new_n639), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n673), .A2(new_n669), .A3(new_n665), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n621), .A3(new_n625), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT90), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n626), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT90), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n333), .A3(new_n698), .A4(new_n694), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n630), .A2(new_n578), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT26), .B1(new_n675), .B2(new_n625), .ZN(new_n702));
  INV_X1    g0502(.A(new_n625), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT26), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n694), .A3(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n702), .A2(new_n692), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n546), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n688), .A2(new_n708), .ZN(G369));
  NAND3_X1  g0509(.A1(new_n302), .A2(new_n216), .A3(G13), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G343), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n580), .A2(new_n716), .ZN(new_n717));
  MUX2_X1   g0517(.A(new_n588), .B(new_n578), .S(new_n717), .Z(new_n718));
  AND2_X1   g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(new_n630), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n627), .A2(new_n715), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n722), .B2(new_n691), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n630), .A2(new_n716), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n719), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n578), .A2(new_n716), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n726), .B1(new_n723), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(G399));
  NOR2_X1   g0532(.A1(new_n649), .A2(G116), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n211), .A2(new_n342), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(G1), .ZN(new_n735));
  INV_X1    g0535(.A(new_n220), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n642), .A2(new_n300), .A3(new_n308), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n574), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n605), .A2(new_n606), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n600), .A2(new_n601), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(KEYINPUT30), .A3(new_n574), .A4(new_n741), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n314), .A2(new_n664), .A3(G179), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n743), .A2(new_n747), .A3(new_n560), .A4(new_n556), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n715), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT31), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n676), .A2(new_n588), .A3(new_n333), .A4(new_n716), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n739), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n715), .B1(new_n701), .B2(new_n706), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n703), .A2(new_n694), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT26), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n703), .A2(new_n704), .A3(new_n658), .A4(new_n674), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n759), .A2(new_n692), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n700), .A2(new_n333), .A3(new_n697), .A4(new_n694), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(KEYINPUT29), .A3(new_n716), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n753), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n738), .B1(new_n765), .B2(G1), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT94), .Z(G364));
  INV_X1    g0567(.A(G13), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G45), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n771), .A2(G1), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n734), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n719), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G330), .B2(new_n718), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n215), .B1(G20), .B2(new_n425), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n446), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n211), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n252), .A2(new_n343), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n343), .C2(new_n220), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n264), .A2(new_n211), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(G116), .B2(new_n211), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n782), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n775), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n216), .A2(new_n310), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n507), .A2(G179), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n550), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n478), .A2(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n216), .A2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G329), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n797), .A2(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n478), .A2(new_n507), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n795), .B(new_n803), .C1(G326), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n799), .A2(new_n793), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G283), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n804), .A2(new_n799), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT33), .B(G317), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n799), .A2(new_n796), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n812), .A2(new_n813), .B1(new_n815), .B2(G311), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n216), .B1(new_n800), .B2(G190), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n264), .B1(G294), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n807), .A2(new_n810), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT96), .B(G159), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n801), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT32), .ZN(new_n823));
  INV_X1    g0623(.A(new_n797), .ZN(new_n824));
  INV_X1    g0624(.A(new_n365), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G50), .A2(new_n806), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n794), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G68), .A2(new_n812), .B1(new_n827), .B2(G87), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n823), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n815), .A2(G77), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n809), .A2(G107), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n818), .A2(G97), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n264), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n820), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT97), .ZN(new_n835));
  INV_X1    g0635(.A(new_n781), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n834), .B2(KEYINPUT97), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n791), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n780), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n718), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n777), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n526), .A2(new_n425), .ZN(new_n843));
  INV_X1    g0643(.A(new_n539), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n542), .A4(new_n715), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT99), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT99), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n541), .A2(new_n847), .A3(new_n542), .A4(new_n715), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n540), .B(new_n543), .C1(new_n539), .C2(new_n716), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT100), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(new_n849), .B2(new_n850), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n754), .B(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n753), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n775), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  INV_X1    g0659(.A(new_n775), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n781), .A2(new_n778), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(G77), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n811), .A2(new_n370), .ZN(new_n864));
  INV_X1    g0664(.A(G143), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n797), .A2(new_n865), .B1(new_n814), .B2(new_n821), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n864), .B(new_n866), .C1(G137), .C2(new_n806), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n446), .B1(new_n365), .B2(new_n817), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n808), .A2(new_n202), .ZN(new_n871));
  INV_X1    g0671(.A(G132), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n794), .A2(new_n219), .B1(new_n801), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n868), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n493), .B1(new_n274), .B2(new_n794), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT98), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n808), .A2(new_n265), .ZN(new_n879));
  INV_X1    g0679(.A(G294), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n805), .A2(new_n550), .B1(new_n797), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n801), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n879), .B(new_n881), .C1(G311), .C2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n876), .A2(new_n877), .ZN(new_n884));
  AOI22_X1  g0684(.A1(G283), .A2(new_n812), .B1(new_n815), .B2(G116), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n883), .A2(new_n884), .A3(new_n832), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n875), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n860), .B(new_n863), .C1(new_n887), .C2(new_n781), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n855), .B2(new_n779), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n859), .A2(new_n889), .ZN(G384));
  NOR2_X1   g0690(.A1(new_n769), .A2(new_n302), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n750), .B1(KEYINPUT105), .B2(KEYINPUT31), .ZN(new_n892));
  NOR2_X1   g0692(.A1(KEYINPUT105), .A2(KEYINPUT31), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n749), .A2(new_n715), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n752), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n408), .A2(new_n716), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n409), .B(new_n898), .C1(new_n421), .C2(new_n408), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n427), .A2(new_n897), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n849), .A2(new_n850), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT100), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n899), .A2(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n444), .A2(new_n447), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT16), .B1(new_n906), .B2(new_n498), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n490), .B1(new_n505), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n713), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n520), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n461), .A2(new_n518), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n512), .A2(new_n908), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n910), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n506), .A2(new_n512), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n506), .A2(new_n909), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT37), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n913), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT102), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n912), .A2(new_n921), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT38), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT102), .A4(KEYINPUT38), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n905), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT40), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT106), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT106), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n930), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n917), .A2(new_n918), .A3(new_n913), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT37), .ZN(new_n938));
  INV_X1    g0738(.A(new_n918), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n920), .A2(new_n938), .B1(new_n520), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n922), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n905), .A2(KEYINPUT40), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n936), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n546), .A2(new_n896), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n739), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT38), .B1(new_n912), .B2(new_n921), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n923), .B2(new_n922), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n951), .B2(new_n928), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n942), .A2(KEYINPUT39), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT104), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n429), .A2(new_n715), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n929), .A2(KEYINPUT39), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n942), .A2(KEYINPUT39), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT104), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n954), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n678), .A2(new_n909), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n543), .A2(new_n715), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n754), .B2(new_n855), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n899), .A2(new_n900), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n961), .B1(new_n966), .B2(new_n929), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n764), .B(new_n546), .C1(new_n754), .C2(new_n756), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n688), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n891), .B1(new_n948), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n971), .B2(new_n948), .ZN(new_n973));
  INV_X1    g0773(.A(new_n613), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT35), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT35), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n975), .A2(G116), .A3(new_n217), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT36), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n736), .A2(new_n224), .A3(new_n438), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n248), .B(KEYINPUT101), .ZN(new_n980));
  OAI211_X1 g0780(.A(G1), .B(new_n768), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(new_n978), .A3(new_n981), .ZN(G367));
  NAND2_X1  g0782(.A1(new_n623), .A2(new_n715), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n697), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n703), .A2(new_n715), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n719), .A2(new_n727), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT108), .Z(new_n988));
  NAND3_X1  g0788(.A1(new_n723), .A2(new_n725), .A3(new_n730), .ZN(new_n989));
  INV_X1    g0789(.A(new_n986), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n989), .A2(KEYINPUT42), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT42), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n625), .B1(new_n984), .B2(new_n720), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n716), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n991), .A2(new_n992), .A3(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n673), .A2(new_n716), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n694), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n692), .B2(new_n999), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n988), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n987), .B(KEYINPUT108), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(new_n1002), .A3(new_n998), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1005), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n734), .B(KEYINPUT41), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n731), .A2(new_n986), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT45), .Z(new_n1014));
  NOR2_X1   g0814(.A1(new_n731), .A2(new_n986), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT44), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n728), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n719), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n718), .A2(G330), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(KEYINPUT109), .A3(new_n989), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n727), .A2(new_n730), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1024), .B(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1014), .A2(new_n1016), .A3(new_n728), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1019), .A2(new_n1027), .A3(new_n765), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1012), .B1(new_n1029), .B2(new_n765), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1008), .B(new_n1011), .C1(new_n1030), .C2(new_n773), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1001), .A2(new_n839), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n784), .A2(new_n243), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n782), .B1(new_n537), .B2(new_n211), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n775), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n808), .A2(new_n565), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1036), .B(new_n446), .C1(G311), .C2(new_n806), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G303), .A2(new_n824), .B1(new_n882), .B2(G317), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G294), .A2(new_n812), .B1(new_n815), .B2(G283), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n794), .A2(new_n280), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1040), .A2(KEYINPUT46), .B1(G107), .B2(new_n818), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1040), .A2(KEYINPUT46), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT110), .Z(new_n1044));
  NAND2_X1  g0844(.A1(new_n882), .A2(G137), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n865), .B2(new_n805), .C1(new_n821), .C2(new_n811), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n493), .B1(G68), .B2(new_n818), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n808), .A2(new_n224), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G50), .B2(new_n815), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n825), .A2(new_n827), .B1(new_n824), .B2(G150), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1042), .A2(new_n1044), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT47), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1035), .B1(new_n1053), .B2(new_n781), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1032), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1031), .A2(new_n1055), .ZN(G387));
  NAND2_X1  g0856(.A1(new_n240), .A2(G45), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT111), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n531), .A2(new_n219), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT50), .Z(new_n1060));
  INV_X1    g0860(.A(new_n733), .ZN(new_n1061));
  AOI211_X1 g0861(.A(G45), .B(new_n1061), .C1(G68), .C2(G77), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n784), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(G107), .B2(new_n211), .C1(new_n733), .C2(new_n787), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n782), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n367), .A2(new_n811), .B1(new_n202), .B2(new_n814), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT113), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n797), .A2(new_n219), .B1(new_n808), .B2(new_n565), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1069), .B(new_n783), .C1(G159), .C2(new_n806), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n655), .A2(new_n818), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n794), .A2(new_n224), .B1(new_n801), .B2(new_n370), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT112), .Z(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G116), .A2(new_n809), .B1(new_n882), .B2(G326), .ZN(new_n1075));
  INV_X1    g0875(.A(G283), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n794), .A2(new_n880), .B1(new_n817), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G311), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n805), .A2(new_n798), .B1(new_n811), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(G317), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n797), .A2(new_n1080), .B1(new_n814), .B2(new_n550), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1077), .B1(new_n1082), .B2(KEYINPUT48), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(KEYINPUT48), .B2(new_n1082), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT49), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n783), .B(new_n1075), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1074), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT114), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n836), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1089), .B2(new_n1088), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1066), .A2(new_n775), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n727), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n780), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1027), .B2(new_n773), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1027), .A2(new_n765), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n774), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1027), .A2(new_n765), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(G393));
  INV_X1    g0899(.A(new_n1028), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n773), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n728), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n990), .A2(new_n780), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n782), .B1(new_n565), .B2(new_n211), .C1(new_n784), .C2(new_n247), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n775), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n815), .A2(new_n531), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n818), .A2(G77), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n219), .C2(new_n811), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT115), .Z(new_n1110));
  INV_X1    g0910(.A(G159), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n805), .A2(new_n370), .B1(new_n797), .B2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT51), .Z(new_n1113));
  AOI21_X1  g0913(.A(new_n879), .B1(G68), .B2(new_n827), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n865), .B2(new_n801), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1110), .A2(new_n783), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n805), .A2(new_n1080), .B1(new_n797), .B2(new_n1078), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT52), .Z(new_n1118));
  OAI22_X1  g0918(.A1(new_n811), .A2(new_n550), .B1(new_n817), .B2(new_n280), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT116), .Z(new_n1120));
  AOI22_X1  g0920(.A1(G294), .A2(new_n815), .B1(new_n882), .B2(G322), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n831), .C1(new_n1076), .C2(new_n794), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n264), .A4(new_n1122), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1106), .B1(new_n1124), .B2(new_n781), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1103), .B1(new_n1104), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1096), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n774), .A3(new_n1029), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(G390));
  AND3_X1   g0929(.A1(new_n896), .A2(G330), .A3(new_n904), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n955), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n707), .A2(new_n716), .A3(new_n855), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n962), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n964), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n954), .A2(new_n959), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n715), .B1(new_n761), .B2(new_n762), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n962), .B1(new_n1137), .B2(new_n855), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1131), .B(new_n942), .C1(new_n1138), .C2(new_n965), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1130), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n958), .B1(new_n956), .B2(new_n957), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1142), .A2(new_n1143), .B1(new_n955), .B2(new_n966), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n753), .A2(new_n855), .A3(new_n964), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n1139), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1141), .A2(new_n1146), .A3(new_n773), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n778), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n860), .B1(new_n367), .B2(new_n861), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n814), .A2(new_n565), .B1(new_n801), .B2(new_n880), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n871), .B(new_n1150), .C1(G87), .C2(new_n827), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n274), .A2(new_n811), .B1(new_n797), .B2(new_n280), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G283), .B2(new_n806), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n493), .A3(new_n1108), .A4(new_n1153), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  INV_X1    g0957(.A(G137), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n805), .A2(new_n1157), .B1(new_n811), .B2(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n797), .A2(new_n872), .B1(new_n808), .B2(new_n219), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  INV_X1    g0961(.A(G125), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n814), .A2(new_n1161), .B1(new_n801), .B2(new_n1162), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n493), .A2(new_n1159), .A3(new_n1160), .A4(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n794), .A2(new_n370), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT53), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(new_n1111), .C2(new_n817), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1155), .A2(new_n1156), .A3(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1148), .B(new_n1149), .C1(new_n836), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1147), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n546), .A2(G330), .A3(new_n896), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n969), .A2(new_n688), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT117), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n739), .B(new_n854), .C1(new_n752), .C2(new_n895), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1145), .B(new_n1138), .C1(new_n1176), .C2(new_n964), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n964), .B1(new_n753), .B2(new_n855), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(new_n1130), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1177), .B1(new_n1179), .B2(new_n963), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n969), .A2(new_n688), .A3(new_n1172), .A4(KEYINPUT117), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1175), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1141), .A2(new_n1146), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n774), .B(new_n1183), .C1(new_n1184), .C2(KEYINPUT118), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(KEYINPUT118), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1171), .B1(new_n1185), .B2(new_n1186), .ZN(G378));
  NAND3_X1  g0987(.A1(new_n936), .A2(G330), .A3(new_n943), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n375), .A2(new_n909), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n386), .B(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n960), .A2(new_n967), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n960), .B2(new_n967), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1188), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1193), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n968), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n943), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n739), .B(new_n1199), .C1(new_n933), .C2(new_n935), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n960), .A2(new_n967), .A3(new_n1193), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1196), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1197), .A2(new_n778), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n775), .B1(G50), .B2(new_n862), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n258), .A2(new_n342), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT120), .ZN(new_n1207));
  INV_X1    g1007(.A(G124), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n808), .A2(new_n821), .B1(new_n801), .B2(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n805), .A2(new_n1162), .B1(new_n811), .B2(new_n872), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1161), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n827), .A2(new_n1211), .B1(new_n815), .B2(G137), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1157), .B2(new_n797), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1210), .B(new_n1213), .C1(G150), .C2(new_n818), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1207), .B(new_n1209), .C1(new_n1215), .C2(KEYINPUT59), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(KEYINPUT59), .B2(new_n1215), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G107), .A2(new_n824), .B1(new_n882), .B2(G283), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n565), .B2(new_n811), .C1(new_n280), .C2(new_n805), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n809), .A2(new_n825), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n202), .B2(new_n817), .C1(new_n224), .C2(new_n794), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n342), .B(new_n783), .C1(new_n537), .C2(new_n814), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1207), .B(new_n219), .C1(new_n446), .C2(G41), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1217), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1205), .B1(new_n1227), .B2(new_n781), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1203), .A2(new_n773), .B1(new_n1204), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1175), .A2(new_n1181), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1183), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1203), .A2(KEYINPUT57), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n774), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1232), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1229), .B1(new_n1234), .B2(new_n1235), .ZN(G375));
  OAI211_X1 g1036(.A(new_n1230), .B(new_n1177), .C1(new_n963), .C2(new_n1179), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1012), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1175), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n565), .A2(new_n794), .B1(new_n797), .B2(new_n1076), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1048), .B(new_n1241), .C1(G294), .C2(new_n806), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n811), .A2(new_n280), .B1(new_n814), .B2(new_n274), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G303), .B2(new_n882), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1242), .A2(new_n493), .A3(new_n1071), .A4(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT121), .B1(new_n1220), .B2(new_n446), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n805), .A2(new_n872), .B1(new_n797), .B2(new_n1158), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G50), .B2(new_n818), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1220), .A2(new_n446), .A3(KEYINPUT121), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G159), .A2(new_n827), .B1(new_n812), .B2(new_n1211), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G150), .A2(new_n815), .B1(new_n882), .B2(G128), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1246), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n781), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1254), .B(new_n775), .C1(G68), .C2(new_n862), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n965), .B2(new_n778), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1180), .B2(new_n773), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1240), .A2(new_n1257), .ZN(G381));
  OR2_X1    g1058(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G378), .B1(G375), .B2(KEYINPUT122), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1262), .A2(G387), .A3(G381), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT123), .ZN(G407));
  INV_X1    g1065(.A(G213), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1261), .B2(new_n714), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G407), .A2(new_n1267), .ZN(G409));
  AND3_X1   g1068(.A1(new_n1031), .A2(new_n1055), .A3(G390), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G390), .B1(new_n1031), .B2(new_n1055), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(G393), .B(G396), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1271), .ZN(new_n1273));
  INV_X1    g1073(.A(G390), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1011), .A2(new_n1008), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1029), .A2(new_n765), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1238), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1277), .B2(new_n1101), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1055), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1274), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1031), .A2(new_n1055), .A3(G390), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1273), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1272), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1266), .A2(G343), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1239), .A2(KEYINPUT60), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1237), .A2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n774), .B1(new_n1237), .B2(new_n1286), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1257), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G384), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G384), .B(new_n1257), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G378), .B(new_n1229), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT118), .B1(new_n1295), .B2(new_n1239), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1183), .A2(new_n774), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1184), .A2(KEYINPUT118), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1170), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1203), .A2(new_n1238), .A3(new_n1232), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1229), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1285), .B(new_n1293), .C1(new_n1294), .C2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT62), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1294), .A2(new_n1303), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1285), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1293), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1305), .A2(new_n1311), .A3(KEYINPUT126), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1285), .A2(G2897), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1293), .B(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1313), .B(new_n1317), .C1(new_n1311), .C2(KEYINPUT126), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1284), .B1(new_n1312), .B2(new_n1318), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1304), .A2(KEYINPUT124), .A3(KEYINPUT63), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT124), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT63), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1309), .B2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1320), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1315), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1293), .B(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1285), .B1(new_n1294), .B2(new_n1303), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1283), .B(new_n1313), .C1(new_n1326), .C2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT125), .B1(new_n1324), .B2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT124), .B1(new_n1304), .B2(KEYINPUT63), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1309), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1317), .A2(new_n1313), .A3(new_n1329), .A4(new_n1283), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT125), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1335), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1319), .B1(new_n1332), .B2(new_n1338), .ZN(G405));
  INV_X1    g1139(.A(G375), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1293), .B1(new_n1340), .B2(G378), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1308), .A2(G375), .A3(new_n1300), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1343), .A2(KEYINPUT127), .A3(new_n1294), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1294), .A2(KEYINPUT127), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1341), .A2(new_n1345), .A3(new_n1342), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1347), .B(new_n1284), .ZN(G402));
endmodule


