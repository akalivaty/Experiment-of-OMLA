//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G127gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G134gat), .ZN(new_n206));
  INV_X1    g005(.A(G134gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G127gat), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT72), .B1(new_n205), .B2(G134gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT73), .B1(new_n207), .B2(G127gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT72), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(new_n207), .A3(G127gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(new_n205), .A3(G134gat), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n210), .A2(new_n211), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n204), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT74), .A3(new_n216), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT70), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT26), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT26), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n227), .A2(new_n222), .A3(new_n223), .A4(KEYINPUT70), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT71), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT27), .B(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT28), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT27), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n234), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  OR3_X1    g039(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT68), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n236), .B1(KEYINPUT68), .B2(new_n240), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n235), .B1(new_n243), .B2(KEYINPUT28), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT71), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n245), .A3(new_n230), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n232), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT23), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(new_n222), .A3(new_n223), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n226), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n254), .A3(new_n226), .ZN(new_n255));
  NAND3_X1  g054(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n257), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n234), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT24), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n230), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n258), .A2(new_n259), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n253), .A2(new_n255), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n256), .B(KEYINPUT67), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT68), .B(G183gat), .Z(new_n267));
  OAI211_X1 g066(.A(new_n266), .B(new_n262), .C1(G190gat), .C2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n226), .B(KEYINPUT66), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n251), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n264), .A2(new_n265), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n221), .B1(new_n247), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n264), .A2(new_n265), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OR3_X1    g074(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n276));
  INV_X1    g075(.A(new_n220), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT74), .B1(new_n204), .B2(new_n216), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n232), .A2(new_n244), .A3(new_n246), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G227gat), .ZN(new_n283));
  INV_X1    g082(.A(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT34), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n282), .A2(new_n286), .B1(KEYINPUT78), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n281), .A3(new_n285), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT32), .ZN(new_n291));
  XOR2_X1   g090(.A(G15gat), .B(G43gat), .Z(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(KEYINPUT75), .B(KEYINPUT76), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n296), .A2(KEYINPUT33), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT33), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(new_n291), .A3(new_n296), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n287), .A2(KEYINPUT78), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n300), .A2(new_n291), .A3(KEYINPUT77), .A4(new_n296), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n303), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n289), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n304), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n288), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT36), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT36), .B1(new_n309), .B2(new_n313), .ZN(new_n315));
  XNOR2_X1  g114(.A(G141gat), .B(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G155gat), .ZN(new_n318));
  INV_X1    g117(.A(G162gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(KEYINPUT2), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n321), .B(new_n320), .C1(new_n316), .C2(KEYINPUT2), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n327), .B(new_n276), .C1(new_n277), .C2(new_n278), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT4), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n221), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT84), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n324), .A2(new_n325), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n279), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT84), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n328), .A2(new_n337), .A3(KEYINPUT4), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(KEYINPUT83), .Z(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n332), .A2(new_n336), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n221), .A2(new_n327), .ZN(new_n343));
  INV_X1    g142(.A(new_n328), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT5), .ZN(new_n346));
  INV_X1    g145(.A(new_n340), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n335), .A2(new_n334), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n221), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n329), .B2(new_n331), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n342), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT0), .ZN(new_n353));
  XNOR2_X1  g152(.A(G57gat), .B(G85gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n351), .B2(new_n356), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n351), .A2(new_n356), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT80), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n275), .A2(new_n280), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G197gat), .B(G204gat), .Z(new_n372));
  NAND2_X1  g171(.A1(G211gat), .A2(G218gat), .ZN(new_n373));
  XOR2_X1   g172(.A(KEYINPUT79), .B(KEYINPUT22), .Z(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G211gat), .ZN(new_n376));
  INV_X1    g175(.A(G218gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n373), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n373), .B(new_n378), .C1(new_n374), .C2(new_n372), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n247), .A2(new_n271), .ZN(new_n383));
  INV_X1    g182(.A(new_n367), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n383), .A2(KEYINPUT81), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n368), .B2(new_n367), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n371), .B(new_n382), .C1(new_n385), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n382), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n383), .A2(new_n384), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n370), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G8gat), .B(G36gat), .Z(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT82), .ZN(new_n393));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n388), .A2(new_n391), .ZN(new_n399));
  INV_X1    g198(.A(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n388), .A2(KEYINPUT30), .A3(new_n391), .A4(new_n395), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n334), .A2(new_n369), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT3), .B1(new_n382), .B2(new_n369), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n407), .B(new_n408), .C1(new_n409), .C2(new_n327), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n381), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n369), .B(new_n413), .C1(new_n382), .C2(KEYINPUT86), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n333), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n415), .A2(new_n326), .B1(new_n389), .B2(new_n406), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n410), .B(new_n411), .C1(new_n416), .C2(new_n408), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT87), .ZN(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT31), .B(G50gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n405), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n421), .ZN(new_n424));
  AOI211_X1 g223(.A(KEYINPUT88), .B(new_n424), .C1(new_n417), .C2(KEYINPUT87), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n410), .B1(new_n416), .B2(new_n408), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G22gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n417), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n422), .B2(new_n425), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n365), .A2(new_n404), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n314), .A2(new_n315), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n400), .B1(new_n399), .B2(KEYINPUT37), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n371), .B(new_n389), .C1(new_n385), .C2(new_n387), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n382), .B1(new_n370), .B2(new_n390), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(KEYINPUT37), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT38), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n396), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n435), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n399), .A2(KEYINPUT37), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(new_n444), .B2(KEYINPUT38), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n351), .A2(KEYINPUT91), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n342), .B(new_n448), .C1(new_n346), .C2(new_n350), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n356), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT92), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n355), .B1(new_n351), .B2(KEYINPUT91), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n449), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n446), .B1(new_n455), .B2(new_n362), .ZN(new_n456));
  AOI211_X1 g255(.A(KEYINPUT93), .B(new_n361), .C1(new_n451), .C2(new_n454), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n359), .B(new_n445), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n338), .A2(new_n336), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n347), .B1(new_n459), .B2(new_n332), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n343), .A2(new_n344), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT39), .B1(new_n461), .B2(new_n340), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT89), .B(KEYINPUT39), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n355), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n463), .A2(new_n355), .A3(new_n465), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n403), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n450), .A2(KEYINPUT92), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n453), .B1(new_n452), .B2(new_n449), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n431), .A2(new_n432), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n434), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n359), .B1(new_n456), .B2(new_n457), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n309), .B2(new_n313), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n403), .A2(KEYINPUT35), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n309), .A2(new_n313), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n431), .A2(new_n432), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n403), .B1(new_n359), .B2(new_n364), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G92gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT101), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT101), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G92gat), .ZN(new_n495));
  INV_X1    g294(.A(G85gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT7), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(G85gat), .A3(G92gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT8), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G99gat), .B(G106gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n497), .A2(new_n502), .A3(new_n506), .A4(new_n504), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT102), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n497), .A2(new_n504), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT102), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n506), .A4(new_n502), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT96), .B(G50gat), .Z(new_n516));
  INV_X1    g315(.A(G43gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT95), .B(G43gat), .ZN(new_n519));
  INV_X1    g318(.A(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT15), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n517), .A2(new_n520), .ZN(new_n523));
  NOR2_X1   g322(.A1(G43gat), .A2(G50gat), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT15), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n525), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(KEYINPUT94), .B2(new_n527), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(KEYINPUT94), .B2(new_n527), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n525), .B1(new_n533), .B2(new_n526), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n515), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G190gat), .B(G218gat), .Z(new_n539));
  AND3_X1   g338(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n540), .B1(new_n535), .B2(new_n514), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT103), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT104), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n538), .A2(new_n541), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(new_n539), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT104), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n544), .A2(new_n552), .A3(new_n547), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n550), .B(new_n539), .Z(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n544), .B2(new_n547), .ZN(new_n556));
  INV_X1    g355(.A(new_n547), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT104), .B(new_n557), .C1(new_n542), .C2(new_n543), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n555), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G57gat), .B(G64gat), .Z(new_n561));
  OR2_X1    g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n563), .B(new_n562), .C1(new_n568), .C2(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G127gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G15gat), .B(G22gat), .ZN(new_n576));
  INV_X1    g375(.A(G1gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT16), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(G1gat), .B2(new_n576), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n580), .A2(G8gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(G8gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(new_n570), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n575), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n318), .ZN(new_n589));
  XOR2_X1   g388(.A(G183gat), .B(G211gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n587), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n510), .A2(new_n570), .A3(new_n513), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n509), .A2(new_n569), .A3(new_n567), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n505), .A2(KEYINPUT105), .A3(new_n507), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT105), .B1(new_n505), .B2(new_n507), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT10), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n594), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n570), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n514), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT106), .B1(new_n607), .B2(new_n600), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT106), .ZN(new_n609));
  AOI211_X1 g408(.A(new_n609), .B(new_n601), .C1(new_n604), .C2(new_n606), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n602), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(new_n600), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n602), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n560), .A2(new_n593), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT107), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G197gat), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT11), .B(G169gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(new_n535), .B2(new_n583), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n531), .A2(new_n534), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n584), .A2(new_n632), .A3(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n535), .A2(new_n583), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT13), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT99), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n583), .B(KEYINPUT97), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n536), .B2(new_n537), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n636), .A3(new_n634), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT18), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n641), .A2(KEYINPUT18), .A3(new_n636), .A4(new_n634), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n629), .B1(new_n639), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n638), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n629), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n649), .A2(new_n650), .A3(new_n644), .A4(new_n645), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n623), .A2(new_n624), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n491), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n365), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g457(.A(KEYINPUT108), .B(KEYINPUT16), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G8gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n403), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n655), .ZN(new_n664));
  OAI21_X1  g463(.A(G8gat), .B1(new_n664), .B2(new_n404), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(G1325gat));
  INV_X1    g466(.A(new_n485), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n664), .A2(G15gat), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n315), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT36), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n664), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n655), .A2(new_n477), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  AOI21_X1  g477(.A(new_n560), .B1(new_n480), .B2(new_n490), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n653), .A2(new_n593), .A3(new_n619), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(G29gat), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n656), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n479), .A2(new_n434), .B1(new_n484), .B2(new_n489), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(new_n560), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n554), .A2(new_n559), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n491), .A2(KEYINPUT44), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n680), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691), .B2(new_n365), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n684), .A2(new_n692), .ZN(G1328gat));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694));
  AOI21_X1  g493(.A(G36gat), .B1(new_n694), .B2(KEYINPUT46), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n681), .A2(new_n403), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(KEYINPUT46), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n691), .B2(new_n404), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1329gat));
  NAND4_X1  g499(.A1(new_n687), .A2(new_n689), .A3(new_n672), .A4(new_n680), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n519), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n668), .A2(new_n519), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n679), .A2(new_n680), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n702), .A2(KEYINPUT111), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n704), .B(KEYINPUT112), .Z(new_n707));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n701), .B2(new_n519), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n705), .B1(new_n710), .B2(new_n711), .ZN(G1330gat));
  NAND4_X1  g511(.A1(new_n687), .A2(new_n689), .A3(new_n477), .A4(new_n680), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n516), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n486), .A2(new_n516), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n681), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT48), .Z(G1331gat));
  NAND4_X1  g517(.A1(new_n560), .A2(new_n653), .A3(new_n593), .A4(new_n619), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n686), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n656), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n403), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT113), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n686), .A2(new_n719), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT114), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n727), .B(new_n728), .Z(G1333gat));
  NAND2_X1  g528(.A1(new_n720), .A2(new_n672), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n668), .A2(G71gat), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(G71gat), .B1(new_n720), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n720), .A2(new_n477), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n652), .A2(new_n593), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n620), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n690), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n365), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n491), .A2(new_n688), .A3(new_n736), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n679), .B2(new_n736), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n656), .A2(new_n496), .A3(new_n619), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(G1336gat));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n404), .A2(new_n620), .A3(G92gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n743), .B2(new_n744), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n687), .A2(new_n689), .A3(new_n403), .A4(new_n738), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n493), .A2(new_n495), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI211_X1 g555(.A(new_n560), .B(new_n737), .C1(new_n480), .C2(new_n490), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n742), .B1(new_n757), .B2(KEYINPUT115), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n759), .A3(KEYINPUT51), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n760), .A3(new_n749), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n754), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n748), .B(new_n756), .C1(new_n762), .C2(new_n755), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n755), .B1(new_n761), .B2(new_n754), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT116), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(G1337gat));
  OAI21_X1  g566(.A(G99gat), .B1(new_n739), .B2(new_n673), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n668), .A2(G99gat), .A3(new_n620), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n745), .B2(new_n769), .ZN(G1338gat));
  NAND4_X1  g569(.A1(new_n687), .A2(new_n689), .A3(new_n477), .A4(new_n738), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(KEYINPUT53), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n743), .A2(new_n744), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n486), .A2(G106gat), .A3(new_n620), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n758), .A2(new_n760), .A3(new_n776), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT53), .B1(new_n780), .B2(new_n772), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1339gat));
  INV_X1    g581(.A(G113gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n617), .A2(new_n609), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n607), .A2(KEYINPUT106), .A3(new_n600), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n607), .B2(new_n600), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n604), .A2(new_n601), .A3(new_n606), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n614), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n618), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT54), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n617), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n615), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n652), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n636), .B1(new_n641), .B2(new_n634), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n635), .A2(new_n637), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n628), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n802), .A2(KEYINPUT118), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(KEYINPUT118), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n651), .A2(new_n803), .A3(new_n619), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n688), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n651), .A2(new_n803), .A3(new_n804), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n807), .A2(new_n688), .A3(new_n798), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n592), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n621), .A2(new_n652), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n477), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n656), .A2(new_n404), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n668), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n783), .B1(new_n814), .B2(new_n652), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT119), .Z(new_n816));
  AOI21_X1  g615(.A(new_n365), .B1(new_n809), .B2(new_n810), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n817), .A2(new_n404), .A3(new_n482), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n783), .A3(new_n652), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(G1340gat));
  AOI21_X1  g619(.A(G120gat), .B1(new_n818), .B2(new_n619), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n619), .A2(G120gat), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n814), .B2(new_n822), .ZN(G1341gat));
  INV_X1    g622(.A(new_n814), .ZN(new_n824));
  OAI21_X1  g623(.A(G127gat), .B1(new_n824), .B2(new_n592), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n818), .A2(new_n205), .A3(new_n593), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1342gat));
  OAI21_X1  g626(.A(G134gat), .B1(new_n824), .B2(new_n560), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n560), .A2(new_n403), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n817), .A2(new_n207), .A3(new_n482), .A4(new_n829), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n828), .A2(new_n831), .A3(new_n832), .ZN(G1343gat));
  NOR2_X1   g632(.A1(new_n672), .A2(new_n812), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n809), .A2(new_n810), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n477), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n836), .B2(KEYINPUT57), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n787), .A2(new_n790), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n793), .ZN(new_n840));
  AOI211_X1 g639(.A(KEYINPUT120), .B(KEYINPUT55), .C1(new_n787), .C2(new_n790), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n792), .B(KEYINPUT121), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n652), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n797), .A2(KEYINPUT120), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n838), .A3(new_n793), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT121), .B1(new_n846), .B2(new_n792), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n805), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT122), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n805), .C1(new_n843), .C2(new_n847), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n560), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n808), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n593), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n810), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n477), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n837), .B1(new_n856), .B2(KEYINPUT57), .ZN(new_n857));
  INV_X1    g656(.A(G141gat), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n653), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n817), .A2(new_n477), .A3(new_n673), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n403), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n652), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n858), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n865), .B(new_n866), .Z(G1344gat));
  INV_X1    g666(.A(G148gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n862), .A2(new_n868), .A3(new_n619), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n486), .A2(KEYINPUT57), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n623), .A2(new_n624), .A3(new_n652), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n854), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n836), .A2(KEYINPUT57), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n619), .A3(new_n834), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n870), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT59), .B(new_n868), .C1(new_n857), .C2(new_n619), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n869), .B1(new_n877), .B2(new_n878), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n318), .A3(new_n593), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n857), .A2(new_n593), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n318), .ZN(G1346gat));
  AND2_X1   g681(.A1(new_n857), .A2(new_n688), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n829), .A2(new_n319), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n883), .A2(new_n319), .B1(new_n861), .B2(new_n884), .ZN(G1347gat));
  NAND2_X1  g684(.A1(new_n365), .A2(new_n403), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n668), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n811), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n222), .A3(new_n653), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n656), .B1(new_n809), .B2(new_n810), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n668), .A2(new_n477), .A3(new_n404), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n652), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n889), .B1(new_n222), .B2(new_n894), .ZN(G1348gat));
  AOI21_X1  g694(.A(G176gat), .B1(new_n893), .B2(new_n619), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n811), .A2(G176gat), .A3(new_n619), .A4(new_n887), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n897), .A2(KEYINPUT124), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(KEYINPUT124), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(G1349gat));
  OAI21_X1  g699(.A(new_n267), .B1(new_n888), .B2(new_n592), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n593), .A2(new_n233), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n892), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n888), .B2(new_n560), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT61), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n893), .A2(new_n234), .A3(new_n688), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1351gat));
  NOR2_X1   g707(.A1(new_n672), .A2(new_n886), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n875), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(G197gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n910), .A2(new_n911), .A3(new_n653), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n672), .A2(new_n486), .A3(new_n404), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n890), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n652), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n912), .A2(new_n915), .ZN(G1352gat));
  NOR2_X1   g715(.A1(new_n620), .A2(G204gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n890), .A2(new_n913), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT125), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n890), .A2(new_n913), .A3(new_n920), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT62), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n873), .A2(new_n619), .A3(new_n874), .A4(new_n909), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G204gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n923), .A2(KEYINPUT126), .A3(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n376), .A3(new_n593), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n873), .A2(new_n593), .A3(new_n874), .A4(new_n909), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n932), .B2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT127), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n937), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n910), .B2(new_n560), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n914), .A2(new_n377), .A3(new_n688), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1355gat));
endmodule


