//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n593, new_n595, new_n596, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1117, new_n1118;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n453), .B2(G2106), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n463), .A2(new_n465), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT69), .Z(new_n476));
  NAND2_X1  g051(.A1(new_n464), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n465), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(G162));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n482));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n461), .B2(new_n462), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(KEYINPUT71), .A3(new_n484), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n487), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n482), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n496), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT71), .B1(new_n488), .B2(new_n484), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n487), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(KEYINPUT72), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  XOR2_X1   g092(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G89), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n509), .A2(new_n523), .B1(new_n511), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G168));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n509), .A2(new_n527), .B1(new_n511), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n515), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n529), .A2(new_n531), .A3(KEYINPUT74), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT74), .B1(new_n529), .B2(new_n531), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G171));
  XOR2_X1   g109(.A(KEYINPUT75), .B(G81), .Z(new_n535));
  INV_X1    g110(.A(G43), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n509), .A2(new_n535), .B1(new_n511), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n515), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  INV_X1    g120(.A(G53), .ZN(new_n546));
  OR3_X1    g121(.A1(new_n511), .A2(KEYINPUT9), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT9), .B1(new_n511), .B2(new_n546), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n507), .A2(new_n508), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n547), .A2(new_n548), .B1(G91), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT5), .B(G543), .Z(new_n552));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n554), .A2(KEYINPUT76), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(KEYINPUT76), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G171), .ZN(G301));
  OR2_X1    g133(.A1(new_n522), .A2(new_n525), .ZN(G286));
  INV_X1    g134(.A(G166), .ZN(G303));
  OAI21_X1  g135(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n561));
  INV_X1    g136(.A(G49), .ZN(new_n562));
  INV_X1    g137(.A(G87), .ZN(new_n563));
  OAI221_X1 g138(.A(new_n561), .B1(new_n511), .B2(new_n562), .C1(new_n563), .C2(new_n509), .ZN(G288));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G61), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n552), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n507), .A2(G543), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n567), .A2(G651), .B1(new_n568), .B2(G48), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n549), .A2(G86), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G305));
  XOR2_X1   g146(.A(KEYINPUT77), .B(G85), .Z(new_n572));
  INV_X1    g147(.A(G47), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n509), .A2(new_n572), .B1(new_n511), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n515), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G290));
  INV_X1    g153(.A(G868), .ZN(new_n579));
  NOR2_X1   g154(.A1(G301), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n549), .A2(G92), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT10), .Z(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n552), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n568), .B2(G54), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n580), .B1(new_n579), .B2(new_n587), .ZN(G321));
  XOR2_X1   g163(.A(G321), .B(KEYINPUT78), .Z(G284));
  NAND2_X1  g164(.A1(G299), .A2(new_n579), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n579), .B2(G168), .ZN(G297));
  OAI21_X1  g166(.A(new_n590), .B1(new_n579), .B2(G168), .ZN(G280));
  INV_X1    g167(.A(G559), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n587), .B1(new_n593), .B2(G860), .ZN(G148));
  NAND2_X1  g169(.A1(new_n587), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G868), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g172(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n598));
  XNOR2_X1  g173(.A(G323), .B(new_n598), .ZN(G282));
  NAND2_X1  g174(.A1(new_n464), .A2(G135), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n474), .A2(G123), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n465), .A2(G111), .ZN(new_n602));
  OAI21_X1  g177(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n600), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT81), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(G2096), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(G2096), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n488), .A2(new_n466), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT80), .B(G2100), .Z(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n610), .B(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n607), .A2(new_n608), .A3(new_n613), .ZN(G156));
  XNOR2_X1  g189(.A(G2427), .B(G2438), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2430), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(KEYINPUT14), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G1341), .B(G1348), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n620), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G2451), .B(G2454), .Z(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G14), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n624), .A2(new_n627), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(G401));
  XOR2_X1   g206(.A(G2072), .B(G2078), .Z(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT83), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT17), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT84), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n638), .B(new_n640), .C1(new_n637), .C2(new_n633), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n633), .A2(new_n635), .A3(new_n639), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT18), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n636), .A2(new_n639), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n641), .B(new_n643), .C1(new_n634), .C2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT85), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(G1971), .B(G1976), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT87), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n657), .B(new_n658), .Z(new_n659));
  NOR3_X1   g234(.A1(new_n650), .A2(new_n653), .A3(new_n656), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n655), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1981), .B(G1986), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G229));
  INV_X1    g242(.A(G16), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G24), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n577), .B2(new_n668), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT89), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n464), .A2(G131), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n474), .A2(G119), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n465), .A2(G107), .ZN(new_n675));
  OAI21_X1  g250(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  MUX2_X1   g252(.A(G25), .B(new_n677), .S(G29), .Z(new_n678));
  XOR2_X1   g253(.A(KEYINPUT35), .B(G1991), .Z(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT88), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n668), .A2(G23), .ZN(new_n682));
  OR2_X1    g257(.A1(G288), .A2(KEYINPUT90), .ZN(new_n683));
  NAND2_X1  g258(.A1(G288), .A2(KEYINPUT90), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n682), .B1(new_n685), .B2(new_n668), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT33), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n668), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n668), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n688), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n672), .B(new_n681), .C1(new_n696), .C2(KEYINPUT34), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(KEYINPUT34), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n699), .A2(KEYINPUT36), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(KEYINPUT36), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n700), .ZN(new_n703));
  NOR2_X1   g278(.A1(G5), .A2(G16), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G171), .B2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT97), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1961), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G27), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G164), .B2(new_n708), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G2078), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n712));
  INV_X1    g287(.A(G34), .ZN(new_n713));
  AOI21_X1  g288(.A(G29), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G160), .B2(new_n708), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G2084), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT93), .Z(new_n718));
  NAND3_X1  g293(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n464), .A2(G139), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(KEYINPUT92), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(KEYINPUT92), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  OAI22_X1  g300(.A1(new_n723), .A2(new_n724), .B1(new_n465), .B2(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G33), .B(new_n726), .S(G29), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2072), .ZN(new_n728));
  NOR4_X1   g303(.A1(new_n707), .A2(new_n711), .A3(new_n718), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n708), .A2(G32), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n474), .A2(G129), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT94), .Z(new_n732));
  AND2_X1   g307(.A1(new_n466), .A2(G105), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT26), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n733), .B(new_n735), .C1(G141), .C2(new_n464), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(new_n708), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT27), .ZN(new_n740));
  INV_X1    g315(.A(G1996), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G35), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G162), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT29), .B(G2090), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n668), .A2(G20), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT23), .Z(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G299), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1956), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G168), .A2(G16), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(KEYINPUT95), .C1(G16), .C2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT95), .B2(new_n752), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT96), .B(G1966), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n708), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n464), .A2(G140), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n474), .A2(G128), .ZN(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(new_n708), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2067), .ZN(new_n766));
  NOR2_X1   g341(.A1(G4), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n587), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G1348), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n716), .A2(G2084), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n605), .A2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G28), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT30), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(KEYINPUT30), .ZN(new_n776));
  OR2_X1    g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  NAND2_X1  g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g354(.A1(new_n772), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n668), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n540), .B2(new_n668), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1341), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n768), .B2(G1348), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n756), .A2(new_n771), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n744), .A2(new_n745), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n742), .A2(new_n751), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n702), .A2(new_n703), .A3(new_n729), .A4(new_n787), .ZN(G150));
  INV_X1    g363(.A(G150), .ZN(G311));
  NAND2_X1  g364(.A1(new_n587), .A2(G559), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT38), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT98), .B(G93), .Z(new_n792));
  INV_X1    g367(.A(G55), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n509), .A2(new_n792), .B1(new_n511), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(new_n515), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n540), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n540), .A2(new_n797), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n791), .B(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT39), .ZN(new_n803));
  INV_X1    g378(.A(G860), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(KEYINPUT39), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n797), .A2(new_n804), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT37), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(G145));
  XOR2_X1   g384(.A(KEYINPUT102), .B(G37), .Z(new_n810));
  INV_X1    g385(.A(KEYINPUT100), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n726), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT99), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(new_n764), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n677), .B(new_n610), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n502), .A2(new_n503), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n737), .B(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(G130), .A2(new_n474), .B1(new_n464), .B2(G142), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT101), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n820), .A2(new_n465), .A3(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n465), .B2(G118), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n818), .B(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n816), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n605), .B(G160), .ZN(new_n827));
  XNOR2_X1  g402(.A(G162), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n816), .A2(new_n825), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n826), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n810), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(G395));
  OAI21_X1  g409(.A(new_n579), .B1(new_n794), .B2(new_n796), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n587), .A2(G299), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n587), .A2(G299), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(KEYINPUT104), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT104), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n587), .A2(new_n839), .A3(G299), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(KEYINPUT41), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n836), .A2(new_n842), .A3(new_n837), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n595), .B(new_n801), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n838), .A2(new_n840), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n685), .B(G305), .ZN(new_n852));
  XOR2_X1   g427(.A(G166), .B(new_n577), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n835), .B1(new_n855), .B2(new_n579), .ZN(G295));
  OAI21_X1  g431(.A(new_n835), .B1(new_n855), .B2(new_n579), .ZN(G331));
  NAND2_X1  g432(.A1(G301), .A2(G168), .ZN(new_n858));
  NAND2_X1  g433(.A1(G171), .A2(G286), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n801), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n836), .A2(new_n837), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT41), .B1(new_n838), .B2(new_n840), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT108), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n800), .B1(new_n858), .B2(new_n859), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(KEYINPUT107), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n861), .B2(KEYINPUT107), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n848), .ZN(new_n870));
  INV_X1    g445(.A(new_n865), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n871), .A2(new_n872), .A3(new_n861), .A4(new_n863), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n866), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n854), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n860), .A2(new_n801), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(new_n867), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n848), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n854), .B(new_n879), .C1(new_n869), .C2(new_n844), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n880), .A2(new_n810), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT43), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n841), .B(new_n843), .C1(new_n887), .C2(new_n868), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n854), .B1(new_n888), .B2(new_n879), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n883), .B(KEYINPUT44), .C1(new_n885), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n876), .A2(new_n881), .A3(new_n884), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n885), .B1(new_n889), .B2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT109), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n899));
  AOI211_X1 g474(.A(new_n899), .B(KEYINPUT44), .C1(new_n894), .C2(new_n895), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n893), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g478(.A(KEYINPUT110), .B(new_n893), .C1(new_n898), .C2(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(G397));
  XNOR2_X1  g480(.A(new_n737), .B(new_n741), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n763), .B(G2067), .Z(new_n907));
  AND2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n677), .B(new_n679), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G1384), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n490), .B2(new_n498), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n577), .B(G1986), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT111), .ZN(new_n921));
  INV_X1    g496(.A(G2084), .ZN(new_n922));
  AOI21_X1  g497(.A(G1384), .B1(new_n502), .B2(new_n503), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n915), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G1384), .B1(new_n499), .B2(new_n504), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT50), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n922), .B(new_n925), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n915), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n923), .B2(KEYINPUT45), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n913), .A2(G1384), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n499), .B2(new_n504), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n755), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(G8), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT119), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT118), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(G286), .B2(G8), .ZN(new_n940));
  INV_X1    g515(.A(G8), .ZN(new_n941));
  NOR3_X1   g516(.A1(G168), .A2(KEYINPUT118), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n936), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n935), .B1(new_n942), .B2(new_n940), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n938), .A2(new_n944), .A3(KEYINPUT51), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n683), .A2(new_n684), .A3(G1976), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n941), .B1(new_n929), .B2(new_n923), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT52), .ZN(new_n950));
  INV_X1    g525(.A(G1976), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT52), .B1(G288), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT114), .B(G86), .Z(new_n954));
  OAI21_X1  g529(.A(new_n569), .B1(new_n509), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G1981), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT113), .B(G1981), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n569), .A2(new_n570), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n948), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n959), .B2(new_n960), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n950), .B(new_n953), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G303), .A2(G8), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT55), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n969), .A2(G2090), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n817), .A2(new_n931), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n929), .B(new_n971), .C1(new_n926), .C2(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n691), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n941), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n965), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n936), .B(new_n943), .C1(new_n937), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n926), .A2(new_n927), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n929), .C1(new_n923), .C2(new_n924), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n973), .B1(new_n979), .B2(G2090), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G8), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n967), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n946), .A2(new_n975), .A3(new_n977), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n972), .B2(G2078), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1961), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n969), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT120), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n930), .A2(new_n933), .ZN(new_n990));
  INV_X1    g565(.A(G2078), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n490), .A2(new_n498), .A3(new_n482), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT72), .B1(new_n502), .B2(new_n503), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n931), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n915), .B1(new_n912), .B2(new_n913), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n989), .A3(new_n996), .A4(new_n991), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT53), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n988), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT121), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(KEYINPUT121), .B(new_n988), .C1(new_n992), .C2(new_n998), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n986), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G301), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n991), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1006));
  INV_X1    g581(.A(new_n467), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n471), .B(new_n1006), .C1(new_n1007), .C2(KEYINPUT122), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(KEYINPUT122), .B2(new_n1007), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(new_n914), .A3(new_n971), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n985), .A2(new_n988), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1005), .B1(new_n1011), .B2(G171), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n983), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1011), .A2(G171), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1002), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n995), .A2(new_n991), .A3(new_n996), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT120), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(KEYINPUT53), .A3(new_n997), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT121), .B1(new_n1018), .B2(new_n988), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n985), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1014), .B1(new_n1020), .B2(G171), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT123), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1021), .A2(new_n1022), .A3(KEYINPUT54), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1014), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n1003), .B2(G301), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT123), .B1(new_n1025), .B2(new_n1005), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1013), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT124), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT124), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n1013), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT61), .ZN(new_n1031));
  INV_X1    g606(.A(G1956), .ZN(new_n1032));
  INV_X1    g607(.A(new_n972), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT56), .B(G2072), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1032), .A2(new_n979), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(G299), .B(KEYINPUT57), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1031), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1038), .B(new_n1039), .Z(new_n1040));
  INV_X1    g615(.A(new_n587), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(KEYINPUT60), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n929), .A2(new_n923), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G2067), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n969), .B2(new_n770), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT58), .B(G1341), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n972), .B2(G1996), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n540), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1051));
  OAI21_X1  g626(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1045), .B(new_n587), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1040), .B(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1036), .B(KEYINPUT116), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(new_n1035), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1045), .A2(new_n1041), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1039), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1028), .A2(new_n1030), .A3(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n974), .A2(new_n968), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n936), .A2(G286), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(new_n975), .A3(KEYINPUT63), .A4(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n975), .A2(new_n982), .A3(new_n1064), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(KEYINPUT63), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n974), .A2(new_n968), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n965), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G288), .A2(G1976), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n963), .B2(new_n964), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n958), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1069), .B1(new_n1072), .B2(new_n948), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT62), .B1(new_n946), .B2(new_n977), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n975), .A2(new_n982), .ZN(new_n1076));
  NOR4_X1   g651(.A1(new_n1075), .A2(new_n1076), .A3(G301), .A4(new_n1003), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(KEYINPUT125), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n946), .A2(KEYINPUT62), .A3(new_n977), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1077), .B2(KEYINPUT125), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1074), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n921), .B1(new_n1062), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n916), .A2(new_n741), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT46), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n738), .A2(new_n907), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n918), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(new_n1088), .B(KEYINPUT47), .Z(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n763), .A2(G2067), .ZN(new_n1091));
  INV_X1    g666(.A(new_n679), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n677), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n908), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(new_n918), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT48), .ZN(new_n1096));
  OR3_X1    g671(.A1(new_n918), .A2(G1986), .A3(G290), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n910), .A2(new_n916), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1097), .A2(new_n1096), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1090), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT126), .B1(new_n1084), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1074), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1076), .A2(new_n1003), .A3(G301), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1075), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1080), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1105), .B1(new_n1110), .B2(new_n1078), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1027), .A2(KEYINPUT124), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1030), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1104), .B(new_n1101), .C1(new_n1113), .C2(new_n921), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1103), .A2(new_n1114), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g690(.A(G319), .B1(new_n629), .B2(new_n630), .ZN(new_n1117));
  NOR3_X1   g691(.A1(G229), .A2(G227), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g692(.A1(new_n832), .A2(new_n896), .A3(new_n1118), .ZN(G225));
  INV_X1    g693(.A(G225), .ZN(G308));
endmodule


