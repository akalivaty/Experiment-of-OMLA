//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G244), .ZN(new_n213));
  AOI22_X1  g0013(.A1(new_n213), .A2(G77), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n206), .C2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G68), .B2(G238), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n205), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n212), .B(new_n226), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n227), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT71), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n228), .A2(G1), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT71), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n202), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n203), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n228), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT70), .B(G58), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT8), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(KEYINPUT8), .B2(G58), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n264), .A2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n262), .B1(new_n263), .B2(new_n265), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n261), .B1(new_n271), .B2(new_n253), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n256), .A2(G13), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n202), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(G1), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n215), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(G274), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT68), .B(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OR3_X1    g0086(.A1(new_n282), .A2(new_n286), .A3(KEYINPUT69), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G222), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G223), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n292), .B(new_n293), .C1(G77), .C2(new_n288), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT69), .B1(new_n282), .B2(new_n286), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n287), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(G179), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n276), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n272), .A2(KEYINPUT9), .A3(new_n275), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT9), .B1(new_n272), .B2(new_n275), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n296), .A2(G200), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n303), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n310), .A2(new_n306), .A3(new_n301), .A4(new_n308), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n300), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT16), .ZN(new_n314));
  INV_X1    g0114(.A(G159), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT77), .B1(new_n265), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G20), .A2(G33), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT77), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(G159), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n201), .B1(new_n266), .B2(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n228), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  OR2_X1    g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n228), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n325), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n323), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n314), .B1(new_n322), .B2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT7), .B1(new_n334), .B2(new_n228), .ZN(new_n335));
  INV_X1    g0135(.A(new_n329), .ZN(new_n336));
  OAI21_X1  g0136(.A(G68), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G58), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT70), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G58), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n341), .A3(G68), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n231), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(G20), .B1(new_n316), .B2(new_n319), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n337), .A2(new_n344), .A3(KEYINPUT16), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n331), .A2(new_n345), .A3(new_n253), .ZN(new_n346));
  MUX2_X1   g0146(.A(new_n260), .B(new_n273), .S(new_n268), .Z(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OR2_X1    g0148(.A1(G223), .A2(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n215), .A2(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n332), .C2(new_n333), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G87), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n293), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  INV_X1    g0155(.A(new_n286), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n278), .A2(G232), .A3(new_n280), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n278), .B1(new_n351), .B2(new_n352), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n360), .A2(new_n286), .A3(new_n357), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n361), .B2(G169), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n348), .A2(KEYINPUT18), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT78), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n346), .A2(new_n347), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(new_n362), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n362), .B1(new_n346), .B2(new_n347), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT78), .A3(KEYINPUT18), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT79), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n360), .A2(new_n286), .ZN(new_n374));
  AOI21_X1  g0174(.A(G200), .B1(new_n374), .B2(new_n358), .ZN(new_n375));
  NOR4_X1   g0175(.A1(new_n360), .A2(new_n286), .A3(new_n357), .A4(G190), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n307), .A3(new_n358), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(KEYINPUT79), .C1(new_n361), .C2(G200), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n368), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n368), .A3(KEYINPUT17), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n372), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n254), .A2(new_n273), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n387), .A2(new_n323), .A3(new_n256), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n317), .A2(G50), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n389), .B(KEYINPUT75), .ZN(new_n390));
  INV_X1    g0190(.A(G77), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n390), .B1(new_n228), .B2(G68), .C1(new_n391), .C2(new_n270), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n253), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT11), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT11), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n395), .A3(new_n253), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n388), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n279), .A2(new_n323), .A3(G13), .A4(G20), .ZN(new_n398));
  XOR2_X1   g0198(.A(new_n398), .B(KEYINPUT12), .Z(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n215), .A2(new_n290), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n288), .B(new_n403), .C1(G232), .C2(new_n290), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n278), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n286), .ZN(new_n407));
  INV_X1    g0207(.A(G238), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n281), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n402), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  NOR4_X1   g0211(.A1(new_n406), .A2(KEYINPUT13), .A3(new_n286), .A4(new_n409), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT14), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(G169), .C1(new_n411), .C2(new_n412), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n407), .A2(new_n410), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n419));
  INV_X1    g0219(.A(new_n412), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(KEYINPUT74), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(new_n422), .A3(KEYINPUT13), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n355), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n401), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n411), .A2(new_n412), .A3(new_n422), .ZN(new_n426));
  INV_X1    g0226(.A(new_n423), .ZN(new_n427));
  OAI21_X1  g0227(.A(G190), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n419), .B2(new_n420), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n428), .A2(new_n431), .A3(new_n400), .A4(new_n397), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n313), .B(new_n386), .C1(KEYINPUT76), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(KEYINPUT76), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n254), .A2(new_n273), .A3(G77), .A4(new_n257), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n273), .A2(G77), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT73), .ZN(new_n438));
  XOR2_X1   g0238(.A(KEYINPUT15), .B(G87), .Z(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n317), .B(KEYINPUT72), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT8), .B(G58), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n270), .A2(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(G20), .B2(G77), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n436), .B(new_n438), .C1(new_n444), .C2(new_n254), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n408), .A2(G1698), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(G232), .B2(G1698), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n278), .B1(new_n447), .B2(new_n288), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(G107), .B2(new_n288), .ZN(new_n449));
  INV_X1    g0249(.A(new_n281), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n213), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n451), .A3(new_n356), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n452), .A2(G200), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n445), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n307), .B2(new_n452), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n298), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n445), .B(new_n456), .C1(G179), .C2(new_n452), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n435), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n434), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT81), .B(G97), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT6), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n460), .A2(new_n206), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n207), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n464), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n228), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n317), .A2(G77), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT82), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n205), .A2(KEYINPUT81), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G97), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n476), .A3(new_n206), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n468), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n462), .A2(new_n464), .B1(new_n207), .B2(new_n466), .ZN(new_n479));
  OAI21_X1  g0279(.A(G20), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT82), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n471), .ZN(new_n482));
  OAI21_X1  g0282(.A(G107), .B1(new_n335), .B2(new_n336), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n473), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n253), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n273), .A2(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n254), .B(new_n273), .C1(G1), .C2(new_n264), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(G97), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G45), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G1), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G274), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n496), .A2(G257), .A3(new_n278), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n290), .A2(G244), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n334), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT83), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n221), .A2(new_n290), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n288), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n500), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n288), .A2(G244), .A3(new_n290), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n498), .B(new_n499), .C1(new_n511), .C2(new_n293), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G179), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n293), .ZN(new_n514));
  INV_X1    g0314(.A(new_n498), .ZN(new_n515));
  INV_X1    g0315(.A(new_n499), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G169), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n490), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n499), .B1(new_n511), .B2(new_n293), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(new_n307), .A3(new_n515), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n512), .B2(G200), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n485), .A3(new_n489), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n288), .A2(new_n525), .A3(new_n228), .A4(G87), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n228), .B(G87), .C1(new_n332), .C2(new_n333), .ZN(new_n527));
  XOR2_X1   g0327(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT23), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n228), .B2(G107), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n531), .A2(new_n532), .B1(new_n269), .B2(G116), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n526), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n526), .A2(new_n529), .A3(KEYINPUT24), .A4(new_n533), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n253), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n279), .A2(new_n206), .A3(G13), .A4(G20), .ZN(new_n539));
  XOR2_X1   g0339(.A(new_n539), .B(KEYINPUT25), .Z(new_n540));
  AND2_X1   g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n221), .A2(new_n290), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n223), .A2(G1698), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n332), .C2(new_n333), .ZN(new_n544));
  INV_X1    g0344(.A(G294), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n264), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n496), .A2(new_n278), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n293), .A2(new_n546), .B1(new_n547), .B2(G264), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(G190), .A3(new_n515), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n488), .A2(G107), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n515), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n541), .A2(new_n549), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n439), .A2(new_n273), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n288), .A2(new_n228), .A3(G68), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n474), .A2(new_n476), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n270), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n460), .A2(G87), .A3(G107), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n405), .A2(new_n556), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(G20), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n555), .B(new_n558), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n554), .B1(new_n562), .B2(new_n253), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n488), .A2(new_n439), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n408), .A2(new_n290), .ZN(new_n565));
  INV_X1    g0365(.A(G244), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G1698), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n567), .C1(new_n332), .C2(new_n333), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G116), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n278), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n279), .A2(G45), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n278), .A2(new_n571), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n572), .A2(new_n221), .B1(new_n497), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n563), .A2(new_n564), .B1(new_n575), .B2(new_n298), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n355), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n487), .A2(new_n220), .ZN(new_n578));
  AOI211_X1 g0378(.A(new_n554), .B(new_n578), .C1(new_n562), .C2(new_n253), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n570), .A2(new_n573), .A3(new_n307), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n575), .B2(G200), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n576), .A2(new_n577), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n520), .A2(new_n524), .A3(new_n553), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n496), .A2(G270), .A3(new_n278), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n223), .A2(new_n290), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n216), .A2(G1698), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n278), .B1(new_n589), .B2(new_n288), .ZN(new_n590));
  INV_X1    g0390(.A(G303), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n324), .A2(new_n591), .A3(new_n325), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT84), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n290), .A2(G264), .ZN(new_n594));
  NOR2_X1   g0394(.A1(G257), .A2(G1698), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(new_n332), .B2(new_n333), .ZN(new_n596));
  AND4_X1   g0396(.A1(KEYINPUT84), .A2(new_n596), .A3(new_n293), .A4(new_n592), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n515), .B(new_n586), .C1(new_n593), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G169), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n274), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n487), .B2(new_n600), .ZN(new_n602));
  AOI21_X1  g0402(.A(G20), .B1(G33), .B2(G283), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n557), .B2(G33), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(G20), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n253), .A2(KEYINPUT85), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT85), .B1(new_n253), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n604), .B(KEYINPUT20), .C1(new_n606), .C2(new_n607), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n602), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT21), .B1(new_n599), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n602), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n253), .A2(new_n605), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n253), .A2(KEYINPUT85), .A3(new_n605), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT20), .B1(new_n619), .B2(new_n604), .ZN(new_n620));
  INV_X1    g0420(.A(new_n611), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(G169), .A4(new_n598), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n613), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n596), .A2(new_n293), .A3(new_n592), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n590), .A2(KEYINPUT84), .A3(new_n592), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n498), .B(new_n585), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n622), .A2(G179), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n598), .A2(G200), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n632), .B(new_n612), .C1(new_n307), .C2(new_n598), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n538), .A2(new_n550), .A3(new_n540), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n551), .A2(new_n298), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n548), .A2(new_n355), .A3(new_n515), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n625), .A2(new_n631), .A3(new_n633), .A4(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n459), .A2(new_n584), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT87), .ZN(G372));
  AND2_X1   g0441(.A1(new_n625), .A2(new_n631), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n583), .B1(new_n642), .B2(new_n637), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n576), .A2(new_n577), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n579), .A2(new_n581), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n644), .B1(new_n520), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n485), .A2(new_n489), .B1(new_n513), .B2(new_n518), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n582), .A3(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n645), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n459), .B1(new_n643), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT88), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n307), .B1(new_n421), .B2(new_n423), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n655), .A2(new_n401), .A3(new_n430), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n425), .B1(new_n656), .B2(new_n457), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n380), .A2(new_n368), .A3(KEYINPUT17), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT17), .B1(new_n380), .B2(new_n368), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(KEYINPUT90), .B(new_n425), .C1(new_n656), .C2(new_n457), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n364), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n370), .A2(KEYINPUT18), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT89), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT89), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n369), .B2(new_n364), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n309), .A2(new_n312), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n300), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n654), .A2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n625), .A2(new_n631), .ZN(new_n677));
  INV_X1    g0477(.A(G13), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n678), .A2(G1), .A3(G20), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT27), .ZN(new_n680));
  OR3_X1    g0480(.A1(new_n679), .A2(KEYINPUT91), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G213), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n679), .B2(new_n680), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT91), .B1(new_n679), .B2(new_n680), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n612), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n677), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n642), .A2(new_n633), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n637), .A2(new_n687), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n634), .A2(new_n687), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n553), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n695), .B1(new_n697), .B2(new_n637), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n637), .ZN(new_n700));
  NOR4_X1   g0500(.A1(new_n642), .A2(new_n697), .A3(new_n700), .A4(new_n687), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n695), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(G399));
  NAND2_X1  g0503(.A1(new_n559), .A2(new_n600), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n210), .A2(new_n285), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n704), .A2(new_n706), .B1(new_n232), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(new_n645), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n648), .B2(new_n650), .ZN(new_n710));
  INV_X1    g0510(.A(new_n490), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n649), .B1(new_n711), .B2(new_n523), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n625), .A2(new_n631), .A3(new_n637), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(new_n553), .A4(new_n582), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n687), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n584), .A2(new_n639), .A3(new_n688), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n546), .A2(new_n293), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n496), .A2(G264), .A3(new_n278), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n571), .A2(new_n497), .ZN(new_n723));
  INV_X1    g0523(.A(new_n572), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(G250), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n568), .A2(new_n569), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n293), .ZN(new_n727));
  AND4_X1   g0527(.A1(new_n721), .A2(new_n722), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n630), .A2(new_n512), .A3(new_n728), .A4(G179), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n521), .A2(G179), .A3(new_n515), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(KEYINPUT30), .A3(new_n630), .A4(new_n728), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n515), .B1(new_n521), .B2(new_n548), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(new_n355), .A3(new_n575), .A4(new_n598), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n731), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n687), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT31), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(new_n739), .A3(new_n687), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n719), .B1(new_n720), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n718), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n708), .B1(new_n745), .B2(G1), .ZN(G364));
  OR2_X1    g0546(.A1(new_n692), .A2(G330), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n678), .A2(G20), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G45), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(G1), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n705), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n747), .A2(new_n693), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n228), .A2(G179), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G329), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n228), .A2(new_n355), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n764), .A2(new_n429), .A3(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  OAI221_X1 g0567(.A(new_n761), .B1(new_n591), .B2(new_n762), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n763), .A2(G190), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G200), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n288), .B(new_n768), .C1(G322), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n769), .A2(new_n429), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G326), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n757), .A2(new_n307), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT98), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G283), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n307), .A2(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n228), .B1(new_n781), .B2(new_n355), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n763), .A2(new_n758), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT97), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n787), .A2(G294), .B1(new_n794), .B2(G311), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n771), .A2(new_n773), .A3(new_n780), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n759), .A2(new_n315), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n787), .A2(G97), .B1(KEYINPUT32), .B2(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n794), .A2(G77), .B1(G68), .B2(new_n765), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n798), .A2(KEYINPUT32), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n779), .B2(G107), .ZN(new_n802));
  INV_X1    g0602(.A(new_n770), .ZN(new_n803));
  INV_X1    g0603(.A(new_n266), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n288), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G50), .B2(new_n772), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n799), .A2(new_n800), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n762), .A2(new_n220), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n796), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n227), .B1(G20), .B2(new_n298), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT95), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT95), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G13), .A2(G33), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n228), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT94), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT96), .ZN(new_n819));
  NAND3_X1  g0619(.A1(G355), .A2(new_n288), .A3(new_n210), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n247), .A2(new_n491), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n334), .A2(new_n210), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT93), .Z(new_n823));
  INV_X1    g0623(.A(new_n284), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n232), .B2(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n820), .B1(G116), .B2(new_n210), .C1(new_n821), .C2(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n809), .A2(new_n813), .B1(new_n819), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n817), .B(KEYINPUT100), .Z(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n692), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n756), .B1(new_n755), .B2(new_n830), .ZN(G396));
  NOR2_X1   g0631(.A1(new_n813), .A2(new_n815), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n391), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n457), .A2(new_n687), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n445), .A2(new_n687), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n455), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(new_n836), .B2(new_n457), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n755), .B1(new_n838), .B2(new_n815), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n334), .B1(new_n759), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n772), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n842), .A2(new_n591), .B1(new_n206), .B2(new_n762), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(G294), .C2(new_n770), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n765), .A2(G283), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n779), .A2(G87), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n787), .A2(G97), .B1(new_n794), .B2(G116), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G150), .A2(new_n765), .B1(new_n770), .B2(G143), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n850), .B2(new_n842), .C1(new_n793), .C2(new_n315), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT34), .Z(new_n852));
  AOI211_X1 g0652(.A(new_n334), .B(new_n852), .C1(G132), .C2(new_n760), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n779), .A2(G68), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(new_n202), .C2(new_n762), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n786), .A2(new_n804), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n848), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT101), .Z(new_n858));
  OAI211_X1 g0658(.A(new_n833), .B(new_n839), .C1(new_n858), .C2(new_n814), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n715), .B(new_n838), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(new_n743), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n755), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n859), .A2(new_n862), .ZN(G384));
  INV_X1    g0663(.A(new_n685), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n672), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n348), .A2(new_n864), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n372), .B2(new_n385), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n348), .B1(new_n363), .B2(new_n864), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n381), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n381), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n662), .B1(new_n667), .B2(new_n670), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n872), .B2(new_n873), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n381), .A2(new_n871), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT102), .B1(new_n880), .B2(new_n870), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n877), .A2(new_n868), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n866), .B(new_n876), .C1(new_n882), .C2(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n869), .B2(new_n875), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n867), .B1(new_n662), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n886), .A2(new_n874), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT39), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(G179), .B1(new_n426), .B2(new_n427), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n414), .A3(new_n416), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n401), .A3(new_n688), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n865), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n884), .A2(new_n888), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n401), .A2(new_n687), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n425), .A2(new_n432), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n892), .A2(new_n401), .A3(new_n687), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n834), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n688), .B1(new_n652), .B2(new_n643), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n902), .B2(new_n838), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n896), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n895), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n459), .A2(new_n717), .A3(new_n716), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n675), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n905), .B(new_n907), .Z(new_n908));
  NAND2_X1  g0708(.A1(new_n459), .A2(new_n742), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n884), .A2(new_n888), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n720), .A2(new_n741), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n837), .A3(new_n900), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n912), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n882), .A2(KEYINPUT38), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n888), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n913), .B1(KEYINPUT40), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n909), .B1(new_n917), .B2(new_n719), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n896), .A2(new_n919), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n879), .A2(new_n881), .ZN(new_n921));
  INV_X1    g0721(.A(new_n877), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n867), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n887), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n912), .B1(new_n924), .B2(new_n876), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n920), .B1(new_n925), .B2(new_n919), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n459), .A3(new_n911), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n918), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n908), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n279), .B2(new_n748), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n465), .A2(new_n469), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n600), .B1(new_n931), .B2(KEYINPUT35), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(new_n230), .C1(KEYINPUT35), .C2(new_n931), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n233), .A2(G77), .A3(new_n342), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(G50), .B2(new_n323), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n678), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(G367));
  NAND3_X1  g0738(.A1(new_n490), .A2(new_n519), .A3(new_n687), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT105), .Z(new_n940));
  OAI21_X1  g0740(.A(new_n712), .B1(new_n711), .B2(new_n688), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n701), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT42), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n579), .A2(new_n688), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n645), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n582), .B2(new_n945), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT103), .Z(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT104), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n942), .A2(new_n700), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n687), .B1(new_n952), .B2(new_n520), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n944), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n948), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n951), .B1(new_n950), .B2(new_n955), .C1(new_n944), .C2(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n699), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n942), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n957), .B(new_n959), .Z(new_n960));
  XOR2_X1   g0760(.A(new_n705), .B(KEYINPUT41), .Z(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n698), .B1(new_n677), .B2(new_n688), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n693), .B1(new_n701), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT106), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n699), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(new_n744), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT107), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n702), .A2(new_n942), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT44), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n702), .A2(new_n942), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT45), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(new_n958), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n967), .A2(KEYINPUT107), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n962), .B1(new_n976), .B2(new_n745), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n960), .B1(new_n977), .B2(new_n752), .ZN(new_n978));
  INV_X1    g0778(.A(new_n818), .ZN(new_n979));
  INV_X1    g0779(.A(new_n823), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n979), .B1(new_n210), .B2(new_n440), .C1(new_n980), .C2(new_n242), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n755), .B1(new_n955), .B2(new_n828), .ZN(new_n982));
  INV_X1    g0782(.A(new_n762), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(G116), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n984), .A2(new_n985), .B1(new_n772), .B2(G311), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n591), .B2(new_n803), .C1(new_n557), .C2(new_n778), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n288), .B1(new_n794), .B2(G283), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n765), .A2(G294), .B1(G317), .B2(new_n760), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(new_n985), .C2(new_n984), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(G107), .C2(new_n787), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n759), .A2(new_n850), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n786), .A2(new_n323), .B1(new_n263), .B2(new_n803), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT108), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n779), .A2(G77), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n288), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n794), .A2(G50), .B1(G143), .B2(new_n772), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n994), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n992), .B(new_n1000), .C1(G159), .C2(new_n765), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n983), .A2(new_n266), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n991), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n981), .B(new_n982), .C1(new_n1004), .C2(new_n814), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n978), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(G387));
  INV_X1    g0807(.A(new_n966), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n752), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n288), .B1(new_n842), .B2(new_n315), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n766), .A2(new_n268), .B1(new_n803), .B2(new_n202), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(G77), .C2(new_n983), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n760), .A2(G150), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n787), .A2(new_n439), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G68), .A2(new_n794), .B1(new_n779), .B2(G97), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(G283), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n786), .A2(new_n1017), .B1(new_n545), .B2(new_n762), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT111), .Z(new_n1019));
  AOI22_X1  g0819(.A1(G311), .A2(new_n765), .B1(new_n770), .B2(G317), .ZN(new_n1020));
  INV_X1    g0820(.A(G322), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n842), .C1(new_n793), .C2(new_n591), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1023), .A2(KEYINPUT48), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(KEYINPUT48), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1019), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT49), .Z(new_n1027));
  NAND2_X1  g0827(.A1(new_n760), .A2(G326), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n334), .B(new_n1028), .C1(new_n778), .C2(new_n600), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1016), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n813), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n704), .A2(new_n210), .A3(new_n288), .ZN(new_n1032));
  AOI211_X1 g0832(.A(G45), .B(new_n704), .C1(G68), .C2(G77), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT110), .Z(new_n1034));
  INV_X1    g0834(.A(new_n442), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n202), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n823), .B1(new_n239), .B2(new_n284), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1032), .B1(G107), .B2(new_n210), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n819), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n698), .A2(new_n829), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1031), .A2(new_n754), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n753), .B1(new_n1008), .B2(new_n745), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1009), .B(new_n1043), .C1(new_n1044), .C2(new_n967), .ZN(G393));
  OR2_X1    g0845(.A1(new_n942), .A2(new_n817), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n979), .B1(new_n210), .B2(new_n557), .C1(new_n980), .C2(new_n250), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n754), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n787), .A2(G77), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G150), .A2(new_n772), .B1(new_n770), .B2(G159), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1052));
  AND4_X1   g0852(.A1(new_n846), .A2(new_n1049), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n983), .A2(G68), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n334), .B1(new_n794), .B2(new_n1035), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n765), .A2(G50), .B1(G143), .B2(new_n760), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n794), .A2(G294), .B1(G303), .B2(new_n765), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n600), .B2(new_n786), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT112), .Z(new_n1060));
  OAI21_X1  g0860(.A(new_n334), .B1(new_n759), .B2(new_n1021), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G283), .B2(new_n983), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(new_n206), .C2(new_n778), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G311), .A2(new_n770), .B1(new_n772), .B2(G317), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1057), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1048), .B1(new_n813), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n974), .B2(new_n752), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n976), .B1(new_n974), .B2(new_n967), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n705), .ZN(G390));
  AND3_X1   g0870(.A1(new_n736), .A2(new_n739), .A3(new_n687), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n739), .B1(new_n736), .B2(new_n687), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n583), .A2(new_n638), .A3(new_n687), .ZN(new_n1074));
  OAI211_X1 g0874(.A(G330), .B(new_n837), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n900), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT115), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n834), .B1(new_n715), .B2(new_n837), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n911), .A2(new_n900), .A3(G330), .A4(new_n837), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1075), .A2(new_n1076), .A3(KEYINPUT115), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(KEYINPUT114), .B(new_n1080), .C1(new_n1081), .C2(new_n1077), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT114), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n903), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n675), .A2(new_n909), .A3(new_n906), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT113), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n883), .A2(new_n889), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n894), .B1(new_n903), .B2(new_n900), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n915), .A2(new_n888), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n883), .A2(new_n889), .A3(KEYINPUT113), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n893), .B1(new_n1080), .B2(new_n1076), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1081), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1095), .A2(new_n1098), .A3(new_n1081), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1090), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1095), .A2(new_n1098), .A3(new_n1081), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1081), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1089), .B(new_n1088), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n753), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n752), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n883), .A2(new_n889), .A3(new_n815), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n854), .B1(new_n545), .B2(new_n759), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT117), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G107), .A2(new_n765), .B1(new_n770), .B2(G116), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1049), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n460), .B2(new_n794), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n808), .A2(new_n288), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1115), .B1(KEYINPUT116), .B2(new_n1116), .C1(new_n1017), .C2(new_n842), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1112), .B(new_n1117), .C1(KEYINPUT116), .C2(new_n1116), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT54), .B(G143), .Z(new_n1119));
  NAND2_X1  g0919(.A1(new_n794), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n779), .A2(G50), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n760), .A2(G125), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n762), .A2(new_n263), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G132), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n803), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n786), .A2(new_n315), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n288), .B1(new_n842), .B2(new_n1129), .C1(new_n850), .C2(new_n766), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n813), .B1(new_n1118), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n832), .A2(new_n268), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1110), .A2(new_n754), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1107), .A2(new_n1109), .A3(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(KEYINPUT120), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n276), .A2(new_n864), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n313), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n313), .A2(new_n1137), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n917), .A2(new_n719), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n926), .B2(G330), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1136), .B(new_n905), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n917), .B2(new_n719), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n926), .A2(G330), .A3(new_n1146), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n905), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1150), .C1(new_n1151), .C2(KEYINPUT120), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n752), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n755), .B1(new_n1146), .B2(new_n815), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n765), .A2(G97), .B1(G283), .B2(new_n760), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n793), .B2(new_n440), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n786), .A2(new_n323), .B1(new_n600), .B2(new_n842), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT118), .Z(new_n1159));
  AOI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(G107), .C2(new_n770), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n779), .A2(new_n266), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G41), .B1(new_n983), .B2(G77), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1160), .A2(new_n334), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT58), .Z(new_n1164));
  INV_X1    g0964(.A(G124), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n264), .B1(new_n759), .B2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n787), .A2(G150), .B1(G125), .B2(new_n772), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n983), .A2(new_n1119), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n766), .B2(new_n1126), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G137), .B2(new_n794), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1167), .B(new_n1170), .C1(new_n1129), .C2(new_n803), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G41), .B(new_n1166), .C1(new_n1171), .C2(KEYINPUT59), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(KEYINPUT59), .B2(new_n1171), .C1(new_n315), .C2(new_n778), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n202), .B1(new_n332), .B2(G41), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n813), .B1(new_n1164), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n832), .A2(new_n202), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1155), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT119), .Z(new_n1179));
  NAND2_X1  g0979(.A1(new_n1154), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1089), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n1108), .C2(new_n1088), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT121), .B1(new_n1106), .B2(new_n1089), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1153), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1090), .B1(new_n1102), .B2(new_n1101), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1181), .B1(new_n1188), .B2(new_n1182), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1106), .A2(KEYINPUT121), .A3(new_n1089), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n905), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1192), .A2(KEYINPUT57), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n705), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1180), .B1(new_n1187), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(G375));
  OR2_X1    g0997(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n961), .A3(new_n1090), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1076), .A2(new_n815), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n770), .A2(G283), .B1(new_n983), .B2(G97), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n545), .B2(new_n842), .C1(new_n793), .C2(new_n206), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n288), .B1(new_n765), .B2(G116), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1014), .A2(new_n995), .A3(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(G303), .C2(new_n760), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n334), .B1(new_n765), .B2(new_n1119), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n1129), .B2(new_n759), .C1(new_n793), .C2(new_n263), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n772), .A2(G132), .B1(new_n983), .B2(G159), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1161), .B(new_n1208), .C1(new_n202), .C2(new_n786), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1207), .B(new_n1209), .C1(G137), .C2(new_n770), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n813), .B1(new_n1205), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n832), .A2(new_n323), .ZN(new_n1212));
  AND4_X1   g1012(.A1(new_n754), .A2(new_n1200), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1088), .B2(new_n752), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1199), .A2(new_n1214), .ZN(G381));
  NOR2_X1   g1015(.A1(G375), .A2(G378), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1218));
  AND4_X1   g1018(.A1(new_n1006), .A2(new_n1218), .A3(new_n1214), .A4(new_n1199), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT122), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1220), .B2(new_n1219), .ZN(G407));
  NOR2_X1   g1022(.A1(new_n682), .A2(G343), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT123), .Z(new_n1224));
  OAI211_X1 g1024(.A(G407), .B(G213), .C1(new_n1217), .C2(new_n1224), .ZN(G409));
  NAND2_X1  g1025(.A1(new_n1006), .A2(G390), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1006), .A2(G390), .ZN(new_n1227));
  XOR2_X1   g1027(.A(G393), .B(G396), .Z(new_n1228));
  AND2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1228), .A2(KEYINPUT127), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1226), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1006), .A2(new_n1230), .A3(G390), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1192), .A2(new_n752), .A3(new_n1193), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1178), .B(new_n1235), .C1(new_n1185), .C2(new_n962), .ZN(new_n1236));
  INV_X1    g1036(.A(G378), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT124), .B1(new_n1196), .B2(G378), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1194), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n753), .B(new_n1240), .C1(new_n1242), .C2(KEYINPUT57), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1180), .ZN(new_n1244));
  AND4_X1   g1044(.A1(KEYINPUT124), .A2(new_n1243), .A3(G378), .A4(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1238), .B1(new_n1239), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1223), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1198), .A2(KEYINPUT125), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT60), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1198), .A2(KEYINPUT125), .A3(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1249), .A2(new_n753), .A3(new_n1090), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1214), .ZN(new_n1253));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(KEYINPUT126), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(KEYINPUT126), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1252), .A2(KEYINPUT126), .A3(new_n1254), .A4(new_n1214), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1246), .A2(new_n1247), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1224), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1243), .A2(G378), .A3(new_n1244), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1196), .A2(KEYINPUT124), .A3(G378), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1262), .B1(new_n1267), .B2(new_n1238), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1259), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(new_n1261), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1260), .A2(new_n1261), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1257), .A2(new_n1258), .B1(G2897), .B2(new_n1223), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1262), .A2(G2897), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1273), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1272), .B1(new_n1268), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1234), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1269), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1280), .B1(new_n1283), .B2(new_n1275), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1260), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1279), .B(new_n1282), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1278), .A2(new_n1286), .ZN(G405));
  OAI21_X1  g1087(.A(new_n1267), .B1(G378), .B2(new_n1196), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1259), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1234), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1288), .A2(new_n1269), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1288), .A2(new_n1269), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1279), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(G402));
endmodule


