//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AND2_X1   g0009(.A1(G68), .A2(G238), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT66), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n210), .B(new_n212), .C1(G77), .C2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT67), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n217), .B(new_n218), .C1(new_n213), .C2(new_n214), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT64), .Z(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n209), .B(new_n221), .C1(new_n225), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(G97), .B(G107), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n248));
  OR2_X1    g0048(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n222), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G50), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n254), .B1(G50), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n203), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n223), .A2(G33), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n257), .B1(new_n258), .B2(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n256), .B1(new_n251), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT9), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n251), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n267), .B(new_n254), .C1(G50), .C2(new_n255), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n277), .A2(G223), .B1(G77), .B2(new_n275), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n276), .ZN(new_n280));
  INV_X1    g0080(.A(G222), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT68), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n281), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n270), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G274), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n270), .A2(new_n287), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(G226), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n266), .A2(new_n269), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(G200), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n248), .B(new_n249), .C1(new_n294), .C2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n285), .A2(new_n291), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n264), .A2(new_n265), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n298), .A2(G190), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n301), .A2(KEYINPUT71), .A3(KEYINPUT10), .A4(new_n295), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n298), .A2(KEYINPUT69), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n292), .B2(G179), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n292), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n304), .A2(new_n306), .A3(new_n308), .A4(new_n268), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n297), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n279), .A2(G226), .A3(new_n276), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G97), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n279), .A2(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(G232), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n311), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n270), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n289), .B1(new_n290), .B2(G238), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n317), .B1(new_n316), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g0121(.A(G200), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n321), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(G190), .A3(new_n319), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n255), .A2(G68), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT12), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(new_n329), .C1(new_n326), .C2(new_n325), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n253), .A2(G68), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n242), .A2(G20), .ZN(new_n332));
  INV_X1    g0132(.A(G77), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n332), .B1(new_n262), .B2(new_n333), .C1(new_n260), .C2(new_n202), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n251), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(KEYINPUT11), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(KEYINPUT11), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n330), .B(new_n331), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n322), .A2(new_n324), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(G169), .B1(new_n320), .B2(new_n321), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT14), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(G169), .C1(new_n320), .C2(new_n321), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n320), .A2(new_n321), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G179), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n340), .B1(new_n347), .B2(new_n338), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n277), .A2(G238), .B1(G107), .B2(new_n275), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n314), .B2(new_n280), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n270), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n289), .B1(new_n290), .B2(G244), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G200), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n253), .A2(G77), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G77), .B2(new_n255), .ZN(new_n356));
  INV_X1    g0156(.A(new_n261), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT70), .ZN(new_n359));
  OR2_X1    g0159(.A1(KEYINPUT15), .A2(G87), .ZN(new_n360));
  NAND2_X1  g0160(.A1(KEYINPUT15), .A2(G87), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(new_n359), .A3(new_n361), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n358), .B1(new_n365), .B2(new_n262), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n356), .B1(new_n366), .B2(new_n251), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n354), .B(new_n367), .C1(new_n293), .C2(new_n353), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n353), .B2(new_n307), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n351), .A2(new_n303), .A3(new_n352), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n310), .A2(new_n348), .A3(new_n368), .A4(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT7), .B1(new_n275), .B2(new_n223), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  AOI211_X1 g0174(.A(new_n374), .B(G20), .C1(new_n272), .C2(new_n274), .ZN(new_n375));
  OAI21_X1  g0175(.A(G68), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G58), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n242), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n201), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n259), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n374), .B1(new_n279), .B2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n242), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n384), .B1(new_n387), .B2(new_n381), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(new_n388), .A3(new_n251), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n261), .A2(new_n255), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n253), .B2(new_n261), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G41), .ZN(new_n393));
  OAI211_X1 g0193(.A(G1), .B(G13), .C1(new_n271), .C2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(G232), .A3(new_n286), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n288), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT74), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT73), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n272), .A2(new_n274), .A3(G223), .A4(new_n276), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n272), .A2(new_n274), .A3(G226), .A4(G1698), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n270), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT74), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n395), .A2(new_n288), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n396), .B1(new_n270), .B2(new_n402), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n406), .A2(G190), .B1(G200), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n392), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT76), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AND4_X1   g0215(.A1(new_n389), .A2(new_n408), .A3(new_n391), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n410), .B1(new_n392), .B2(new_n408), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT76), .B1(new_n419), .B2(new_n416), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n406), .A2(G179), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n407), .A2(G169), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n389), .A2(new_n391), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n418), .A2(new_n420), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n372), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n255), .A2(G97), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n251), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n252), .A2(G33), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n255), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G97), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G107), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n385), .B2(new_n386), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(G97), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(G107), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT6), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n445), .B2(new_n443), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n439), .B1(new_n449), .B2(new_n251), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n252), .B(G45), .C1(new_n393), .C2(KEYINPUT5), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n393), .A2(KEYINPUT5), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n394), .B(G257), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n272), .A2(new_n274), .A3(G244), .A4(new_n276), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT4), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n276), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n454), .B1(new_n461), .B2(new_n270), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT77), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(KEYINPUT5), .C2(new_n393), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n451), .A2(KEYINPUT77), .ZN(new_n467));
  INV_X1    g0267(.A(G274), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(KEYINPUT5), .B2(new_n393), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n394), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n462), .A2(G190), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n461), .A2(new_n270), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n472), .A2(new_n470), .A3(new_n453), .ZN(new_n473));
  INV_X1    g0273(.A(G200), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n450), .B(new_n471), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n443), .A2(new_n445), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n445), .B2(new_n239), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n477), .A2(new_n223), .B1(new_n333), .B2(new_n260), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n251), .B1(new_n478), .B2(new_n441), .ZN(new_n479));
  INV_X1    g0279(.A(new_n439), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n462), .A2(new_n303), .A3(new_n470), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n481), .B(new_n482), .C1(new_n473), .C2(G169), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT19), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n223), .B1(new_n312), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G87), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(new_n438), .A3(new_n440), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n272), .A2(new_n274), .A3(new_n223), .A4(G68), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n485), .B1(new_n262), .B2(new_n438), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n251), .ZN(new_n493));
  INV_X1    g0293(.A(new_n255), .ZN(new_n494));
  INV_X1    g0294(.A(new_n364), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n362), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n435), .A2(G87), .A3(new_n255), .A4(new_n436), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n252), .A2(G45), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G250), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n270), .A2(new_n500), .B1(new_n468), .B2(new_n499), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n272), .A2(new_n274), .A3(G238), .A4(new_n276), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n272), .A2(new_n274), .A3(G244), .A4(G1698), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G116), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n501), .B1(new_n505), .B2(new_n270), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G190), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n498), .B(new_n507), .C1(new_n506), .C2(new_n474), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n493), .B(new_n496), .C1(new_n365), .C2(new_n437), .ZN(new_n509));
  AOI211_X1 g0309(.A(new_n303), .B(new_n501), .C1(new_n270), .C2(new_n505), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(new_n270), .ZN(new_n511));
  INV_X1    g0311(.A(new_n501), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n307), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n509), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n484), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n279), .A2(G250), .A3(new_n276), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n272), .A2(new_n274), .A3(G257), .A4(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G294), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n521), .A2(new_n270), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n394), .B(G264), .C1(new_n451), .C2(new_n452), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n470), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n517), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n524), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n270), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(KEYINPUT81), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G169), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT82), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n470), .A3(new_n523), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n303), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n307), .B1(new_n525), .B2(new_n528), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT82), .B1(new_n536), .B2(new_n533), .ZN(new_n537));
  INV_X1    g0337(.A(new_n437), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G107), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT25), .B1(new_n255), .B2(G107), .ZN(new_n540));
  OR3_X1    g0340(.A1(new_n255), .A2(KEYINPUT25), .A3(G107), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n539), .A2(KEYINPUT80), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n541), .C1(new_n437), .C2(new_n440), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n440), .A2(G20), .ZN(new_n547));
  AND2_X1   g0347(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n548));
  NOR2_X1   g0348(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(G20), .A3(new_n440), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n223), .A2(G33), .A3(G116), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT79), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT79), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n550), .A2(new_n556), .A3(new_n552), .A4(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n279), .A2(new_n223), .A3(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT22), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT22), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n279), .A2(new_n560), .A3(new_n223), .A4(G87), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n555), .A2(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n251), .B1(new_n562), .B2(KEYINPUT24), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n555), .A2(new_n557), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n561), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n564), .A2(KEYINPUT24), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n546), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n535), .A2(new_n537), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n272), .A2(new_n274), .A3(G257), .A4(new_n276), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n272), .A2(new_n274), .A3(G264), .A4(G1698), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n279), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n270), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n394), .B(G270), .C1(new_n451), .C2(new_n452), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n470), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n435), .A2(G116), .A3(new_n255), .A4(new_n436), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n494), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n250), .A2(new_n222), .B1(G20), .B2(new_n577), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n459), .B(new_n223), .C1(G33), .C2(new_n438), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(KEYINPUT20), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT20), .B1(new_n579), .B2(new_n580), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n576), .B(new_n578), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n575), .A2(KEYINPUT21), .A3(G169), .A4(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n470), .A2(new_n574), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n585), .A2(new_n583), .A3(G179), .A4(new_n573), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n307), .B1(new_n585), .B2(new_n573), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT21), .B1(new_n588), .B2(new_n583), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n583), .B1(new_n575), .B2(G200), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n293), .B2(new_n575), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n525), .A2(new_n528), .A3(new_n293), .ZN(new_n594));
  INV_X1    g0394(.A(new_n532), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(G200), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n567), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n516), .A2(new_n568), .A3(new_n593), .A4(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n432), .A2(new_n599), .ZN(G372));
  INV_X1    g0400(.A(new_n309), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n341), .A2(KEYINPUT14), .B1(new_n345), .B2(G179), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n339), .B1(new_n602), .B2(new_n344), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n370), .B2(new_n369), .ZN(new_n604));
  INV_X1    g0404(.A(new_n340), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n418), .A2(new_n420), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n429), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n297), .A2(new_n302), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n475), .A2(new_n483), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT83), .B1(new_n510), .B2(new_n513), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n506), .A2(G179), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n307), .C2(new_n506), .ZN(new_n614));
  INV_X1    g0414(.A(new_n365), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n538), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n365), .A2(new_n494), .B1(new_n492), .B2(new_n251), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n611), .A2(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n508), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n610), .A2(new_n598), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n567), .B1(new_n536), .B2(new_n533), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT84), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n622), .A2(new_n623), .A3(new_n590), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n622), .B2(new_n590), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NOR4_X1   g0426(.A1(new_n618), .A2(new_n483), .A3(new_n619), .A4(KEYINPUT26), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT26), .B1(new_n483), .B2(new_n515), .ZN(new_n628));
  INV_X1    g0428(.A(new_n618), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n609), .B1(new_n432), .B2(new_n632), .ZN(G369));
  AND2_X1   g0433(.A1(new_n223), .A2(G13), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n252), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n568), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n568), .B(new_n598), .C1(new_n597), .C2(new_n641), .ZN(new_n643));
  INV_X1    g0443(.A(new_n590), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n641), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n640), .A2(new_n583), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n590), .A2(new_n592), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n647), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(G330), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n568), .A2(new_n598), .A3(new_n644), .A4(new_n641), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n622), .A2(new_n640), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(G399));
  INV_X1    g0457(.A(new_n207), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G41), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n488), .A2(G116), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G1), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n226), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n568), .A2(new_n590), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n484), .B1(new_n596), .B2(new_n597), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n620), .A3(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n483), .A2(new_n515), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n629), .B1(new_n668), .B2(KEYINPUT26), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  INV_X1    g0470(.A(new_n483), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(new_n620), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n640), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT29), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n622), .A2(new_n590), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT84), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n622), .A2(new_n590), .A3(new_n623), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n666), .A2(new_n677), .A3(new_n620), .A4(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n627), .A2(new_n630), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n640), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n675), .B1(KEYINPUT29), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n473), .A2(new_n595), .ZN(new_n683));
  INV_X1    g0483(.A(new_n506), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n575), .A2(new_n684), .A3(KEYINPUT86), .A4(new_n303), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n575), .A2(new_n303), .A3(new_n684), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT86), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n683), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n532), .A2(new_n684), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n575), .A2(new_n303), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(new_n462), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT85), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n694), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n690), .A2(new_n691), .A3(new_n462), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n689), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT87), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n640), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(KEYINPUT87), .A3(new_n702), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n649), .A2(new_n484), .A3(new_n515), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n598), .A3(new_n568), .A4(new_n641), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n682), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n664), .B1(new_n710), .B2(G1), .ZN(G364));
  AOI21_X1  g0511(.A(new_n252), .B1(new_n634), .B2(G45), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n659), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n651), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(G330), .B2(new_n650), .ZN(new_n716));
  INV_X1    g0516(.A(new_n714), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n279), .A2(G355), .A3(new_n207), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n658), .A2(new_n279), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n246), .A2(new_n463), .ZN(new_n720));
  OAI221_X1 g0520(.A(new_n719), .B1(G45), .B2(new_n227), .C1(new_n720), .C2(KEYINPUT88), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n720), .A2(KEYINPUT88), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n718), .B1(G116), .B2(new_n207), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n222), .B1(G20), .B2(new_n307), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n293), .A2(G20), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n303), .A2(new_n474), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(KEYINPUT33), .B(G317), .Z(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n474), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G283), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n275), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n731), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n735), .B(new_n739), .C1(G329), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n223), .A2(new_n293), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n736), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n744), .A2(new_n732), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n746), .A2(G303), .B1(new_n747), .B2(G326), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(G179), .A3(new_n474), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n730), .A2(new_n303), .A3(G200), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n750), .A2(G322), .B1(G311), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n223), .B1(new_n740), .B2(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G294), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n743), .A2(new_n748), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n741), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT89), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(KEYINPUT32), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT90), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n737), .A2(new_n440), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n745), .A2(new_n487), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n762), .A2(new_n763), .A3(new_n275), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n759), .A2(KEYINPUT32), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n747), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n768), .A2(new_n202), .B1(new_n733), .B2(new_n242), .ZN(new_n769));
  INV_X1    g0569(.A(new_n751), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n770), .A2(new_n333), .B1(new_n377), .B2(new_n749), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n754), .A2(G97), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(new_n761), .C2(new_n764), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n756), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n717), .B(new_n729), .C1(new_n727), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n726), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n650), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n716), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(G396));
  NOR2_X1   g0580(.A1(new_n371), .A2(new_n640), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n368), .B1(new_n367), .B2(new_n641), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n782), .B2(new_n371), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n681), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n714), .B1(new_n784), .B2(new_n709), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n709), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n727), .A2(new_n724), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n714), .B1(new_n788), .B2(G77), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT91), .ZN(new_n790));
  INV_X1    g0590(.A(new_n727), .ZN(new_n791));
  INV_X1    g0591(.A(G143), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n258), .A2(new_n733), .B1(new_n749), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n770), .A2(new_n757), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(G137), .C2(new_n747), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n279), .B1(new_n745), .B2(new_n202), .ZN(new_n798));
  INV_X1    g0598(.A(G132), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n737), .A2(new_n242), .B1(new_n741), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n798), .B(new_n800), .C1(G58), .C2(new_n754), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n796), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n275), .B1(new_n745), .B2(new_n440), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT92), .Z(new_n804));
  OAI22_X1  g0604(.A1(new_n768), .A2(new_n571), .B1(new_n737), .B2(new_n487), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n770), .A2(new_n577), .B1(new_n741), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n733), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G283), .A2(new_n809), .B1(new_n750), .B2(G294), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n804), .A2(new_n773), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n802), .A2(new_n811), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n790), .B1(new_n791), .B2(new_n812), .C1(new_n783), .C2(new_n725), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n786), .A2(new_n813), .ZN(G384));
  OAI211_X1 g0614(.A(new_n225), .B(G116), .C1(KEYINPUT35), .C2(new_n447), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(KEYINPUT35), .B2(new_n447), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT36), .ZN(new_n817));
  OR3_X1    g0617(.A1(new_n378), .A2(new_n226), .A3(new_n333), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n252), .B(G13), .C1(new_n818), .C2(new_n241), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT40), .ZN(new_n821));
  INV_X1    g0621(.A(new_n391), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n387), .A2(new_n384), .A3(new_n381), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n388), .A2(new_n251), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT93), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n388), .A2(KEYINPUT93), .A3(new_n251), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n822), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n638), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n430), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n638), .B(KEYINPUT95), .Z(new_n831));
  NAND2_X1  g0631(.A1(new_n424), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n409), .A2(new_n425), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n408), .A2(new_n389), .A3(new_n391), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT16), .B1(new_n376), .B2(new_n382), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n825), .B1(new_n837), .B2(new_n435), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(new_n383), .A3(new_n827), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n391), .ZN(new_n840));
  INV_X1    g0640(.A(new_n638), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n423), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n835), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT94), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n834), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n409), .B1(new_n828), .B2(new_n638), .ZN(new_n847));
  INV_X1    g0647(.A(new_n423), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n828), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n845), .B(KEYINPUT37), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(KEYINPUT38), .B(new_n830), .C1(new_n846), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n833), .B(new_n835), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n412), .A2(new_n417), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n832), .B1(new_n855), .B2(new_n429), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n853), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n703), .B(new_n699), .C1(new_n599), .C2(new_n640), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n338), .A2(new_n640), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n348), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n603), .A2(new_n640), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(new_n783), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n821), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n859), .A2(new_n821), .A3(new_n863), .A4(new_n783), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n830), .B1(new_n846), .B2(new_n851), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n853), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n869), .B2(new_n852), .ZN(new_n870));
  OAI21_X1  g0670(.A(G330), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n431), .A2(G330), .A3(new_n859), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n852), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n847), .B2(new_n849), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT94), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n850), .A3(new_n834), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n877), .B2(new_n830), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n864), .B1(new_n852), .B2(new_n857), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n879), .A2(new_n867), .B1(new_n880), .B2(new_n821), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n431), .A3(new_n859), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n675), .B(new_n431), .C1(KEYINPUT29), .C2(new_n681), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n609), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n883), .B(new_n885), .Z(new_n886));
  INV_X1    g0686(.A(new_n863), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n641), .B(new_n783), .C1(new_n626), .C2(new_n631), .ZN(new_n888));
  INV_X1    g0688(.A(new_n781), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n874), .B2(new_n878), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n429), .A2(new_n831), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT96), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n891), .A2(KEYINPUT96), .A3(new_n892), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n869), .B2(new_n852), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n852), .A2(new_n897), .A3(new_n857), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n603), .B(new_n641), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n886), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n252), .B2(new_n634), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n886), .A2(new_n903), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n820), .B1(new_n905), .B2(new_n906), .ZN(G367));
  NOR2_X1   g0707(.A1(new_n641), .A2(new_n498), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n629), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n620), .B2(new_n908), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT97), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n726), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n768), .A2(new_n792), .B1(new_n745), .B2(new_n377), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n753), .A2(new_n242), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n737), .A2(new_n333), .ZN(new_n915));
  OR4_X1    g0715(.A1(new_n275), .A2(new_n913), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n750), .A2(G150), .B1(G50), .B2(new_n751), .ZN(new_n917));
  INV_X1    g0717(.A(G137), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n917), .B1(new_n918), .B2(new_n741), .C1(new_n757), .C2(new_n733), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n750), .A2(G303), .B1(new_n747), .B2(G311), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n279), .B1(new_n751), .B2(G283), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n920), .B(new_n921), .C1(new_n440), .C2(new_n753), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT100), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n745), .B2(new_n577), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT46), .ZN(new_n925));
  AOI22_X1  g0725(.A1(G294), .A2(new_n809), .B1(new_n742), .B2(G317), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(KEYINPUT46), .ZN(new_n927));
  INV_X1    g0727(.A(new_n737), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(G97), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n916), .A2(new_n919), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT47), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n791), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(new_n934));
  INV_X1    g0734(.A(new_n719), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n728), .B1(new_n365), .B2(new_n207), .C1(new_n236), .C2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n912), .A2(new_n714), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n610), .B1(new_n450), .B2(new_n641), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n653), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(KEYINPUT42), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n483), .B1(new_n938), .B2(new_n568), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n939), .A2(KEYINPUT42), .B1(new_n641), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT43), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n911), .A2(new_n944), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n943), .A2(KEYINPUT98), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT98), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n911), .A2(new_n944), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n943), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n671), .A2(new_n640), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n938), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n652), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n950), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n655), .A2(new_n953), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT44), .Z(new_n958));
  INV_X1    g0758(.A(KEYINPUT45), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n655), .A2(new_n959), .A3(new_n953), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT45), .B1(new_n656), .B2(new_n952), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n646), .A2(new_n651), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n963), .A2(new_n652), .A3(new_n653), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(KEYINPUT99), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n710), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n659), .B(KEYINPUT41), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n713), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n937), .B1(new_n956), .B2(new_n968), .ZN(G387));
  AOI22_X1  g0769(.A1(new_n742), .A2(G150), .B1(new_n746), .B2(G77), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(new_n279), .A3(new_n929), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT104), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n770), .A2(new_n242), .B1(new_n261), .B2(new_n733), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT105), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n615), .A2(new_n754), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n750), .A2(G50), .B1(new_n747), .B2(G159), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n972), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n279), .B1(new_n742), .B2(G326), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n746), .A2(G294), .B1(new_n754), .B2(G283), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n747), .A2(G322), .B1(new_n751), .B2(G303), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n980), .B1(new_n806), .B2(new_n733), .C1(new_n981), .C2(new_n749), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT48), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT106), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n983), .B2(new_n982), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n978), .B1(new_n577), .B2(new_n737), .C1(new_n986), .C2(KEYINPUT49), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(KEYINPUT49), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n727), .ZN(new_n990));
  INV_X1    g0790(.A(new_n661), .ZN(new_n991));
  AOI211_X1 g0791(.A(G45), .B(new_n991), .C1(G68), .C2(G77), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(KEYINPUT102), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n261), .A2(G50), .ZN(new_n995));
  XNOR2_X1  g0795(.A(KEYINPUT103), .B(KEYINPUT50), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT102), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n719), .B1(new_n463), .B2(new_n233), .C1(new_n994), .C2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n991), .A2(new_n207), .A3(new_n279), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(G107), .B2(new_n207), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT101), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n717), .B1(new_n1004), .B2(new_n728), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n990), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n642), .A2(new_n643), .A3(new_n726), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1006), .A2(new_n1007), .B1(new_n964), .B2(new_n713), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n964), .A2(new_n682), .A3(new_n709), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n659), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT107), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n710), .A2(new_n964), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1008), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT108), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1013), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1021), .A2(KEYINPUT108), .A3(new_n1008), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1022), .ZN(G393));
  XOR2_X1   g0823(.A(new_n962), .B(new_n652), .Z(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n712), .B2(new_n1010), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n240), .A2(new_n935), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n728), .B1(new_n438), .B2(new_n207), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n714), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n768), .A2(new_n258), .B1(new_n749), .B2(new_n757), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT51), .Z(new_n1030));
  NOR2_X1   g0830(.A1(new_n753), .A2(new_n333), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n275), .B(new_n1031), .C1(G87), .C2(new_n928), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n742), .A2(G143), .B1(new_n746), .B2(G68), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n809), .A2(G50), .B1(new_n751), .B2(new_n357), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n279), .B(new_n762), .C1(G116), .C2(new_n754), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n742), .A2(G322), .B1(G294), .B2(new_n751), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n809), .A2(G303), .B1(new_n746), .B2(G283), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n750), .A2(G311), .B1(new_n747), .B2(G317), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT52), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1030), .A2(new_n1035), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1028), .B1(new_n1042), .B2(new_n727), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n952), .B2(new_n777), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n962), .A2(KEYINPUT99), .A3(new_n652), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1045), .A2(new_n659), .A3(new_n710), .A4(new_n964), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n652), .B1(new_n962), .B2(KEYINPUT99), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1025), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(G390));
  INV_X1    g0850(.A(KEYINPUT109), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT39), .B1(new_n874), .B2(new_n878), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n603), .A2(new_n641), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n781), .B1(new_n681), .B2(new_n783), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n887), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n899), .A3(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n708), .A2(G330), .A3(new_n783), .A4(new_n863), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n782), .A2(new_n371), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n781), .B1(new_n674), .B2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n858), .B(new_n1053), .C1(new_n887), .C2(new_n1059), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n865), .A2(G330), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n884), .A2(new_n609), .A3(new_n872), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n783), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n887), .B1(new_n709), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1054), .B1(new_n1066), .B2(new_n1062), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n859), .A2(G330), .A3(new_n783), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n887), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1064), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1061), .A2(new_n1063), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1051), .B1(new_n1073), .B2(new_n660), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n884), .A2(new_n609), .A3(new_n872), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1066), .A2(new_n1062), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1054), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1078), .B2(new_n1070), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1079), .B(new_n1080), .C1(new_n1081), .C2(new_n1062), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(KEYINPUT109), .A3(new_n659), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1072), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1074), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1061), .A2(new_n1063), .A3(new_n712), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n898), .A2(new_n900), .A3(new_n725), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n714), .B1(new_n788), .B2(new_n357), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT110), .Z(new_n1089));
  AOI22_X1  g0889(.A1(G294), .A2(new_n742), .B1(new_n750), .B2(G116), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n242), .B2(new_n737), .C1(new_n738), .C2(new_n768), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1091), .A2(new_n279), .A3(new_n763), .A4(new_n1031), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n770), .A2(new_n438), .B1(new_n440), .B2(new_n733), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT111), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n746), .A2(G150), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1095), .A2(KEYINPUT53), .B1(new_n757), .B2(new_n753), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(KEYINPUT53), .B2(new_n1095), .ZN(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT54), .B(G143), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n750), .A2(G132), .B1(new_n751), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n918), .B2(new_n733), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n279), .B1(new_n768), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n737), .A2(new_n202), .B1(new_n741), .B2(new_n1103), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1092), .A2(new_n1094), .B1(new_n1097), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1089), .B1(new_n1106), .B2(new_n791), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1087), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT112), .B1(new_n1086), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n713), .B(new_n1080), .C1(new_n1081), .C2(new_n1062), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT112), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1108), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1085), .A2(KEYINPUT113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT113), .B1(new_n1085), .B2(new_n1114), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(KEYINPUT118), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n268), .A2(new_n841), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n1120));
  XNOR2_X1  g0920(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n310), .B(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1122), .B(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n881), .B2(G330), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n1125), .C1(new_n866), .C2(new_n870), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n902), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT96), .B1(new_n891), .B2(new_n892), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1053), .B1(new_n1052), .B2(new_n899), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1125), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n871), .A2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n896), .A2(new_n1132), .B1(new_n1134), .B2(new_n1127), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1118), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1082), .A2(new_n1064), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n902), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1132), .A2(new_n1134), .A3(new_n896), .A4(new_n1127), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT118), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT57), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT119), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT57), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1078), .A2(new_n1070), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1075), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1144), .B(new_n659), .C1(new_n1145), .C2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n659), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1143), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1136), .A2(new_n713), .A3(new_n1140), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n799), .A2(new_n733), .B1(new_n749), .B2(new_n1101), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n746), .A2(new_n1098), .B1(new_n751), .B2(G137), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1103), .B2(new_n768), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G150), .C2(new_n754), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT59), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(G33), .A2(G41), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT114), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n737), .A2(new_n757), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(G124), .C2(new_n742), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n809), .A2(G97), .B1(new_n747), .B2(G116), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n440), .B2(new_n749), .C1(new_n365), .C2(new_n770), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n393), .B(new_n275), .C1(new_n745), .C2(new_n333), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n737), .A2(new_n377), .B1(new_n741), .B2(new_n738), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1167), .A2(new_n914), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT58), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(KEYINPUT58), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1162), .B(new_n202), .C1(G41), .C2(new_n279), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1165), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n727), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT115), .Z(new_n1176));
  OAI211_X1 g0976(.A(new_n1176), .B(new_n714), .C1(G50), .C2(new_n788), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1125), .B2(new_n724), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1153), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1152), .A2(new_n1181), .ZN(G375));
  NAND3_X1  g0982(.A1(new_n1078), .A2(new_n1075), .A3(new_n1070), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n967), .A3(new_n1072), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n863), .A2(new_n725), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT120), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(KEYINPUT120), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n714), .B1(new_n788), .B2(G68), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n733), .A2(new_n577), .B1(new_n741), .B2(new_n571), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1190), .A2(new_n279), .A3(new_n915), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n747), .A2(G294), .B1(new_n751), .B2(G107), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n750), .A2(G283), .B1(new_n746), .B2(G97), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n975), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT121), .Z(new_n1195));
  OAI22_X1  g0995(.A1(new_n768), .A2(new_n799), .B1(new_n741), .B2(new_n1101), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n275), .B(new_n1196), .C1(G58), .C2(new_n928), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n750), .A2(G137), .B1(G150), .B2(new_n751), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n809), .A2(new_n1098), .B1(new_n746), .B2(G159), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n754), .A2(G50), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1195), .A2(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1202), .A2(KEYINPUT122), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n791), .B1(new_n1202), .B2(KEYINPUT122), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1189), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1187), .A2(new_n1188), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1147), .B2(new_n713), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1184), .A2(new_n1207), .ZN(G381));
  AOI22_X1  g1008(.A1(new_n1142), .A2(new_n1141), .B1(new_n1150), .B2(KEYINPUT119), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1180), .B1(new_n1209), .B2(new_n1149), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT123), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(KEYINPUT123), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1085), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1019), .A2(new_n1022), .A3(new_n779), .ZN(new_n1215));
  OR4_X1    g1015(.A1(G384), .A2(G390), .A3(G387), .A4(G381), .ZN(new_n1216));
  OR3_X1    g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n639), .A2(G213), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT124), .Z(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G407), .B(G213), .C1(new_n1214), .C2(new_n1220), .ZN(G409));
  NAND3_X1  g1021(.A1(new_n1138), .A2(new_n1139), .A3(new_n713), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n967), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1179), .B(new_n1222), .C1(new_n1141), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1213), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(G375), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1183), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n659), .A3(new_n1072), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1183), .A2(new_n1228), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1207), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(KEYINPUT125), .B2(G384), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1232), .A2(KEYINPUT125), .A3(G384), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1227), .A2(new_n1220), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT62), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1219), .A2(G2897), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1235), .A2(new_n1236), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G378), .A2(new_n1210), .B1(new_n1213), .B2(new_n1224), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(new_n1219), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT62), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1227), .A2(new_n1247), .A3(new_n1220), .A4(new_n1237), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1239), .A2(new_n1240), .A3(new_n1246), .A4(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1049), .B(G387), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT127), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1019), .A2(new_n1022), .A3(new_n779), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n779), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT126), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT108), .B1(new_n1021), .B2(new_n1008), .ZN(new_n1257));
  OAI21_X1  g1057(.A(G396), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1215), .A3(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1251), .A2(new_n1252), .A3(new_n1255), .A4(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1255), .A2(new_n1260), .A3(new_n1252), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1250), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1252), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1249), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1238), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1262), .A2(new_n1250), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1262), .A2(new_n1250), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1264), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1227), .A2(new_n1220), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1244), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1238), .A2(new_n1267), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1268), .A2(new_n1272), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1266), .A2(new_n1276), .ZN(G405));
  NAND2_X1  g1077(.A1(G378), .A2(new_n1210), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G375), .A2(new_n1213), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1272), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1237), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1265), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(G402));
endmodule


