//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  INV_X1    g037(.A(G101), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G2104), .ZN(new_n464));
  OAI22_X1  g039(.A1(new_n461), .A2(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n459), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  OR2_X1    g044(.A1(new_n461), .A2(KEYINPUT65), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n461), .A2(KEYINPUT65), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n459), .A2(G2105), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  AND2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  OAI211_X1 g058(.A(G126), .B(G2105), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n487), .A3(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n482), .B2(new_n483), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n483), .C2(new_n482), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT67), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OR3_X1    g079(.A1(new_n503), .A2(KEYINPUT69), .A3(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(KEYINPUT66), .A3(G50), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n499), .A2(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n513));
  XOR2_X1   g088(.A(KEYINPUT68), .B(G88), .Z(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n503), .B2(new_n504), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n505), .A2(new_n515), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n508), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(new_n513), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n519), .B(new_n520), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(G168));
  XNOR2_X1  g104(.A(KEYINPUT71), .B(G52), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n508), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n504), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  AND2_X1   g111(.A1(new_n502), .A2(G56), .ZN(new_n537));
  AND2_X1   g112(.A1(G68), .A2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(G651), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n513), .A2(G81), .B1(new_n508), .B2(G43), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  AOI22_X1  g123(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n504), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n508), .A2(G53), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n513), .A2(G91), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT73), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(G299));
  XNOR2_X1  g132(.A(G171), .B(KEYINPUT74), .ZN(G301));
  INV_X1    g133(.A(G168), .ZN(G286));
  NAND2_X1  g134(.A1(new_n508), .A2(G49), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n506), .A2(new_n507), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n502), .A2(G87), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(KEYINPUT75), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n513), .B2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n560), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n499), .A2(new_n568), .A3(new_n501), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT76), .B1(new_n569), .B2(G651), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(KEYINPUT76), .A3(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n567), .A2(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n502), .A2(G86), .A3(new_n561), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT77), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n513), .A2(new_n577), .A3(G86), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n499), .B2(new_n501), .ZN(new_n580));
  AND2_X1   g155(.A1(G73), .A2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n576), .A2(new_n578), .B1(new_n582), .B2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n508), .A2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n513), .A2(G85), .B1(new_n508), .B2(G47), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n504), .B2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(new_n513), .A2(G92), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(G54), .B2(new_n508), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n504), .B1(new_n592), .B2(KEYINPUT78), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(KEYINPUT78), .B2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  MUX2_X1   g171(.A(G301), .B(new_n595), .S(new_n596), .Z(G284));
  MUX2_X1   g172(.A(G301), .B(new_n595), .S(new_n596), .Z(G321));
  NAND2_X1  g173(.A1(G299), .A2(new_n596), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n596), .B2(G168), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(new_n596), .B2(G168), .ZN(G280));
  INV_X1    g176(.A(new_n595), .ZN(new_n602));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G860), .ZN(G148));
  NOR2_X1   g179(.A1(new_n543), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n603), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n473), .A2(G135), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  INV_X1    g186(.A(G111), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G2105), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n478), .B2(G123), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G2096), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT80), .B(G2100), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n615), .A2(G2096), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n616), .A2(new_n621), .A3(new_n622), .A4(new_n623), .ZN(G156));
  INV_X1    g199(.A(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n627), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n630), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(G401));
  INV_X1    g214(.A(KEYINPUT18), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT81), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT20), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n653), .A2(new_n655), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n662), .A2(new_n658), .A3(new_n656), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n663), .C1(new_n658), .C2(new_n662), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT82), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(G229));
  MUX2_X1   g247(.A(G6), .B(G305), .S(G16), .Z(new_n673));
  XOR2_X1   g248(.A(KEYINPUT32), .B(G1981), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G22), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G166), .B2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT33), .B(G1976), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(G16), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(new_n572), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(new_n570), .ZN(new_n686));
  OAI21_X1  g261(.A(KEYINPUT84), .B1(new_n566), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n562), .A2(KEYINPUT75), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n513), .A2(new_n564), .A3(G87), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n573), .A2(new_n690), .A3(new_n691), .A4(new_n560), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n684), .B1(new_n693), .B2(new_n676), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n681), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n683), .B2(new_n694), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  MUX2_X1   g274(.A(G24), .B(G290), .S(G16), .Z(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(G1986), .Z(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n473), .A2(G131), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(G107), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G2105), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n478), .B2(G119), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(new_n702), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(KEYINPUT85), .A2(KEYINPUT36), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n478), .A2(G129), .ZN(new_n717));
  INV_X1    g292(.A(G105), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT86), .B(KEYINPUT26), .Z(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n717), .B1(new_n718), .B2(new_n464), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G141), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n472), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n702), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n702), .B2(G32), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2072), .ZN(new_n732));
  OR2_X1    g307(.A1(G29), .A2(G33), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  AOI22_X1  g310(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n736));
  INV_X1    g311(.A(G139), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n735), .B1(new_n460), .B2(new_n736), .C1(new_n472), .C2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n733), .B1(new_n738), .B2(new_n702), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n731), .B1(new_n732), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G168), .A2(new_n676), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n676), .B2(G21), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G171), .A2(new_n676), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G5), .B2(new_n676), .ZN(new_n746));
  INV_X1    g321(.A(G1961), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n740), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G164), .A2(G29), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G27), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n610), .A2(G29), .A3(new_n614), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT31), .B(G11), .Z(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n702), .B1(new_n757), .B2(G28), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT87), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(KEYINPUT87), .B1(new_n757), .B2(G28), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n762), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n729), .A2(new_n730), .B1(new_n747), .B2(new_n746), .ZN(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n765), .A2(KEYINPUT24), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(KEYINPUT24), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n702), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G160), .B2(new_n702), .ZN(new_n769));
  INV_X1    g344(.A(G2084), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n764), .B(new_n771), .C1(new_n732), .C2(new_n739), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n742), .A2(new_n743), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n749), .A2(new_n763), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT88), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(KEYINPUT88), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n702), .A2(G35), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G162), .B2(new_n702), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT29), .B(G2090), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n702), .A2(G26), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n473), .A2(G140), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n785));
  INV_X1    g360(.A(G116), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G2105), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n478), .B2(G128), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n676), .A2(G20), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT23), .Z(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT89), .B(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n781), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n676), .A2(G4), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n602), .B2(new_n676), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1348), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n676), .A2(G19), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n543), .B2(new_n676), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1341), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n797), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  AND4_X1   g379(.A1(new_n716), .A2(new_n776), .A3(new_n777), .A4(new_n804), .ZN(G311));
  NAND4_X1  g380(.A1(new_n716), .A2(new_n776), .A3(new_n777), .A4(new_n804), .ZN(G150));
  AOI22_X1  g381(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(new_n504), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n513), .A2(G93), .B1(new_n508), .B2(G55), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G860), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT91), .B(KEYINPUT37), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n595), .A2(new_n603), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n543), .B(new_n810), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n817), .B(new_n818), .Z(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n811), .B1(new_n820), .B2(KEYINPUT39), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n814), .B1(new_n821), .B2(new_n822), .ZN(G145));
  XNOR2_X1  g398(.A(new_n709), .B(KEYINPUT94), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n618), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n726), .B(new_n738), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n495), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n494), .B1(new_n459), .B2(new_n491), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n484), .B(new_n488), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n789), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n478), .A2(G130), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n460), .A2(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n473), .B2(G142), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n831), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n827), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n480), .B(new_n615), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G160), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(G37), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n838), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n693), .B(G166), .ZN(new_n847));
  XNOR2_X1  g422(.A(G305), .B(G290), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n846), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(KEYINPUT42), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n852), .B(KEYINPUT42), .C1(new_n846), .C2(new_n850), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n818), .B(new_n606), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n595), .B(G299), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(KEYINPUT41), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n853), .B2(new_n854), .ZN(new_n861));
  OAI21_X1  g436(.A(G868), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(G868), .B2(new_n810), .ZN(G295));
  OAI21_X1  g438(.A(new_n862), .B1(G868), .B2(new_n810), .ZN(G331));
  OR2_X1    g439(.A1(G168), .A2(G171), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(G286), .B2(G301), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n818), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n868), .B1(new_n856), .B2(new_n867), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(KEYINPUT97), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n873), .B2(new_n850), .ZN(new_n874));
  INV_X1    g449(.A(new_n868), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n867), .A2(new_n856), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n870), .B1(new_n877), .B2(new_n869), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n849), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT43), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n850), .B(new_n870), .C1(new_n877), .C2(new_n869), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n877), .B2(new_n850), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n872), .A2(KEYINPUT98), .A3(new_n849), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n881), .A2(new_n883), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT44), .B1(new_n880), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n874), .B2(new_n879), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n889), .B1(new_n892), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(G164), .B2(G1384), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT99), .B(G40), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n465), .A2(new_n468), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(G1996), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT100), .Z(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n726), .ZN(new_n902));
  INV_X1    g477(.A(G2067), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n789), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT101), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n899), .B1(new_n905), .B2(new_n727), .ZN(new_n906));
  INV_X1    g481(.A(G1996), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n902), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n899), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n710), .A2(new_n712), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n710), .A2(new_n712), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(G290), .B(G1986), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n828), .A2(new_n829), .ZN(new_n918));
  OAI211_X1 g493(.A(KEYINPUT45), .B(new_n917), .C1(new_n918), .C2(new_n489), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n895), .A2(new_n898), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n895), .A2(new_n919), .A3(KEYINPUT102), .A4(new_n898), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n679), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n897), .ZN(new_n925));
  NAND2_X1  g500(.A1(G160), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n830), .A2(new_n917), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n927), .B2(KEYINPUT50), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(KEYINPUT50), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(KEYINPUT103), .B(G2090), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G303), .A2(G8), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT55), .Z(new_n937));
  NAND3_X1  g512(.A1(new_n924), .A2(KEYINPUT104), .A3(new_n932), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n935), .A2(G8), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n926), .A2(new_n927), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT105), .B(G8), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(G651), .B1(new_n580), .B2(new_n581), .ZN(new_n944));
  AOI21_X1  g519(.A(G1981), .B1(new_n508), .B2(G48), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n575), .A2(KEYINPUT77), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n577), .B1(new_n513), .B2(G86), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n576), .A2(new_n578), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(KEYINPUT108), .A3(new_n944), .A4(new_n945), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n575), .A2(new_n584), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT109), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n575), .A2(new_n584), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n944), .A3(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n950), .A2(new_n952), .B1(G1981), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n943), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n962));
  AOI221_X4 g537(.A(new_n962), .B1(new_n957), .B2(G1981), .C1(new_n950), .C2(new_n952), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n940), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(G1981), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT108), .B1(new_n583), .B2(new_n945), .ZN(new_n966));
  INV_X1    g541(.A(new_n952), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n959), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n958), .A2(KEYINPUT49), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(KEYINPUT111), .A3(new_n970), .A4(new_n943), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n687), .A2(G1976), .A3(new_n692), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n973), .A2(KEYINPUT106), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n687), .A2(new_n975), .A3(new_n692), .A4(G1976), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n943), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT52), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(KEYINPUT106), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT107), .B(G1976), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT52), .B1(G288), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n979), .A2(new_n981), .A3(new_n943), .A4(new_n976), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT112), .B1(new_n972), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n978), .A2(new_n982), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n964), .A2(new_n971), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n939), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(G288), .A2(G1976), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n966), .A2(new_n967), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n942), .B(new_n941), .C1(new_n991), .C2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT113), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n939), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n972), .A2(KEYINPUT112), .A3(new_n983), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n986), .B1(new_n985), .B2(new_n987), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n991), .A2(new_n993), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n943), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n995), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n937), .ZN(new_n1005));
  INV_X1    g580(.A(new_n942), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n933), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n939), .A2(new_n985), .A3(new_n987), .A4(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n928), .A2(new_n930), .A3(new_n770), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n920), .A2(new_n743), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n1006), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(G286), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n937), .B1(new_n1006), .B2(new_n933), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n924), .A2(KEYINPUT104), .A3(new_n932), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT104), .B1(new_n924), .B2(new_n932), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1017), .B1(new_n1021), .B2(new_n937), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n972), .A2(new_n983), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1014), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1016), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n939), .A2(KEYINPUT63), .A3(new_n1014), .ZN(new_n1028));
  OAI221_X1 g603(.A(new_n1028), .B1(new_n937), .B2(new_n1021), .C1(new_n997), .C2(new_n998), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G301), .ZN(new_n1031));
  OR3_X1    g606(.A1(new_n920), .A2(KEYINPUT123), .A3(G2078), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT123), .B1(new_n920), .B2(G2078), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(KEYINPUT53), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n928), .A2(new_n930), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n747), .ZN(new_n1037));
  AOI21_X1  g612(.A(G2078), .B1(new_n922), .B2(new_n923), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(KEYINPUT53), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1031), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G168), .A2(new_n942), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1013), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1020), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT51), .B1(new_n1045), .B2(new_n1042), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1012), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(new_n1043), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1012), .A2(KEYINPUT122), .A3(new_n1042), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1040), .B1(new_n1053), .B2(KEYINPUT62), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1009), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1054), .B(new_n1055), .C1(KEYINPUT62), .C2(new_n1053), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1004), .A2(new_n1030), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT126), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G164), .A2(G1384), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n898), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n929), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(G1961), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n922), .A2(new_n923), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n752), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G301), .B1(new_n1068), .B2(new_n1034), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT124), .B(G2078), .Z(new_n1070));
  AND3_X1   g645(.A1(new_n1070), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n895), .A2(new_n919), .A3(G160), .A4(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1037), .B(new_n1072), .C1(new_n1038), .C2(KEYINPUT53), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n1031), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1059), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(new_n1022), .A3(new_n1053), .A4(new_n1024), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1059), .B1(new_n1073), .B2(G171), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(G301), .A3(new_n1037), .A4(new_n1034), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1058), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT125), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1040), .B1(new_n1031), .B2(new_n1073), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1089), .A2(new_n1059), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1088), .A2(new_n1090), .A3(KEYINPUT126), .A4(new_n1055), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT58), .B(G1341), .ZN(new_n1092));
  OAI22_X1  g667(.A1(G1996), .A2(new_n920), .B1(new_n941), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n543), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(KEYINPUT59), .Z(new_n1095));
  INV_X1    g670(.A(G1956), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(new_n732), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n920), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1036), .A2(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AND2_X1   g676(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT117), .B1(new_n920), .B2(new_n1098), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(KEYINPUT61), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1104), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1095), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n595), .B(KEYINPUT121), .ZN(new_n1111));
  INV_X1    g686(.A(G1348), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1036), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n941), .A2(new_n903), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT118), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1063), .B2(G1348), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT60), .B(new_n1111), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(KEYINPUT118), .A3(new_n1114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n602), .A2(KEYINPUT121), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1119), .B(new_n1123), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT61), .B1(new_n1108), .B2(KEYINPUT120), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1106), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1127), .B1(new_n1108), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1110), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1115), .A2(new_n1118), .A3(new_n595), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1132), .B(new_n1106), .C1(new_n1133), .C2(new_n1108), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1106), .B1(new_n1133), .B2(new_n1108), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT119), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1131), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1084), .A2(new_n1091), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n916), .B1(new_n1057), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n906), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT46), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT47), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n909), .A2(new_n911), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n784), .A2(new_n903), .A3(new_n788), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n899), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n899), .A2(G1986), .A3(G290), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT48), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n914), .A2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1143), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1139), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1139), .A2(KEYINPUT127), .A3(new_n1150), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g730(.A(G319), .ZN(new_n1157));
  NOR4_X1   g731(.A1(G229), .A2(new_n1157), .A3(G401), .A4(G227), .ZN(new_n1158));
  OAI211_X1 g732(.A(new_n844), .B(new_n1158), .C1(new_n890), .C2(new_n891), .ZN(G225));
  INV_X1    g733(.A(G225), .ZN(G308));
endmodule


