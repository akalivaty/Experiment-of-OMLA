//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G127gat), .B(G134gat), .Z(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT1), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G113gat), .A2(G120gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT69), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n211), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n210), .B1(new_n218), .B2(new_n219), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G141gat), .B(G148gat), .Z(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT2), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G155gat), .B(G162gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n224), .A2(new_n229), .A3(new_n227), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n223), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n220), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n218), .A2(new_n219), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n210), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n222), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n232), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n209), .B1(new_n234), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n239), .B2(new_n240), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n233), .A3(KEYINPUT4), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n239), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT76), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n240), .B(new_n248), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT76), .A3(new_n239), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n247), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n241), .A2(new_n208), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n243), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT4), .B1(new_n223), .B2(new_n233), .ZN(new_n260));
  NOR4_X1   g059(.A1(new_n221), .A2(new_n240), .A3(new_n244), .A4(new_n222), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT76), .B1(new_n254), .B2(new_n239), .ZN(new_n263));
  AND4_X1   g062(.A1(KEYINPUT76), .A2(new_n249), .A3(new_n239), .A4(new_n250), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n208), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n207), .B1(new_n259), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n256), .A2(new_n266), .A3(new_n208), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n265), .A2(new_n257), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n270), .B(new_n206), .C1(new_n271), .C2(new_n243), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(KEYINPUT6), .B(new_n207), .C1(new_n259), .C2(new_n268), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT23), .Z(new_n278));
  AOI21_X1  g077(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT64), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(G183gat), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n282), .B1(new_n281), .B2(new_n286), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n278), .B(new_n279), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n280), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT66), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n278), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT25), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n277), .A2(KEYINPUT68), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT68), .B1(new_n277), .B2(new_n295), .ZN(new_n297));
  OAI221_X1 g096(.A(new_n291), .B1(new_n295), .B2(new_n277), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n285), .ZN(new_n300));
  XOR2_X1   g099(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n301));
  AOI22_X1  g100(.A1(new_n300), .A2(new_n301), .B1(G183gat), .B2(G190gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n285), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n294), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n309), .B(KEYINPUT74), .Z(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n294), .A2(new_n305), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n312), .B2(new_n289), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(G211gat), .ZN(new_n316));
  INV_X1    g115(.A(G218gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(KEYINPUT22), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G211gat), .B(G218gat), .Z(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n311), .A2(new_n314), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n320), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n319), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n310), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n306), .B2(new_n307), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n326), .B2(new_n313), .ZN(new_n327));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G64gat), .ZN(new_n329));
  INV_X1    g128(.A(G92gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n322), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n322), .A2(new_n327), .A3(KEYINPUT30), .A4(new_n331), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n322), .A2(new_n327), .ZN(new_n337));
  INV_X1    g136(.A(new_n331), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI211_X1 g138(.A(KEYINPUT75), .B(new_n331), .C1(new_n322), .C2(new_n327), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n334), .B(new_n335), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(G228gat), .A2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n307), .B1(new_n240), .B2(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n324), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n321), .A2(new_n307), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n233), .B1(new_n350), .B2(new_n248), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n346), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n353));
  INV_X1    g152(.A(G22gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT77), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n324), .A2(KEYINPUT29), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n240), .B1(new_n358), .B2(KEYINPUT3), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n359), .A2(new_n348), .B1(KEYINPUT78), .B2(new_n345), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n355), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n343), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT31), .B(G50gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n355), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n352), .A2(new_n356), .ZN(new_n365));
  INV_X1    g164(.A(new_n343), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT77), .A4(new_n366), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n362), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n363), .B1(new_n362), .B2(new_n367), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT83), .B(KEYINPUT35), .Z(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AND4_X1   g171(.A1(new_n276), .A2(new_n342), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT70), .B1(new_n306), .B2(new_n239), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n312), .A2(new_n375), .A3(new_n223), .A4(new_n289), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n306), .A2(new_n239), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT32), .ZN(new_n382));
  XNOR2_X1  g181(.A(G15gat), .B(G43gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n386), .B2(KEYINPUT33), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(KEYINPUT33), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT71), .B1(new_n390), .B2(new_n386), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n378), .A2(new_n380), .B1(new_n382), .B2(KEYINPUT33), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n392), .A2(new_n393), .A3(new_n385), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n388), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n374), .A2(new_n376), .A3(new_n377), .A4(new_n379), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT34), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(KEYINPUT73), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n390), .A2(KEYINPUT71), .A3(new_n386), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n393), .B1(new_n392), .B2(new_n385), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n402), .A2(new_n403), .B1(new_n381), .B2(new_n387), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n373), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n400), .A2(KEYINPUT72), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n410), .ZN(new_n411));
  OAI221_X1 g210(.A(new_n388), .B1(new_n400), .B2(KEYINPUT72), .C1(new_n391), .C2(new_n394), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n370), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n342), .A2(new_n276), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT35), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n370), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT80), .B(KEYINPUT39), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n256), .A2(KEYINPUT79), .A3(new_n208), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n265), .B2(new_n209), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT79), .B1(new_n256), .B2(new_n208), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n265), .A2(new_n421), .A3(new_n209), .ZN(new_n425));
  OR3_X1    g224(.A1(new_n234), .A2(new_n241), .A3(new_n209), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT39), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n427), .A3(new_n206), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT40), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n423), .A2(new_n427), .A3(KEYINPUT40), .A4(new_n206), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n430), .A2(new_n269), .A3(new_n341), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n370), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT38), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT37), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n322), .A2(new_n327), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n322), .B2(new_n327), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(new_n331), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n439), .B2(KEYINPUT82), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n438), .B2(new_n331), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n434), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n337), .A2(KEYINPUT37), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n444), .A2(new_n434), .A3(new_n338), .A4(new_n436), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n439), .A2(KEYINPUT81), .A3(new_n434), .A4(new_n436), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n274), .A2(new_n275), .A3(new_n332), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n443), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n418), .B1(new_n433), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT36), .B1(new_n401), .B2(new_n407), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n411), .B2(new_n412), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n416), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G229gat), .A2(G233gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n458), .B(KEYINPUT88), .Z(new_n459));
  XOR2_X1   g258(.A(new_n459), .B(KEYINPUT13), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n462));
  XOR2_X1   g261(.A(G43gat), .B(G50gat), .Z(new_n463));
  INV_X1    g262(.A(KEYINPUT15), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT15), .ZN(new_n467));
  NAND2_X1  g266(.A1(G29gat), .A2(G36gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT14), .ZN(new_n469));
  INV_X1    g268(.A(G29gat), .ZN(new_n470));
  INV_X1    g269(.A(G36gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NOR4_X1   g275(.A1(KEYINPUT85), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  NOR2_X1   g277(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(new_n471), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n473), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT86), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(KEYINPUT86), .B(new_n473), .C1(new_n477), .C2(new_n480), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n468), .ZN(new_n485));
  INV_X1    g284(.A(new_n467), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n476), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488));
  INV_X1    g287(.A(G1gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT16), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT87), .B1(new_n488), .B2(G1gat), .ZN(new_n493));
  OAI21_X1  g292(.A(G8gat), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n488), .A2(G1gat), .ZN(new_n495));
  INV_X1    g294(.A(G8gat), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n495), .A2(KEYINPUT87), .A3(new_n496), .A4(new_n491), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n462), .B1(new_n487), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n468), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n481), .B2(new_n482), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n467), .B1(new_n502), .B2(new_n484), .ZN(new_n503));
  OAI211_X1 g302(.A(KEYINPUT89), .B(new_n498), .C1(new_n503), .C2(new_n476), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506));
  INV_X1    g305(.A(new_n473), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n472), .A2(KEYINPUT85), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n479), .A2(new_n478), .A3(new_n471), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n468), .B1(new_n510), .B2(KEYINPUT86), .ZN(new_n511));
  INV_X1    g310(.A(new_n484), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n486), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n475), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n506), .B1(new_n514), .B2(new_n498), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n487), .A2(KEYINPUT90), .A3(new_n499), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n461), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n503), .B2(new_n476), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(KEYINPUT17), .A3(new_n475), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n499), .ZN(new_n522));
  INV_X1    g321(.A(new_n459), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n514), .A2(new_n498), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n522), .A2(KEYINPUT18), .A3(new_n523), .A4(new_n524), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n518), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G169gat), .B(G197gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT12), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n518), .A2(new_n527), .A3(new_n528), .A4(new_n535), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G57gat), .B(G64gat), .Z(new_n540));
  INV_X1    g339(.A(KEYINPUT9), .ZN(new_n541));
  INV_X1    g340(.A(G71gat), .ZN(new_n542));
  INV_X1    g341(.A(G78gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G71gat), .B(G78gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(new_n546), .A3(new_n544), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n498), .B1(KEYINPUT21), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT21), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G127gat), .B(G155gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n316), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n550), .B2(new_n553), .ZN(new_n560));
  AOI211_X1 g359(.A(KEYINPUT21), .B(new_n555), .C1(new_n548), .C2(new_n549), .ZN(new_n561));
  OAI21_X1  g360(.A(G211gat), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n565), .B1(new_n559), .B2(new_n562), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n552), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n559), .A2(new_n562), .ZN(new_n570));
  INV_X1    g369(.A(new_n565), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n552), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n566), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT91), .B(G183gat), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n575), .B1(new_n569), .B2(new_n574), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT41), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n579), .B(new_n582), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT7), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT92), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(KEYINPUT92), .A3(new_n589), .ZN(new_n592));
  NOR2_X1   g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT8), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT93), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n591), .B2(new_n597), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n587), .A2(KEYINPUT7), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n593), .B1(new_n604), .B2(new_n585), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n605), .A2(new_n606), .A3(new_n599), .A4(new_n596), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n520), .A2(new_n521), .A3(new_n600), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OAI22_X1  g410(.A1(new_n611), .A2(KEYINPUT94), .B1(new_n581), .B2(new_n580), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n600), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n514), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(KEYINPUT94), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n609), .B2(new_n614), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n584), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n583), .A3(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n550), .A3(new_n600), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n602), .A2(new_n548), .A3(new_n549), .A4(new_n607), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n551), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n627), .A2(KEYINPUT95), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT95), .B1(new_n627), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n623), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n624), .A2(new_n626), .ZN(new_n632));
  INV_X1    g431(.A(new_n623), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G176gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G204gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n627), .A2(new_n628), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n623), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n634), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n637), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n578), .A2(new_n622), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n457), .A2(new_n539), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n276), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n489), .ZN(G1324gat));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n342), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT96), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n496), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT97), .Z(new_n656));
  OAI221_X1 g455(.A(new_n656), .B1(new_n654), .B2(new_n653), .C1(new_n496), .C2(new_n650), .ZN(G1325gat));
  NOR2_X1   g456(.A1(new_n453), .A2(new_n455), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n647), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n408), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(G15gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n647), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT98), .ZN(G1326gat));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n370), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  OAI211_X1 g465(.A(new_n658), .B(new_n418), .C1(new_n451), .C2(new_n433), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n622), .B1(new_n667), .B2(new_n416), .ZN(new_n668));
  INV_X1    g467(.A(new_n539), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n669), .A2(new_n578), .A3(new_n644), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n276), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n470), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n583), .B1(new_n620), .B2(new_n616), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n617), .A2(new_n584), .A3(new_n618), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n619), .A2(new_n621), .A3(KEYINPUT99), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n457), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n668), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n672), .A3(new_n670), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n674), .B1(new_n686), .B2(new_n470), .ZN(G1328gat));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n471), .A3(new_n341), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT46), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n670), .ZN(new_n690));
  OAI21_X1  g489(.A(G36gat), .B1(new_n690), .B2(new_n342), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(G1329gat));
  OAI21_X1  g491(.A(G43gat), .B1(new_n690), .B2(new_n658), .ZN(new_n693));
  INV_X1    g492(.A(G43gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n671), .A2(new_n694), .A3(new_n408), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  INV_X1    g497(.A(new_n622), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n683), .B1(new_n457), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n681), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n667), .B2(new_n416), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n417), .B(new_n670), .C1(new_n700), .C2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n684), .A2(KEYINPUT101), .A3(new_n417), .A4(new_n670), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(G50gat), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n370), .A2(G50gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT100), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n671), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n698), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n703), .A2(G50gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n698), .A3(new_n710), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT102), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n716));
  INV_X1    g515(.A(G50gat), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n703), .B2(new_n704), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n718), .A2(new_n706), .B1(new_n671), .B2(new_n709), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n716), .B(new_n713), .C1(new_n719), .C2(new_n698), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n715), .A2(new_n720), .ZN(G1331gat));
  INV_X1    g520(.A(new_n578), .ZN(new_n722));
  NOR4_X1   g521(.A1(new_n722), .A2(new_n539), .A3(new_n699), .A4(new_n645), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n457), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n276), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(G57gat), .Z(G1332gat));
  XOR2_X1   g525(.A(new_n724), .B(KEYINPUT103), .Z(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n341), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT49), .B(G64gat), .Z(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(G1333gat));
  OAI21_X1  g530(.A(new_n542), .B1(new_n724), .B2(new_n660), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n658), .A2(new_n542), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n727), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n733), .B1(new_n727), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n727), .A2(new_n417), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT105), .B(G78gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  NAND2_X1  g540(.A1(new_n669), .A2(new_n722), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n645), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n684), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n672), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n205), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n746), .B2(new_n745), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n457), .A2(new_n699), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(KEYINPUT51), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n749), .A2(new_n742), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(KEYINPUT107), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n750), .B(KEYINPUT51), .C1(new_n749), .C2(new_n742), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(new_n644), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n205), .A3(new_n672), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n748), .A2(new_n757), .ZN(G1336gat));
  NOR2_X1   g557(.A1(new_n342), .A2(G92gat), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n754), .A2(new_n644), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n684), .A2(new_n341), .A3(new_n743), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(KEYINPUT52), .A3(G92gat), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT108), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n760), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n330), .B1(new_n761), .B2(KEYINPUT109), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(KEYINPUT109), .B2(new_n761), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(new_n760), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n765), .B1(new_n769), .B2(new_n763), .ZN(G1337gat));
  AOI21_X1  g569(.A(G99gat), .B1(new_n756), .B2(new_n408), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n456), .A2(G99gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n744), .B2(new_n772), .ZN(G1338gat));
  NOR2_X1   g572(.A1(new_n370), .A2(G106gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n744), .A2(new_n417), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n756), .A2(new_n774), .B1(new_n775), .B2(G106gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1339gat));
  AOI21_X1  g577(.A(KEYINPUT110), .B1(new_n646), .B2(new_n669), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n578), .A2(new_n622), .A3(new_n645), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(new_n539), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT90), .B1(new_n487), .B2(new_n499), .ZN(new_n784));
  NOR4_X1   g583(.A1(new_n503), .A2(new_n498), .A3(new_n506), .A4(new_n476), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n500), .A2(new_n504), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n460), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n522), .A2(new_n524), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n459), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n534), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n538), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n678), .A3(new_n679), .ZN(new_n794));
  AOI211_X1 g593(.A(KEYINPUT54), .B(new_n633), .C1(new_n627), .C2(new_n628), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT112), .B1(new_n795), .B2(new_n638), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n797), .B(new_n637), .C1(new_n641), .C2(KEYINPUT54), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT111), .B1(new_n640), .B2(new_n623), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n627), .A2(new_n628), .A3(new_n800), .A4(new_n633), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT95), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n640), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n627), .A2(KEYINPUT95), .A3(new_n628), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n633), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n796), .B(new_n798), .C1(new_n802), .C2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n801), .A2(KEYINPUT54), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n631), .A2(new_n799), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n796), .A4(new_n798), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n639), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n794), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n644), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n460), .B1(new_n786), .B2(new_n787), .ZN(new_n816));
  AND4_X1   g615(.A1(KEYINPUT18), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n535), .B1(new_n818), .B2(new_n527), .ZN(new_n819));
  INV_X1    g618(.A(new_n538), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n809), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n812), .A2(new_n639), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n815), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n814), .B1(new_n680), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n783), .B1(new_n824), .B2(new_n578), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n370), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n276), .A2(new_n341), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n408), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n212), .A3(new_n669), .ZN(new_n831));
  INV_X1    g630(.A(new_n413), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n825), .A2(new_n672), .A3(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(KEYINPUT113), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(KEYINPUT113), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(new_n341), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n539), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n831), .B1(new_n837), .B2(new_n212), .ZN(G1340gat));
  NOR3_X1   g637(.A1(new_n830), .A2(new_n213), .A3(new_n645), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n644), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n213), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n836), .A2(new_n842), .A3(new_n578), .ZN(new_n843));
  OAI21_X1  g642(.A(G127gat), .B1(new_n830), .B2(new_n722), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n836), .A2(new_n846), .A3(new_n699), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n829), .B2(new_n699), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT114), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(G1343gat));
  INV_X1    g651(.A(G141gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n658), .A2(new_n827), .ZN(new_n854));
  XNOR2_X1  g653(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n825), .B2(new_n417), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n370), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n823), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n815), .B(KEYINPUT116), .C1(new_n821), .C2(new_n822), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n622), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n814), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n578), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n782), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n781), .B1(new_n780), .B2(new_n539), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n859), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n857), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT117), .B(new_n859), .C1(new_n865), .C2(new_n868), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n854), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n853), .B1(new_n873), .B2(new_n539), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n453), .A2(new_n455), .A3(new_n370), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n823), .A2(new_n680), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n578), .B1(new_n876), .B2(new_n864), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n875), .B(new_n672), .C1(new_n877), .C2(new_n868), .ZN(new_n878));
  NOR4_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n341), .A4(new_n669), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT58), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n644), .A2(new_n538), .A3(new_n792), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n537), .A2(new_n538), .B1(new_n807), .B2(new_n808), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n812), .A2(new_n639), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n622), .B1(new_n885), .B2(KEYINPUT116), .ZN(new_n886));
  INV_X1    g685(.A(new_n862), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n864), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n868), .B1(new_n888), .B2(new_n722), .ZN(new_n889));
  INV_X1    g688(.A(new_n859), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n870), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n857), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n872), .ZN(new_n893));
  INV_X1    g692(.A(new_n854), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n539), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G141gat), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n669), .A2(G141gat), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n825), .A2(KEYINPUT118), .A3(new_n672), .A4(new_n875), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n898), .A2(new_n342), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n881), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT119), .B(new_n903), .C1(new_n895), .C2(G141gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n880), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n880), .B(KEYINPUT120), .C1(new_n905), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1344gat));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  INV_X1    g711(.A(new_n873), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n912), .B(G148gat), .C1(new_n913), .C2(new_n645), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n825), .A2(new_n417), .A3(new_n856), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n780), .A2(new_n539), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n699), .B1(new_n823), .B2(new_n860), .ZN(new_n919));
  INV_X1    g718(.A(new_n813), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n793), .A2(new_n699), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n919), .A2(new_n862), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n922), .B2(new_n578), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n417), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n916), .B1(new_n924), .B2(KEYINPUT121), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926));
  AOI211_X1 g725(.A(new_n926), .B(KEYINPUT57), .C1(new_n923), .C2(new_n417), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n644), .B(new_n894), .C1(new_n925), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G148gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n915), .B1(new_n929), .B2(KEYINPUT59), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT122), .B(new_n912), .C1(new_n928), .C2(G148gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n914), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n898), .A2(new_n342), .A3(new_n900), .ZN(new_n933));
  INV_X1    g732(.A(G148gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n644), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(G1345gat));
  OAI21_X1  g735(.A(G155gat), .B1(new_n913), .B2(new_n722), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n225), .A3(new_n578), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1346gat));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n226), .A3(new_n699), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT123), .ZN(new_n941));
  OAI21_X1  g740(.A(G162gat), .B1(new_n913), .B2(new_n680), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n672), .A2(new_n342), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n408), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n826), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G169gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(new_n669), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n825), .A2(new_n276), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n341), .A3(new_n832), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT124), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n539), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n952), .B2(new_n947), .ZN(G1348gat));
  INV_X1    g752(.A(G176gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n954), .A3(new_n644), .ZN(new_n955));
  OAI21_X1  g754(.A(G176gat), .B1(new_n946), .B2(new_n645), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1349gat));
  NAND2_X1  g756(.A1(new_n578), .A2(new_n299), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(G183gat), .B1(new_n946), .B2(new_n722), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT125), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g762(.A(new_n680), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n951), .A2(new_n285), .A3(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(new_n946), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n285), .B1(new_n966), .B2(new_n699), .ZN(new_n967));
  OR2_X1    g766(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g767(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n965), .B(new_n970), .C1(new_n967), .C2(new_n968), .ZN(G1351gat));
  AND2_X1   g770(.A1(new_n875), .A2(new_n341), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n949), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(G197gat), .B1(new_n974), .B2(new_n539), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n920), .A2(new_n921), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n863), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n917), .B1(new_n977), .B2(new_n722), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n858), .B1(new_n978), .B2(new_n370), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n926), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n924), .A2(KEYINPUT121), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n980), .A2(new_n981), .A3(new_n916), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n658), .A2(new_n944), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n539), .A2(G197gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n975), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  NAND3_X1  g786(.A1(new_n982), .A2(new_n644), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G204gat), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n973), .A2(G204gat), .A3(new_n645), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(G1353gat));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n316), .A3(new_n578), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n982), .A2(new_n578), .A3(new_n984), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(KEYINPUT127), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n982), .A2(new_n996), .A3(new_n578), .A4(new_n984), .ZN(new_n997));
  AND4_X1   g796(.A1(KEYINPUT63), .A2(new_n995), .A3(G211gat), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n316), .B1(new_n994), .B2(KEYINPUT127), .ZN(new_n999));
  AOI21_X1  g798(.A(KEYINPUT63), .B1(new_n999), .B2(new_n997), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n993), .B1(new_n998), .B2(new_n1000), .ZN(G1354gat));
  AOI21_X1  g800(.A(G218gat), .B1(new_n974), .B2(new_n964), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n622), .A2(new_n317), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1002), .B1(new_n985), .B2(new_n1003), .ZN(G1355gat));
endmodule


