

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745;

  NOR2_X1 U372 ( .A1(n533), .A2(n546), .ZN(n625) );
  XNOR2_X2 U373 ( .A(n550), .B(n549), .ZN(n553) );
  NOR2_X2 U374 ( .A1(n565), .A2(n656), .ZN(n536) );
  XNOR2_X2 U375 ( .A(n514), .B(KEYINPUT22), .ZN(n565) );
  XNOR2_X2 U376 ( .A(n419), .B(G125), .ZN(n454) );
  AND2_X2 U377 ( .A1(n557), .A2(n652), .ZN(n648) );
  NOR2_X1 U378 ( .A1(n637), .A2(n626), .ZN(n563) );
  XNOR2_X2 U379 ( .A(n444), .B(n427), .ZN(n701) );
  XNOR2_X2 U380 ( .A(n417), .B(G131), .ZN(n475) );
  XNOR2_X1 U381 ( .A(n735), .B(n419), .ZN(n444) );
  XNOR2_X2 U382 ( .A(n418), .B(n455), .ZN(n735) );
  NOR2_X2 U383 ( .A1(n745), .A2(n579), .ZN(n580) );
  INV_X1 U384 ( .A(n525), .ZN(n638) );
  AND2_X1 U385 ( .A1(n369), .A2(n368), .ZN(n367) );
  NOR2_X1 U386 ( .A1(n552), .A2(n551), .ZN(n554) );
  NOR2_X1 U387 ( .A1(n381), .A2(n511), .ZN(n512) );
  XNOR2_X1 U388 ( .A(n483), .B(n482), .ZN(n533) );
  BUF_X1 U389 ( .A(n498), .Z(n594) );
  NOR2_X1 U390 ( .A1(G902), .A2(n707), .ZN(n483) );
  XNOR2_X1 U391 ( .A(n438), .B(G104), .ZN(n470) );
  XNOR2_X1 U392 ( .A(n379), .B(G110), .ZN(n451) );
  INV_X2 U393 ( .A(G113), .ZN(n438) );
  XOR2_X1 U394 ( .A(G137), .B(G140), .Z(n420) );
  INV_X2 U395 ( .A(G953), .ZN(n738) );
  INV_X1 U396 ( .A(KEYINPUT70), .ZN(n417) );
  OR2_X1 U397 ( .A1(n390), .A2(n383), .ZN(n382) );
  NOR2_X2 U398 ( .A1(n538), .A2(n537), .ZN(n552) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n466) );
  XOR2_X1 U400 ( .A(KEYINPUT98), .B(KEYINPUT96), .Z(n468) );
  NOR2_X1 U401 ( .A1(n673), .A2(n564), .ZN(n569) );
  XNOR2_X1 U402 ( .A(n394), .B(n454), .ZN(n472) );
  XOR2_X1 U403 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n394) );
  NAND2_X1 U404 ( .A1(n350), .A2(n355), .ZN(n386) );
  XNOR2_X1 U405 ( .A(n454), .B(n453), .ZN(n393) );
  XNOR2_X1 U406 ( .A(n392), .B(KEYINPUT78), .ZN(n391) );
  NAND2_X1 U407 ( .A1(n738), .A2(G224), .ZN(n392) );
  INV_X1 U408 ( .A(n533), .ZN(n547) );
  NAND2_X1 U409 ( .A1(n620), .A2(n616), .ZN(n368) );
  AND2_X1 U410 ( .A1(n359), .A2(n352), .ZN(n737) );
  XNOR2_X1 U411 ( .A(G116), .B(G101), .ZN(n435) );
  INV_X1 U412 ( .A(KEYINPUT76), .ZN(n379) );
  XNOR2_X1 U413 ( .A(n472), .B(n420), .ZN(n736) );
  XNOR2_X1 U414 ( .A(n403), .B(n395), .ZN(n404) );
  XNOR2_X1 U415 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n401) );
  XOR2_X1 U416 ( .A(KEYINPUT92), .B(G110), .Z(n398) );
  XOR2_X1 U417 ( .A(n481), .B(n480), .Z(n707) );
  XOR2_X1 U418 ( .A(G107), .B(G104), .Z(n421) );
  INV_X1 U419 ( .A(G101), .ZN(n423) );
  BUF_X1 U420 ( .A(n535), .Z(n656) );
  BUF_X1 U421 ( .A(n539), .Z(n584) );
  INV_X1 U422 ( .A(n722), .ZN(n371) );
  INV_X1 U423 ( .A(G237), .ZN(n446) );
  XNOR2_X1 U424 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U425 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U426 ( .A(G122), .ZN(n476) );
  NAND2_X1 U427 ( .A1(G234), .A2(G237), .ZN(n432) );
  OR2_X1 U428 ( .A1(n559), .A2(n528), .ZN(n448) );
  XNOR2_X1 U429 ( .A(KEYINPUT5), .B(G137), .ZN(n440) );
  XNOR2_X1 U430 ( .A(n377), .B(G122), .ZN(n488) );
  INV_X1 U431 ( .A(G107), .ZN(n377) );
  INV_X1 U432 ( .A(KEYINPUT16), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n361), .B(n353), .ZN(n726) );
  XOR2_X1 U434 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n400) );
  NAND2_X1 U435 ( .A1(n350), .A2(KEYINPUT64), .ZN(n383) );
  NAND2_X1 U436 ( .A1(n356), .A2(n386), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n393), .B(n391), .ZN(n457) );
  NAND2_X1 U438 ( .A1(n726), .A2(n737), .ZN(n614) );
  NOR2_X1 U439 ( .A1(n595), .A2(n571), .ZN(n463) );
  NAND2_X1 U440 ( .A1(n366), .A2(n351), .ZN(n365) );
  XNOR2_X1 U441 ( .A(n452), .B(n374), .ZN(n723) );
  XNOR2_X1 U442 ( .A(n378), .B(n375), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n488), .B(n376), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n451), .B(n470), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n736), .B(n404), .ZN(n405) );
  XNOR2_X1 U446 ( .A(G119), .B(G128), .ZN(n397) );
  XNOR2_X1 U447 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U448 ( .A(n424), .B(n423), .ZN(n425) );
  AND2_X1 U449 ( .A1(n621), .A2(G953), .ZN(n722) );
  NOR2_X1 U450 ( .A1(n581), .A2(n594), .ZN(n582) );
  XOR2_X1 U451 ( .A(n613), .B(KEYINPUT65), .Z(n350) );
  AND2_X1 U452 ( .A1(n373), .A2(G472), .ZN(n351) );
  AND2_X1 U453 ( .A1(n610), .A2(n609), .ZN(n352) );
  BUF_X1 U454 ( .A(n614), .Z(n645) );
  XOR2_X1 U455 ( .A(KEYINPUT85), .B(KEYINPUT45), .Z(n353) );
  XNOR2_X1 U456 ( .A(KEYINPUT87), .B(KEYINPUT48), .ZN(n354) );
  OR2_X1 U457 ( .A1(n612), .A2(n389), .ZN(n355) );
  INV_X1 U458 ( .A(KEYINPUT64), .ZN(n389) );
  OR2_X1 U459 ( .A1(n350), .A2(n389), .ZN(n356) );
  AND2_X1 U460 ( .A1(n612), .A2(n389), .ZN(n357) );
  XOR2_X1 U461 ( .A(n622), .B(KEYINPUT88), .Z(n358) );
  NAND2_X1 U462 ( .A1(n548), .A2(n597), .ZN(n550) );
  NOR2_X2 U463 ( .A1(n710), .A2(n722), .ZN(n712) );
  NAND2_X1 U464 ( .A1(n718), .A2(G475), .ZN(n709) );
  NOR2_X4 U465 ( .A1(n388), .A2(n615), .ZN(n718) );
  XNOR2_X1 U466 ( .A(n360), .B(n354), .ZN(n359) );
  NAND2_X1 U467 ( .A1(n608), .A2(n607), .ZN(n360) );
  NAND2_X1 U468 ( .A1(n363), .A2(n362), .ZN(n361) );
  XNOR2_X1 U469 ( .A(n570), .B(KEYINPUT102), .ZN(n362) );
  XNOR2_X1 U470 ( .A(n555), .B(n364), .ZN(n363) );
  INV_X1 U471 ( .A(KEYINPUT44), .ZN(n364) );
  NAND2_X1 U472 ( .A1(n367), .A2(n365), .ZN(n372) );
  INV_X1 U473 ( .A(n617), .ZN(n366) );
  NAND2_X1 U474 ( .A1(n617), .A2(n620), .ZN(n369) );
  XNOR2_X1 U475 ( .A(n370), .B(n358), .ZN(G57) );
  NAND2_X1 U476 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U477 ( .A(n620), .ZN(n373) );
  XNOR2_X1 U478 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U479 ( .A1(n589), .A2(n381), .ZN(n380) );
  XNOR2_X1 U480 ( .A(n499), .B(KEYINPUT19), .ZN(n381) );
  NAND2_X2 U481 ( .A1(n384), .A2(n382), .ZN(n388) );
  AND2_X2 U482 ( .A1(n387), .A2(n385), .ZN(n384) );
  NAND2_X1 U483 ( .A1(n390), .A2(n357), .ZN(n387) );
  INV_X1 U484 ( .A(n614), .ZN(n390) );
  BUF_X1 U485 ( .A(n515), .Z(n576) );
  XOR2_X1 U486 ( .A(n402), .B(n401), .Z(n395) );
  AND2_X1 U487 ( .A1(n413), .A2(G217), .ZN(n396) );
  INV_X1 U488 ( .A(n470), .ZN(n471) );
  XNOR2_X1 U489 ( .A(G475), .B(KEYINPUT13), .ZN(n482) );
  XNOR2_X1 U490 ( .A(n462), .B(n461), .ZN(n498) );
  XNOR2_X1 U491 ( .A(n709), .B(n708), .ZN(n710) );
  XOR2_X1 U492 ( .A(n398), .B(n397), .Z(n406) );
  INV_X2 U493 ( .A(G146), .ZN(n419) );
  NAND2_X1 U494 ( .A1(G234), .A2(n738), .ZN(n399) );
  XNOR2_X1 U495 ( .A(n400), .B(n399), .ZN(n492) );
  NAND2_X1 U496 ( .A1(G221), .A2(n492), .ZN(n403) );
  XOR2_X1 U497 ( .A(KEYINPUT83), .B(KEYINPUT73), .Z(n402) );
  XNOR2_X1 U498 ( .A(n406), .B(n405), .ZN(n719) );
  NOR2_X1 U499 ( .A1(n719), .A2(G902), .ZN(n412) );
  XOR2_X1 U500 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n410) );
  XNOR2_X1 U501 ( .A(G902), .B(KEYINPUT89), .ZN(n408) );
  INV_X1 U502 ( .A(KEYINPUT15), .ZN(n407) );
  XNOR2_X1 U503 ( .A(n408), .B(n407), .ZN(n611) );
  NAND2_X1 U504 ( .A1(n611), .A2(G234), .ZN(n409) );
  XNOR2_X1 U505 ( .A(n409), .B(KEYINPUT20), .ZN(n413) );
  XNOR2_X1 U506 ( .A(n410), .B(n396), .ZN(n411) );
  XNOR2_X1 U507 ( .A(n412), .B(n411), .ZN(n522) );
  INV_X1 U508 ( .A(n522), .ZN(n416) );
  AND2_X1 U509 ( .A1(n413), .A2(G221), .ZN(n415) );
  XNOR2_X1 U510 ( .A(KEYINPUT93), .B(KEYINPUT21), .ZN(n414) );
  XNOR2_X1 U511 ( .A(n415), .B(n414), .ZN(n649) );
  INV_X1 U512 ( .A(n649), .ZN(n523) );
  NAND2_X1 U513 ( .A1(n416), .A2(n523), .ZN(n655) );
  XNOR2_X1 U514 ( .A(n475), .B(G134), .ZN(n418) );
  XNOR2_X2 U515 ( .A(G143), .B(G128), .ZN(n486) );
  XNOR2_X1 U516 ( .A(n486), .B(KEYINPUT4), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n420), .B(n451), .ZN(n422) );
  XNOR2_X1 U518 ( .A(n422), .B(n421), .ZN(n426) );
  NAND2_X1 U519 ( .A1(G227), .A2(n738), .ZN(n424) );
  XNOR2_X1 U520 ( .A(n426), .B(n425), .ZN(n427) );
  INV_X1 U521 ( .A(G902), .ZN(n501) );
  NAND2_X1 U522 ( .A1(n701), .A2(n501), .ZN(n429) );
  XOR2_X1 U523 ( .A(KEYINPUT71), .B(G469), .Z(n428) );
  XNOR2_X2 U524 ( .A(n429), .B(n428), .ZN(n515) );
  NAND2_X1 U525 ( .A1(G953), .A2(G902), .ZN(n503) );
  NOR2_X1 U526 ( .A1(G900), .A2(n503), .ZN(n431) );
  NAND2_X1 U527 ( .A1(n738), .A2(G952), .ZN(n505) );
  INV_X1 U528 ( .A(n505), .ZN(n430) );
  OR2_X1 U529 ( .A1(n431), .A2(n430), .ZN(n433) );
  XNOR2_X1 U530 ( .A(n432), .B(KEYINPUT14), .ZN(n646) );
  AND2_X1 U531 ( .A1(n433), .A2(n646), .ZN(n521) );
  NAND2_X1 U532 ( .A1(n576), .A2(n521), .ZN(n434) );
  NOR2_X1 U533 ( .A1(n655), .A2(n434), .ZN(n450) );
  XNOR2_X1 U534 ( .A(n435), .B(KEYINPUT3), .ZN(n437) );
  XOR2_X1 U535 ( .A(KEYINPUT72), .B(G119), .Z(n436) );
  XNOR2_X1 U536 ( .A(n437), .B(n436), .ZN(n452) );
  NAND2_X1 U537 ( .A1(n466), .A2(G210), .ZN(n439) );
  XNOR2_X1 U538 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U539 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U540 ( .A(n452), .B(n442), .ZN(n443) );
  XNOR2_X1 U541 ( .A(n444), .B(n443), .ZN(n619) );
  OR2_X1 U542 ( .A1(n619), .A2(G902), .ZN(n445) );
  INV_X1 U543 ( .A(G472), .ZN(n616) );
  XNOR2_X2 U544 ( .A(n445), .B(n616), .ZN(n559) );
  NAND2_X1 U545 ( .A1(n501), .A2(n446), .ZN(n459) );
  AND2_X1 U546 ( .A1(n459), .A2(G214), .ZN(n528) );
  INV_X1 U547 ( .A(KEYINPUT30), .ZN(n447) );
  XNOR2_X1 U548 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U549 ( .A1(n450), .A2(n449), .ZN(n595) );
  XNOR2_X1 U550 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n453) );
  INV_X1 U551 ( .A(n455), .ZN(n456) );
  XNOR2_X1 U552 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U553 ( .A(n723), .B(n458), .ZN(n693) );
  NAND2_X1 U554 ( .A1(n693), .A2(n611), .ZN(n462) );
  NAND2_X1 U555 ( .A1(n459), .A2(G210), .ZN(n460) );
  XNOR2_X1 U556 ( .A(n460), .B(KEYINPUT90), .ZN(n461) );
  XOR2_X1 U557 ( .A(KEYINPUT38), .B(n594), .Z(n571) );
  XOR2_X1 U558 ( .A(KEYINPUT39), .B(n463), .Z(n534) );
  XOR2_X1 U559 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n465) );
  XNOR2_X1 U560 ( .A(G140), .B(KEYINPUT11), .ZN(n464) );
  XNOR2_X1 U561 ( .A(n465), .B(n464), .ZN(n481) );
  NAND2_X1 U562 ( .A1(G214), .A2(n466), .ZN(n467) );
  XNOR2_X1 U563 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U564 ( .A(KEYINPUT12), .B(n469), .Z(n474) );
  XNOR2_X1 U565 ( .A(n474), .B(n473), .ZN(n479) );
  XNOR2_X1 U566 ( .A(G143), .B(n475), .ZN(n477) );
  XOR2_X1 U567 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n485) );
  XNOR2_X1 U568 ( .A(G116), .B(G134), .ZN(n484) );
  XNOR2_X1 U569 ( .A(n485), .B(n484), .ZN(n491) );
  XOR2_X1 U570 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n487) );
  XOR2_X1 U571 ( .A(n487), .B(n486), .Z(n489) );
  XNOR2_X1 U572 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U573 ( .A(n491), .B(n490), .Z(n494) );
  NAND2_X1 U574 ( .A1(G217), .A2(n492), .ZN(n493) );
  XNOR2_X1 U575 ( .A(n494), .B(n493), .ZN(n713) );
  NOR2_X1 U576 ( .A1(G902), .A2(n713), .ZN(n495) );
  XNOR2_X1 U577 ( .A(n495), .B(G478), .ZN(n546) );
  NAND2_X1 U578 ( .A1(n533), .A2(n546), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n534), .A2(n638), .ZN(n497) );
  XNOR2_X1 U580 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n496) );
  XNOR2_X1 U581 ( .A(n497), .B(n496), .ZN(n579) );
  XOR2_X1 U582 ( .A(G131), .B(n579), .Z(G33) );
  NAND2_X1 U583 ( .A1(n547), .A2(n546), .ZN(n671) );
  NOR2_X1 U584 ( .A1(n671), .A2(n649), .ZN(n513) );
  NOR2_X1 U585 ( .A1(n498), .A2(n528), .ZN(n499) );
  NOR2_X1 U586 ( .A1(G898), .A2(n738), .ZN(n725) );
  NAND2_X1 U587 ( .A1(n725), .A2(KEYINPUT91), .ZN(n500) );
  NOR2_X1 U588 ( .A1(n501), .A2(n500), .ZN(n508) );
  NAND2_X1 U589 ( .A1(n508), .A2(n646), .ZN(n502) );
  AND2_X1 U590 ( .A1(n502), .A2(KEYINPUT91), .ZN(n510) );
  OR2_X1 U591 ( .A1(n503), .A2(G898), .ZN(n504) );
  NAND2_X1 U592 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U593 ( .A1(n506), .A2(n646), .ZN(n507) );
  NOR2_X1 U594 ( .A1(n508), .A2(n507), .ZN(n509) );
  NOR2_X1 U595 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X2 U596 ( .A(n512), .B(KEYINPUT0), .ZN(n562) );
  NAND2_X1 U597 ( .A1(n513), .A2(n562), .ZN(n514) );
  XNOR2_X1 U598 ( .A(n515), .B(KEYINPUT1), .ZN(n535) );
  INV_X1 U599 ( .A(n535), .ZN(n539) );
  NOR2_X1 U600 ( .A1(n416), .A2(n584), .ZN(n517) );
  XNOR2_X1 U601 ( .A(n559), .B(KEYINPUT6), .ZN(n566) );
  XNOR2_X1 U602 ( .A(n566), .B(KEYINPUT81), .ZN(n516) );
  NAND2_X1 U603 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U604 ( .A1(n565), .A2(n518), .ZN(n519) );
  XNOR2_X1 U605 ( .A(n519), .B(KEYINPUT32), .ZN(n551) );
  XNOR2_X1 U606 ( .A(G119), .B(KEYINPUT127), .ZN(n520) );
  XNOR2_X1 U607 ( .A(n551), .B(n520), .ZN(G21) );
  AND2_X1 U608 ( .A1(n522), .A2(n521), .ZN(n573) );
  NAND2_X1 U609 ( .A1(n523), .A2(n573), .ZN(n524) );
  NOR2_X1 U610 ( .A1(n525), .A2(n524), .ZN(n526) );
  AND2_X1 U611 ( .A1(n526), .A2(n566), .ZN(n527) );
  XNOR2_X1 U612 ( .A(n527), .B(KEYINPUT104), .ZN(n529) );
  INV_X1 U613 ( .A(n528), .ZN(n667) );
  NAND2_X1 U614 ( .A1(n529), .A2(n667), .ZN(n581) );
  XNOR2_X1 U615 ( .A(KEYINPUT105), .B(n581), .ZN(n530) );
  NAND2_X1 U616 ( .A1(n530), .A2(n584), .ZN(n531) );
  XNOR2_X1 U617 ( .A(n531), .B(KEYINPUT43), .ZN(n532) );
  NAND2_X1 U618 ( .A1(n532), .A2(n594), .ZN(n610) );
  XNOR2_X1 U619 ( .A(n610), .B(G140), .ZN(G42) );
  NAND2_X1 U620 ( .A1(n534), .A2(n625), .ZN(n609) );
  XNOR2_X1 U621 ( .A(n609), .B(G134), .ZN(G36) );
  XNOR2_X1 U622 ( .A(n536), .B(KEYINPUT103), .ZN(n538) );
  INV_X1 U623 ( .A(n416), .ZN(n650) );
  NAND2_X1 U624 ( .A1(n650), .A2(n559), .ZN(n537) );
  XOR2_X1 U625 ( .A(n552), .B(G110), .Z(G12) );
  NOR2_X2 U626 ( .A1(n539), .A2(n655), .ZN(n541) );
  INV_X1 U627 ( .A(KEYINPUT75), .ZN(n540) );
  XNOR2_X1 U628 ( .A(n541), .B(n540), .ZN(n557) );
  NAND2_X1 U629 ( .A1(n557), .A2(n566), .ZN(n543) );
  XNOR2_X1 U630 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n542) );
  XNOR2_X2 U631 ( .A(n543), .B(n542), .ZN(n676) );
  NAND2_X1 U632 ( .A1(n676), .A2(n562), .ZN(n545) );
  XOR2_X1 U633 ( .A(KEYINPUT80), .B(KEYINPUT34), .Z(n544) );
  XNOR2_X1 U634 ( .A(n545), .B(n544), .ZN(n548) );
  NOR2_X1 U635 ( .A1(n547), .A2(n546), .ZN(n597) );
  XNOR2_X1 U636 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n549) );
  XNOR2_X1 U637 ( .A(n553), .B(G122), .ZN(G24) );
  NAND2_X1 U638 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U639 ( .A1(n638), .A2(n625), .ZN(n556) );
  XNOR2_X1 U640 ( .A(KEYINPUT101), .B(n556), .ZN(n587) );
  INV_X1 U641 ( .A(n587), .ZN(n673) );
  INV_X1 U642 ( .A(n559), .ZN(n652) );
  NAND2_X1 U643 ( .A1(n648), .A2(n562), .ZN(n558) );
  XNOR2_X2 U644 ( .A(n558), .B(KEYINPUT31), .ZN(n637) );
  NAND2_X1 U645 ( .A1(n576), .A2(n559), .ZN(n560) );
  NOR2_X1 U646 ( .A1(n655), .A2(n560), .ZN(n561) );
  AND2_X1 U647 ( .A1(n562), .A2(n561), .ZN(n626) );
  XNOR2_X1 U648 ( .A(n563), .B(KEYINPUT94), .ZN(n564) );
  NOR2_X1 U649 ( .A1(n650), .A2(n566), .ZN(n567) );
  NAND2_X1 U650 ( .A1(n567), .A2(n584), .ZN(n568) );
  NOR2_X1 U651 ( .A1(n565), .A2(n568), .ZN(n623) );
  NOR2_X2 U652 ( .A1(n569), .A2(n623), .ZN(n570) );
  INV_X1 U653 ( .A(n571), .ZN(n668) );
  NAND2_X1 U654 ( .A1(n668), .A2(n667), .ZN(n672) );
  NOR2_X1 U655 ( .A1(n671), .A2(n672), .ZN(n572) );
  XNOR2_X1 U656 ( .A(n572), .B(KEYINPUT41), .ZN(n647) );
  NAND2_X1 U657 ( .A1(n573), .A2(n652), .ZN(n574) );
  NOR2_X1 U658 ( .A1(n649), .A2(n574), .ZN(n575) );
  XNOR2_X1 U659 ( .A(n575), .B(KEYINPUT28), .ZN(n577) );
  NAND2_X1 U660 ( .A1(n577), .A2(n576), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n647), .A2(n589), .ZN(n578) );
  XNOR2_X1 U662 ( .A(n578), .B(KEYINPUT42), .ZN(n745) );
  XNOR2_X1 U663 ( .A(n580), .B(KEYINPUT46), .ZN(n608) );
  INV_X1 U664 ( .A(KEYINPUT36), .ZN(n583) );
  XNOR2_X1 U665 ( .A(n583), .B(n582), .ZN(n585) );
  NOR2_X1 U666 ( .A1(n585), .A2(n584), .ZN(n642) );
  INV_X1 U667 ( .A(KEYINPUT82), .ZN(n586) );
  OR2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n588) );
  AND2_X1 U669 ( .A1(n588), .A2(KEYINPUT47), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n590), .A2(n380), .ZN(n593) );
  INV_X1 U671 ( .A(KEYINPUT47), .ZN(n591) );
  NAND2_X1 U672 ( .A1(n591), .A2(KEYINPUT82), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n593), .A2(n592), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT106), .ZN(n598) );
  AND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n633) );
  INV_X1 U677 ( .A(n633), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT47), .B(KEYINPUT67), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n380), .A2(n599), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n600), .A2(KEYINPUT82), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n587), .A2(n601), .ZN(n602) );
  AND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n642), .A2(n606), .ZN(n607) );
  INV_X1 U685 ( .A(n611), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n612), .A2(KEYINPUT2), .ZN(n613) );
  AND2_X1 U687 ( .A1(n390), .A2(KEYINPUT2), .ZN(n615) );
  INV_X1 U688 ( .A(n718), .ZN(n617) );
  XOR2_X1 U689 ( .A(KEYINPUT108), .B(KEYINPUT62), .Z(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n620) );
  INV_X1 U691 ( .A(G952), .ZN(n621) );
  XNOR2_X1 U692 ( .A(KEYINPUT109), .B(KEYINPUT63), .ZN(n622) );
  XOR2_X1 U693 ( .A(G101), .B(n623), .Z(G3) );
  NAND2_X1 U694 ( .A1(n626), .A2(n638), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(G104), .ZN(G6) );
  XNOR2_X1 U696 ( .A(G107), .B(KEYINPUT26), .ZN(n630) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT110), .Z(n628) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(G9) );
  XOR2_X1 U701 ( .A(G128), .B(KEYINPUT29), .Z(n632) );
  NAND2_X1 U702 ( .A1(n625), .A2(n380), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(G30) );
  XOR2_X1 U704 ( .A(G143), .B(n633), .Z(G45) );
  XOR2_X1 U705 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n635) );
  NAND2_X1 U706 ( .A1(n638), .A2(n380), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U708 ( .A(G146), .B(n636), .ZN(G48) );
  NAND2_X1 U709 ( .A1(n637), .A2(n638), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n639), .B(G113), .ZN(G15) );
  XOR2_X1 U711 ( .A(G116), .B(KEYINPUT113), .Z(n641) );
  NAND2_X1 U712 ( .A1(n637), .A2(n625), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(G18) );
  XNOR2_X1 U714 ( .A(G125), .B(n642), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U716 ( .A(KEYINPUT2), .B(KEYINPUT84), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n689) );
  NAND2_X1 U718 ( .A1(G952), .A2(n646), .ZN(n683) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U720 ( .A(KEYINPUT49), .B(n651), .ZN(n653) );
  NOR2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT114), .ZN(n661) );
  INV_X1 U723 ( .A(n655), .ZN(n657) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n659) );
  XNOR2_X1 U725 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U728 ( .A(KEYINPUT116), .B(n662), .Z(n663) );
  NOR2_X1 U729 ( .A1(n648), .A2(n663), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n664), .B(KEYINPUT51), .ZN(n665) );
  XNOR2_X1 U731 ( .A(KEYINPUT117), .B(n665), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n647), .A2(n666), .ZN(n680) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U734 ( .A(n669), .B(KEYINPUT118), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n678) );
  INV_X1 U738 ( .A(n676), .ZN(n677) );
  NOR2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U741 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U743 ( .A(KEYINPUT119), .B(n684), .ZN(n687) );
  INV_X1 U744 ( .A(n647), .ZN(n685) );
  NAND2_X1 U745 ( .A1(n685), .A2(n676), .ZN(n686) );
  NAND2_X1 U746 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U747 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U748 ( .A(KEYINPUT120), .B(n690), .Z(n691) );
  NOR2_X1 U749 ( .A1(G953), .A2(n691), .ZN(n692) );
  XNOR2_X1 U750 ( .A(KEYINPUT53), .B(n692), .ZN(G75) );
  NAND2_X1 U751 ( .A1(n718), .A2(G210), .ZN(n696) );
  XOR2_X1 U752 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n694) );
  XOR2_X1 U753 ( .A(n694), .B(n693), .Z(n695) );
  XNOR2_X1 U754 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X2 U755 ( .A1(n697), .A2(n722), .ZN(n700) );
  XOR2_X1 U756 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n698) );
  XNOR2_X1 U757 ( .A(KEYINPUT86), .B(n698), .ZN(n699) );
  XNOR2_X1 U758 ( .A(n700), .B(n699), .ZN(G51) );
  NAND2_X1 U759 ( .A1(n718), .A2(G469), .ZN(n704) );
  XOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  XOR2_X1 U761 ( .A(n702), .B(n701), .Z(n703) );
  XNOR2_X1 U762 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U763 ( .A1(n722), .A2(n705), .ZN(G54) );
  XOR2_X1 U764 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n706) );
  XNOR2_X1 U765 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n711) );
  XNOR2_X1 U766 ( .A(n712), .B(n711), .ZN(G60) );
  NAND2_X1 U767 ( .A1(n718), .A2(G478), .ZN(n715) );
  XOR2_X1 U768 ( .A(n713), .B(KEYINPUT123), .Z(n714) );
  XNOR2_X1 U769 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X2 U770 ( .A1(n716), .A2(n722), .ZN(n717) );
  XNOR2_X1 U771 ( .A(n717), .B(KEYINPUT124), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n718), .A2(G217), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n722), .A2(n721), .ZN(G66) );
  XOR2_X1 U775 ( .A(n723), .B(KEYINPUT126), .Z(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n734) );
  BUF_X1 U777 ( .A(n726), .Z(n727) );
  NAND2_X1 U778 ( .A1(n727), .A2(n738), .ZN(n732) );
  XOR2_X1 U779 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n729) );
  NAND2_X1 U780 ( .A1(G224), .A2(G953), .ZN(n728) );
  XNOR2_X1 U781 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U782 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(n733), .ZN(G69) );
  XOR2_X1 U785 ( .A(n736), .B(n735), .Z(n740) );
  XNOR2_X1 U786 ( .A(n737), .B(n740), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n739), .A2(n738), .ZN(n744) );
  XOR2_X1 U788 ( .A(n740), .B(G227), .Z(n741) );
  NAND2_X1 U789 ( .A1(n741), .A2(G900), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(G953), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n744), .A2(n743), .ZN(G72) );
  XOR2_X1 U792 ( .A(G137), .B(n745), .Z(G39) );
endmodule

