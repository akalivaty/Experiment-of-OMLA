

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(n728), .ZN(n722) );
  NOR2_X2 U556 ( .A1(n532), .A2(n531), .ZN(G160) );
  NOR2_X1 U557 ( .A1(G651), .A2(n631), .ZN(n650) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n696) );
  NOR2_X1 U559 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U560 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U561 ( .A(KEYINPUT23), .ZN(n523) );
  NOR2_X1 U562 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U563 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U564 ( .A(n757), .B(KEYINPUT65), .ZN(n758) );
  XNOR2_X1 U565 ( .A(KEYINPUT67), .B(G651), .ZN(n548) );
  NAND2_X1 U566 ( .A1(G160), .A2(G40), .ZN(n695) );
  XNOR2_X1 U567 ( .A(KEYINPUT78), .B(KEYINPUT13), .ZN(n577) );
  NOR2_X2 U568 ( .A1(n631), .A2(n548), .ZN(n657) );
  INV_X1 U569 ( .A(G2105), .ZN(n522) );
  XNOR2_X1 U570 ( .A(n578), .B(n577), .ZN(n579) );
  AND2_X2 U571 ( .A1(n522), .A2(G2104), .ZN(n881) );
  INV_X1 U572 ( .A(KEYINPUT99), .ZN(n539) );
  XNOR2_X1 U573 ( .A(KEYINPUT79), .B(n581), .ZN(n967) );
  NOR2_X2 U574 ( .A1(G2104), .A2(n522), .ZN(n877) );
  NAND2_X1 U575 ( .A1(n877), .A2(G125), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n881), .A2(G101), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U578 ( .A(KEYINPUT66), .B(n527), .ZN(n532) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n535) );
  NAND2_X1 U580 ( .A1(G113), .A2(n535), .ZN(n530) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XOR2_X2 U582 ( .A(KEYINPUT17), .B(n528), .Z(n880) );
  NAND2_X1 U583 ( .A1(G137), .A2(n880), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G138), .A2(n880), .ZN(n534) );
  NAND2_X1 U586 ( .A1(G102), .A2(n881), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n542) );
  NAND2_X1 U588 ( .A1(G126), .A2(n877), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n535), .A2(G114), .ZN(n536) );
  XNOR2_X1 U590 ( .A(n536), .B(KEYINPUT98), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U592 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U593 ( .A1(n542), .A2(n541), .ZN(G164) );
  NOR2_X2 U594 ( .A1(G651), .A2(G543), .ZN(n656) );
  NAND2_X1 U595 ( .A1(n656), .A2(G89), .ZN(n543) );
  XNOR2_X1 U596 ( .A(n543), .B(KEYINPUT4), .ZN(n545) );
  XOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .Z(n631) );
  NAND2_X1 U598 ( .A1(G76), .A2(n657), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U600 ( .A(n546), .B(KEYINPUT5), .ZN(n556) );
  NAND2_X1 U601 ( .A1(n650), .A2(G51), .ZN(n547) );
  XNOR2_X1 U602 ( .A(n547), .B(KEYINPUT82), .ZN(n553) );
  XNOR2_X1 U603 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n551) );
  NOR2_X1 U604 ( .A1(n548), .A2(G543), .ZN(n549) );
  XNOR2_X1 U605 ( .A(n549), .B(KEYINPUT1), .ZN(n550) );
  XNOR2_X2 U606 ( .A(n551), .B(n550), .ZN(n652) );
  NAND2_X1 U607 ( .A1(G63), .A2(n652), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U609 ( .A(KEYINPUT6), .B(n554), .Z(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U611 ( .A(n557), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(G111), .A2(n535), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G99), .A2(n881), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n564) );
  XOR2_X1 U617 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n561) );
  NAND2_X1 U618 ( .A1(G123), .A2(n877), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U620 ( .A(KEYINPUT86), .B(n562), .Z(n563) );
  NOR2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n880), .A2(G135), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n921) );
  XNOR2_X1 U624 ( .A(G2096), .B(n921), .ZN(n567) );
  OR2_X1 U625 ( .A1(G2100), .A2(n567), .ZN(G156) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G69), .ZN(G235) );
  INV_X1 U628 ( .A(G108), .ZN(G238) );
  INV_X1 U629 ( .A(G120), .ZN(G236) );
  INV_X1 U630 ( .A(G132), .ZN(G219) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n823) );
  NAND2_X1 U634 ( .A1(n823), .A2(G567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U636 ( .A1(n652), .A2(G56), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT14), .ZN(n572) );
  NAND2_X1 U638 ( .A1(G43), .A2(n650), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G68), .A2(n657), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT77), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n656), .A2(G81), .ZN(n574) );
  XOR2_X1 U643 ( .A(n574), .B(KEYINPUT12), .Z(n575) );
  NOR2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n578) );
  INV_X1 U645 ( .A(G860), .ZN(n612) );
  OR2_X1 U646 ( .A1(n967), .A2(n612), .ZN(G153) );
  NAND2_X1 U647 ( .A1(G64), .A2(n652), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G52), .A2(n650), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G90), .A2(n656), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G77), .A2(n657), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U653 ( .A(KEYINPUT9), .B(n586), .ZN(n587) );
  XNOR2_X1 U654 ( .A(KEYINPUT73), .B(n587), .ZN(n588) );
  NOR2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U656 ( .A(KEYINPUT74), .B(n590), .ZN(G171) );
  XOR2_X1 U657 ( .A(KEYINPUT80), .B(G171), .Z(G301) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U659 ( .A1(G54), .A2(n650), .ZN(n597) );
  NAND2_X1 U660 ( .A1(G66), .A2(n652), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G92), .A2(n656), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G79), .A2(n657), .ZN(n593) );
  XNOR2_X1 U664 ( .A(KEYINPUT81), .B(n593), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT15), .ZN(n975) );
  INV_X1 U668 ( .A(n975), .ZN(n893) );
  INV_X1 U669 ( .A(G868), .ZN(n674) );
  NAND2_X1 U670 ( .A1(n893), .A2(n674), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G65), .A2(n652), .ZN(n602) );
  NAND2_X1 U673 ( .A1(G78), .A2(n657), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G53), .A2(n650), .ZN(n603) );
  XNOR2_X1 U676 ( .A(KEYINPUT75), .B(n603), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n656), .A2(G91), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(G299) );
  XNOR2_X1 U680 ( .A(KEYINPUT83), .B(G868), .ZN(n608) );
  NOR2_X1 U681 ( .A1(G286), .A2(n608), .ZN(n610) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U684 ( .A(KEYINPUT84), .B(n611), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n612), .A2(G559), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n613), .A2(n975), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G559), .A2(n674), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n975), .A2(n615), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT85), .ZN(n618) );
  NOR2_X1 U691 ( .A1(n967), .A2(G868), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G559), .A2(n975), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(n967), .ZN(n671) );
  NOR2_X1 U695 ( .A1(n671), .A2(G860), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G67), .A2(n652), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G55), .A2(n650), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G93), .A2(n656), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G80), .A2(n657), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n673) );
  XOR2_X1 U703 ( .A(n626), .B(n673), .Z(G145) );
  NAND2_X1 U704 ( .A1(G49), .A2(n650), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U707 ( .A(KEYINPUT88), .B(n629), .ZN(n630) );
  NOR2_X1 U708 ( .A1(n652), .A2(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G86), .A2(n656), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G48), .A2(n650), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n657), .A2(G73), .ZN(n636) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n652), .A2(G61), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U719 ( .A1(n657), .A2(G72), .ZN(n641) );
  XNOR2_X1 U720 ( .A(n641), .B(KEYINPUT68), .ZN(n648) );
  NAND2_X1 U721 ( .A1(G85), .A2(n656), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G47), .A2(n650), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G60), .A2(n652), .ZN(n644) );
  XNOR2_X1 U725 ( .A(KEYINPUT71), .B(n644), .ZN(n645) );
  NOR2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(KEYINPUT72), .B(n649), .ZN(G290) );
  NAND2_X1 U729 ( .A1(G50), .A2(n650), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(KEYINPUT90), .ZN(n655) );
  NAND2_X1 U731 ( .A1(G62), .A2(n652), .ZN(n653) );
  XOR2_X1 U732 ( .A(KEYINPUT89), .B(n653), .Z(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n662) );
  NAND2_X1 U734 ( .A1(G88), .A2(n656), .ZN(n659) );
  NAND2_X1 U735 ( .A1(G75), .A2(n657), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT91), .B(n660), .Z(n661) );
  NOR2_X1 U738 ( .A1(n662), .A2(n661), .ZN(G166) );
  INV_X1 U739 ( .A(G166), .ZN(G303) );
  XOR2_X1 U740 ( .A(KEYINPUT19), .B(KEYINPUT92), .Z(n663) );
  XNOR2_X1 U741 ( .A(G288), .B(n663), .ZN(n664) );
  XNOR2_X1 U742 ( .A(KEYINPUT93), .B(n664), .ZN(n666) );
  XNOR2_X1 U743 ( .A(G305), .B(KEYINPUT94), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n667), .B(n673), .ZN(n669) );
  INV_X1 U746 ( .A(G299), .ZN(n968) );
  XNOR2_X1 U747 ( .A(n968), .B(G290), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U749 ( .A(n670), .B(G303), .ZN(n895) );
  XNOR2_X1 U750 ( .A(n671), .B(n895), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n672), .A2(G868), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n676), .A2(n675), .ZN(G295) );
  XOR2_X1 U754 ( .A(KEYINPUT21), .B(KEYINPUT95), .Z(n680) );
  NAND2_X1 U755 ( .A1(G2084), .A2(G2078), .ZN(n677) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U757 ( .A1(n678), .A2(G2090), .ZN(n679) );
  XNOR2_X1 U758 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U759 ( .A1(G2072), .A2(n681), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U761 ( .A(KEYINPUT76), .B(G82), .Z(G220) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U764 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(G96), .A2(n684), .ZN(n827) );
  NAND2_X1 U766 ( .A1(n827), .A2(G2106), .ZN(n689) );
  NOR2_X1 U767 ( .A1(G236), .A2(G238), .ZN(n686) );
  NOR2_X1 U768 ( .A1(G235), .A2(G237), .ZN(n685) );
  NAND2_X1 U769 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U770 ( .A(KEYINPUT96), .B(n687), .ZN(n828) );
  NAND2_X1 U771 ( .A1(n828), .A2(G567), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n829) );
  NAND2_X1 U773 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U774 ( .A1(n829), .A2(n690), .ZN(n826) );
  NAND2_X1 U775 ( .A1(n826), .A2(G36), .ZN(n691) );
  XOR2_X1 U776 ( .A(KEYINPUT97), .B(n691), .Z(G176) );
  NOR2_X1 U777 ( .A1(n696), .A2(n695), .ZN(n819) );
  NAND2_X1 U778 ( .A1(G1986), .A2(G290), .ZN(n971) );
  NOR2_X1 U779 ( .A1(G1986), .A2(G290), .ZN(n983) );
  INV_X1 U780 ( .A(n983), .ZN(n692) );
  NAND2_X1 U781 ( .A1(n971), .A2(n692), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n819), .A2(n693), .ZN(n694) );
  XOR2_X1 U783 ( .A(KEYINPUT100), .B(n694), .Z(n778) );
  INV_X1 U784 ( .A(n695), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X2 U786 ( .A(n698), .B(KEYINPUT64), .ZN(n728) );
  AND2_X1 U787 ( .A1(n728), .A2(G1341), .ZN(n699) );
  NOR2_X1 U788 ( .A1(n699), .A2(n967), .ZN(n702) );
  NAND2_X1 U789 ( .A1(n722), .A2(G1996), .ZN(n700) );
  XNOR2_X1 U790 ( .A(n700), .B(KEYINPUT26), .ZN(n701) );
  AND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n703) );
  OR2_X1 U792 ( .A1(n703), .A2(n975), .ZN(n709) );
  NAND2_X1 U793 ( .A1(n703), .A2(n975), .ZN(n707) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n722), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n728), .A2(G1348), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n715) );
  NAND2_X1 U799 ( .A1(n722), .A2(G2072), .ZN(n711) );
  XNOR2_X1 U800 ( .A(KEYINPUT102), .B(KEYINPUT27), .ZN(n710) );
  XNOR2_X1 U801 ( .A(n711), .B(n710), .ZN(n713) );
  INV_X1 U802 ( .A(G1956), .ZN(n997) );
  NOR2_X1 U803 ( .A1(n722), .A2(n997), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n716), .A2(n968), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U806 ( .A1(n716), .A2(n968), .ZN(n717) );
  XOR2_X1 U807 ( .A(n717), .B(KEYINPUT28), .Z(n718) );
  NAND2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U809 ( .A(KEYINPUT29), .B(KEYINPUT103), .ZN(n720) );
  XNOR2_X1 U810 ( .A(n721), .B(n720), .ZN(n726) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n941) );
  NAND2_X1 U812 ( .A1(n722), .A2(n941), .ZN(n724) );
  OR2_X1 U813 ( .A1(n722), .A2(G1961), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U815 ( .A1(n727), .A2(G171), .ZN(n725) );
  NAND2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n746) );
  NOR2_X1 U817 ( .A1(G171), .A2(n727), .ZN(n733) );
  NAND2_X1 U818 ( .A1(n728), .A2(G8), .ZN(n771) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n771), .ZN(n748) );
  NOR2_X1 U820 ( .A1(n728), .A2(G2084), .ZN(n744) );
  NOR2_X1 U821 ( .A1(n748), .A2(n744), .ZN(n729) );
  NAND2_X1 U822 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U824 ( .A1(G168), .A2(n731), .ZN(n732) );
  NOR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n735) );
  XOR2_X1 U826 ( .A(KEYINPUT31), .B(KEYINPUT104), .Z(n734) );
  XNOR2_X1 U827 ( .A(n735), .B(n734), .ZN(n745) );
  NAND2_X1 U828 ( .A1(n746), .A2(n745), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n736), .A2(G286), .ZN(n741) );
  NOR2_X1 U830 ( .A1(n728), .A2(G2090), .ZN(n738) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n771), .ZN(n737) );
  NOR2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U833 ( .A1(G303), .A2(n739), .ZN(n740) );
  NAND2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U835 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U836 ( .A(n743), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U837 ( .A1(G8), .A2(n744), .ZN(n750) );
  AND2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n769) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n759) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U844 ( .A1(n759), .A2(n753), .ZN(n976) );
  NAND2_X1 U845 ( .A1(n769), .A2(n976), .ZN(n756) );
  INV_X1 U846 ( .A(n771), .ZN(n754) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n972) );
  AND2_X1 U848 ( .A1(n754), .A2(n972), .ZN(n755) );
  NOR2_X1 U849 ( .A1(KEYINPUT33), .A2(n758), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n759), .A2(KEYINPUT33), .ZN(n760) );
  NOR2_X1 U851 ( .A1(n760), .A2(n771), .ZN(n761) );
  NOR2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U853 ( .A(KEYINPUT105), .B(G1981), .ZN(n763) );
  XNOR2_X1 U854 ( .A(n763), .B(G305), .ZN(n964) );
  NAND2_X1 U855 ( .A1(n764), .A2(n964), .ZN(n776) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XOR2_X1 U857 ( .A(n765), .B(KEYINPUT24), .Z(n766) );
  OR2_X1 U858 ( .A1(n771), .A2(n766), .ZN(n774) );
  NOR2_X1 U859 ( .A1(G2090), .A2(G303), .ZN(n767) );
  NAND2_X1 U860 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U863 ( .A(n772), .B(KEYINPUT106), .ZN(n773) );
  AND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  AND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n806) );
  NAND2_X1 U867 ( .A1(G129), .A2(n877), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G141), .A2(n880), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n881), .A2(G105), .ZN(n781) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n535), .A2(G117), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n867) );
  NAND2_X1 U875 ( .A1(G1996), .A2(n867), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G131), .A2(n880), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G95), .A2(n881), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G119), .A2(n877), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G107), .A2(n535), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n868) );
  NAND2_X1 U883 ( .A1(G1991), .A2(n868), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n932) );
  NAND2_X1 U885 ( .A1(n932), .A2(n819), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G140), .A2(n880), .ZN(n795) );
  NAND2_X1 U887 ( .A1(G104), .A2(n881), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n797) );
  XOR2_X1 U889 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n796) );
  XNOR2_X1 U890 ( .A(n797), .B(n796), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G128), .A2(n877), .ZN(n799) );
  NAND2_X1 U892 ( .A1(G116), .A2(n535), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U894 ( .A(KEYINPUT35), .B(n800), .Z(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U896 ( .A(KEYINPUT36), .B(n803), .Z(n889) );
  XOR2_X1 U897 ( .A(G2067), .B(KEYINPUT37), .Z(n818) );
  AND2_X1 U898 ( .A1(n889), .A2(n818), .ZN(n920) );
  NAND2_X1 U899 ( .A1(n920), .A2(n819), .ZN(n807) );
  AND2_X1 U900 ( .A1(n804), .A2(n807), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n817) );
  INV_X1 U902 ( .A(n807), .ZN(n815) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n867), .ZN(n917) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n868), .ZN(n924) );
  XOR2_X1 U905 ( .A(n983), .B(KEYINPUT107), .Z(n808) );
  NOR2_X1 U906 ( .A1(n924), .A2(n808), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n809), .A2(n932), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n917), .A2(n810), .ZN(n811) );
  XNOR2_X1 U909 ( .A(n811), .B(KEYINPUT108), .ZN(n812) );
  XNOR2_X1 U910 ( .A(n812), .B(KEYINPUT39), .ZN(n813) );
  NAND2_X1 U911 ( .A1(n813), .A2(n819), .ZN(n814) );
  OR2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  AND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n889), .A2(n818), .ZN(n933) );
  NAND2_X1 U915 ( .A1(n933), .A2(n819), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(KEYINPUT40), .B(n822), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U920 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(G188) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(G325) );
  XOR2_X1 U924 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  INV_X1 U927 ( .A(n829), .ZN(G319) );
  XNOR2_X1 U928 ( .A(G2078), .B(G2072), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n830), .B(KEYINPUT42), .ZN(n840) );
  XOR2_X1 U930 ( .A(G2678), .B(KEYINPUT43), .Z(n832) );
  XNOR2_X1 U931 ( .A(KEYINPUT112), .B(G2096), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U933 ( .A(G2100), .B(G2090), .Z(n834) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2084), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT113), .B(KEYINPUT111), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U940 ( .A(G1986), .B(G1961), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1976), .B(G1971), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n843), .B(KEYINPUT41), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(G2474), .B(G1956), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1981), .B(G1966), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n877), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n850), .B(KEYINPUT44), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n851), .B(KEYINPUT114), .ZN(n853) );
  NAND2_X1 U953 ( .A1(G112), .A2(n535), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U955 ( .A1(G136), .A2(n880), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G100), .A2(n881), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U958 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G127), .A2(n877), .ZN(n859) );
  NAND2_X1 U960 ( .A1(G115), .A2(n535), .ZN(n858) );
  NAND2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n860), .B(KEYINPUT47), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G139), .A2(n880), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n881), .A2(G103), .ZN(n863) );
  XOR2_X1 U966 ( .A(KEYINPUT116), .B(n863), .Z(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n928) );
  XOR2_X1 U968 ( .A(G160), .B(n928), .Z(n866) );
  XNOR2_X1 U969 ( .A(n921), .B(n866), .ZN(n871) );
  XNOR2_X1 U970 ( .A(G162), .B(n867), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U972 ( .A(n871), .B(n870), .Z(n876) );
  XOR2_X1 U973 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n873) );
  XNOR2_X1 U974 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U976 ( .A(KEYINPUT118), .B(n874), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n888) );
  NAND2_X1 U978 ( .A1(G130), .A2(n877), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G118), .A2(n535), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G142), .A2(n880), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G106), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n884), .Z(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U986 ( .A(n888), .B(n887), .Z(n891) );
  XNOR2_X1 U987 ( .A(n889), .B(G164), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U989 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U990 ( .A(G286), .B(G171), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n967), .B(n895), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U994 ( .A1(G37), .A2(n898), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2454), .B(G2435), .Z(n900) );
  XNOR2_X1 U996 ( .A(G2438), .B(G2427), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n907) );
  XOR2_X1 U998 ( .A(KEYINPUT109), .B(G2446), .Z(n902) );
  XNOR2_X1 U999 ( .A(G2443), .B(G2430), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n903), .B(G2451), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n908), .A2(G14), .ZN(n915) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n909) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n909), .Z(n910) );
  XNOR2_X1 U1009 ( .A(n910), .B(KEYINPUT119), .ZN(n911) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(n915), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n918), .B(KEYINPUT51), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n927) );
  XNOR2_X1 U1019 ( .A(G160), .B(G2084), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n925), .B(KEYINPUT120), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n937) );
  XOR2_X1 U1024 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(KEYINPUT50), .B(n931), .ZN(n935) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  INV_X1 U1032 ( .A(KEYINPUT55), .ZN(n960) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n960), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n940), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1035 ( .A(G2090), .B(G35), .ZN(n955) );
  XOR2_X1 U1036 ( .A(n941), .B(G27), .Z(n943) );
  XNOR2_X1 U1037 ( .A(G32), .B(G1996), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(KEYINPUT122), .B(n944), .ZN(n950) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1041 ( .A1(n945), .A2(G28), .ZN(n948) );
  XOR2_X1 U1042 ( .A(KEYINPUT121), .B(G2072), .Z(n946) );
  XNOR2_X1 U1043 ( .A(G33), .B(n946), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G26), .B(G2067), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n953), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1050 ( .A(G2084), .B(G34), .Z(n956) );
  XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(n960), .B(n959), .ZN(n962) );
  INV_X1 U1054 ( .A(G29), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n963), .ZN(n1020) );
  XNOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT57), .ZN(n988) );
  XNOR2_X1 U1061 ( .A(n967), .B(G1341), .ZN(n986) );
  XNOR2_X1 U1062 ( .A(G1956), .B(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n981) );
  XNOR2_X1 U1067 ( .A(G1348), .B(n975), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n979) );
  XOR2_X1 U1069 ( .A(G1961), .B(G171), .Z(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(KEYINPUT123), .B(n984), .ZN(n985) );
  NOR2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1076 ( .A1(n990), .A2(n989), .ZN(n1018) );
  INV_X1 U1077 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1078 ( .A(G1976), .B(G23), .Z(n992) );
  XOR2_X1 U1079 ( .A(G1971), .B(G22), .Z(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(G24), .B(G1986), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1083 ( .A(KEYINPUT58), .B(n995), .Z(n1013) );
  XNOR2_X1 U1084 ( .A(G1961), .B(G5), .ZN(n1010) );
  XOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .Z(n996) );
  XNOR2_X1 U1086 ( .A(G4), .B(n996), .ZN(n1004) );
  XOR2_X1 U1087 ( .A(G1981), .B(G6), .Z(n999) );
  XNOR2_X1 U1088 ( .A(n997), .B(G20), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G19), .B(G1341), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(KEYINPUT124), .B(n1002), .Z(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT125), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(KEYINPUT126), .B(n1011), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

