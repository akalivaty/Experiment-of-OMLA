//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G68), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n218), .A2(G238), .B1(G50), .B2(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n213), .B(new_n224), .C1(G116), .C2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  AOI22_X1  g0027(.A1(new_n225), .A2(new_n227), .B1(G1), .B2(G20), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n202), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n210), .B(new_n229), .C1(new_n232), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n244), .B(KEYINPUT68), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n230), .B1(new_n207), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT69), .Z(new_n256));
  INV_X1    g0056(.A(G50), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n231), .B1(new_n201), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT70), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n254), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n231), .A2(new_n254), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n260), .A2(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n256), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n257), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n255), .B(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n268), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n266), .B(new_n271), .C1(new_n257), .C2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT9), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G222), .A2(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G223), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n280), .B(new_n283), .C1(G77), .C2(new_n276), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G226), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n282), .A2(new_n285), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n284), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n275), .B(new_n292), .C1(new_n293), .C2(new_n291), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT77), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT77), .B1(new_n254), .B2(KEYINPUT3), .ZN(new_n301));
  OAI211_X1 g0101(.A(KEYINPUT7), .B(new_n231), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT7), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n276), .B2(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n218), .ZN(new_n306));
  INV_X1    g0106(.A(G159), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n264), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n215), .A2(new_n217), .A3(G58), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT76), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT76), .A4(G58), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n202), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n308), .B1(new_n313), .B2(G20), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT16), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(G20), .B1(new_n298), .B2(new_n297), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT75), .B1(new_n318), .B2(KEYINPUT7), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(KEYINPUT7), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n321), .B(new_n303), .C1(new_n276), .C2(G20), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G68), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n314), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n317), .A2(new_n256), .A3(new_n325), .ZN(new_n326));
  OR2_X1    g0126(.A1(G223), .A2(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n289), .A2(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n298), .A2(new_n327), .A3(new_n297), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G87), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n283), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n282), .A2(G232), .A3(new_n285), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n288), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT78), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n332), .A2(KEYINPUT78), .A3(new_n288), .A4(new_n334), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n282), .B1(new_n329), .B2(new_n330), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n341), .A2(new_n287), .A3(new_n333), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n293), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n260), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n270), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n273), .B2(new_n345), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n326), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(KEYINPUT79), .B2(KEYINPUT17), .ZN(new_n350));
  XOR2_X1   g0150(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n325), .A2(new_n256), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT16), .B1(new_n306), .B2(new_n314), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n348), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n335), .A2(G179), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n342), .A2(KEYINPUT78), .ZN(new_n358));
  NOR4_X1   g0158(.A1(new_n341), .A2(new_n336), .A3(new_n333), .A4(new_n287), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n356), .A2(new_n362), .A3(KEYINPUT18), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n353), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n291), .A2(new_n361), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n274), .B(new_n368), .C1(G179), .C2(new_n291), .ZN(new_n369));
  XOR2_X1   g0169(.A(KEYINPUT15), .B(G87), .Z(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n262), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n260), .A2(new_n264), .B1(new_n231), .B2(new_n220), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n256), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n272), .A2(G77), .A3(new_n268), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n270), .A2(new_n220), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n276), .A2(G238), .A3(G1698), .ZN(new_n379));
  INV_X1    g0179(.A(G107), .ZN(new_n380));
  INV_X1    g0180(.A(G232), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n276), .A2(new_n278), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n379), .B1(new_n380), .B2(new_n276), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n287), .B1(new_n383), .B2(new_n283), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n290), .A2(new_n221), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT71), .B(new_n378), .C1(new_n387), .C2(new_n338), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(G190), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT71), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n338), .B1(new_n384), .B2(new_n386), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n377), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n388), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n295), .A2(new_n367), .A3(new_n369), .A4(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n282), .A2(G238), .A3(new_n285), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G226), .A2(G1698), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n381), .B2(G1698), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n276), .B1(G33), .B2(G97), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n395), .B(new_n288), .C1(new_n398), .C2(new_n282), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT72), .ZN(new_n402));
  OR3_X1    g0202(.A1(new_n399), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n293), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n272), .A2(G68), .A3(new_n268), .ZN(new_n405));
  XOR2_X1   g0205(.A(new_n405), .B(KEYINPUT73), .Z(new_n406));
  INV_X1    g0206(.A(new_n264), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(G50), .B1(G77), .B2(new_n261), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n231), .B2(new_n218), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n256), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT11), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT12), .B1(new_n270), .B2(new_n214), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT12), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n218), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n412), .B1(new_n414), .B2(new_n270), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n338), .B1(new_n400), .B2(new_n401), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n404), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n404), .A2(new_n416), .A3(KEYINPUT74), .A4(new_n417), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n361), .B1(new_n400), .B2(new_n401), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G179), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n402), .B2(new_n403), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n416), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n387), .A2(new_n426), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n377), .C1(G169), .C2(new_n387), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n394), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G283), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n231), .C1(G33), .C2(new_n211), .ZN(new_n435));
  XOR2_X1   g0235(.A(KEYINPUT83), .B(G116), .Z(new_n436));
  OAI211_X1 g0236(.A(new_n255), .B(new_n435), .C1(new_n436), .C2(new_n231), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT20), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n270), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n254), .A2(G1), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT82), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n270), .B1(KEYINPUT82), .B2(new_n443), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n272), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n439), .B(new_n441), .C1(new_n442), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G41), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(G45), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(G1), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n453), .A2(new_n286), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n282), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G270), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n298), .A2(new_n297), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G303), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n276), .A2(G1698), .ZN(new_n459));
  INV_X1    g0259(.A(G264), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n457), .A2(G1698), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(G257), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n454), .B(new_n456), .C1(new_n463), .C2(new_n282), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n447), .A2(G169), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT21), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n464), .A2(new_n426), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n447), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n447), .A2(KEYINPUT21), .A3(G169), .A4(new_n464), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n276), .A2(new_n231), .A3(G87), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT22), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT22), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n276), .A2(new_n474), .A3(new_n231), .A4(G87), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n436), .A2(new_n261), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n231), .A2(G107), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT23), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT24), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n476), .A2(KEYINPUT24), .A3(new_n477), .A4(new_n479), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n256), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n446), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n270), .A2(new_n380), .ZN(new_n487));
  XOR2_X1   g0287(.A(new_n487), .B(KEYINPUT25), .Z(new_n488));
  NAND3_X1  g0288(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT85), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n459), .B2(new_n212), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n276), .A2(KEYINPUT85), .A3(G257), .A4(G1698), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G294), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n382), .A2(new_n223), .B1(new_n254), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n283), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n455), .A2(G264), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n426), .A3(new_n454), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(new_n454), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n361), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n489), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n464), .A2(G200), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n293), .B2(new_n464), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n504), .A2(new_n447), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n471), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n270), .A2(new_n211), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n485), .A2(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n305), .A2(G107), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n380), .A2(KEYINPUT6), .A3(G97), .ZN(new_n512));
  XOR2_X1   g0312(.A(G97), .B(G107), .Z(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(G20), .B1(G77), .B2(new_n407), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n305), .A2(KEYINPUT80), .A3(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n256), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n517), .B2(new_n256), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n507), .B(new_n508), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n462), .A2(KEYINPUT4), .A3(G244), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n382), .B2(new_n221), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n434), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n283), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n455), .A2(G257), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n528), .A2(new_n454), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n426), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT86), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n500), .A2(G200), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(new_n486), .A3(new_n488), .A4(new_n484), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n500), .A2(new_n293), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n539));
  INV_X1    g0339(.A(new_n537), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(KEYINPUT86), .A3(new_n540), .A4(new_n535), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n221), .A2(G1698), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n276), .B(new_n543), .C1(G238), .C2(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n436), .A2(G33), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n282), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(G274), .B2(new_n451), .ZN(new_n547));
  INV_X1    g0347(.A(new_n451), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(G250), .A3(new_n282), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n361), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n276), .A2(new_n231), .A3(G68), .ZN(new_n552));
  NAND3_X1  g0352(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n231), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n205), .B2(G87), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n262), .A2(new_n211), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n552), .B(new_n555), .C1(new_n556), .C2(KEYINPUT19), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n256), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n371), .A2(new_n270), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n446), .C2(new_n371), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n547), .A2(new_n426), .A3(new_n549), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n551), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n558), .A2(new_n559), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n446), .A2(new_n222), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n547), .A2(G190), .A3(new_n549), .ZN(new_n566));
  INV_X1    g0366(.A(new_n549), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n567), .B(new_n546), .C1(G274), .C2(new_n451), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n565), .B(new_n566), .C1(new_n568), .C2(new_n338), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n562), .A2(KEYINPUT84), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT84), .B1(new_n562), .B2(new_n569), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n521), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n519), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n530), .A2(new_n293), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G200), .B2(new_n530), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n574), .A2(new_n576), .A3(new_n507), .A4(new_n508), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n533), .A2(new_n542), .A3(new_n572), .A4(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n433), .A2(new_n506), .A3(new_n578), .ZN(G372));
  INV_X1    g0379(.A(new_n430), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n422), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n353), .B1(new_n581), .B2(new_n428), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT88), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n356), .A2(KEYINPUT18), .A3(new_n362), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT18), .B1(new_n356), .B2(new_n362), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n365), .A2(KEYINPUT88), .A3(new_n366), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n295), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n589), .A2(new_n369), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n533), .A2(new_n577), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n471), .A2(new_n502), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(new_n542), .A3(new_n569), .A4(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n551), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n551), .A2(new_n561), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n560), .B(new_n595), .C1(new_n596), .C2(new_n594), .ZN(new_n597));
  INV_X1    g0397(.A(new_n533), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n572), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT26), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n569), .ZN(new_n601));
  OR3_X1    g0401(.A1(new_n601), .A2(new_n533), .A3(KEYINPUT26), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n593), .A2(new_n597), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n432), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n590), .A2(new_n604), .ZN(G369));
  NAND2_X1  g0405(.A1(new_n471), .A2(new_n505), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT90), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n269), .A2(G20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n267), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n609), .A2(KEYINPUT27), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(KEYINPUT27), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(G213), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(G343), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n447), .A2(new_n614), .ZN(new_n615));
  OR3_X1    g0415(.A1(new_n607), .A2(KEYINPUT89), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n607), .B1(KEYINPUT89), .B2(new_n615), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(G330), .ZN(new_n618));
  INV_X1    g0418(.A(new_n502), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n489), .A2(new_n614), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n542), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n502), .A2(new_n614), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n471), .A2(new_n614), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n622), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(G399));
  INV_X1    g0429(.A(new_n208), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(G41), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G1), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n233), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT28), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT29), .ZN(new_n637));
  INV_X1    g0437(.A(new_n614), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n603), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n578), .A2(new_n506), .A3(new_n614), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n528), .A2(new_n529), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(new_n568), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(KEYINPUT30), .A3(new_n498), .A4(new_n468), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n468), .A2(new_n498), .A3(new_n568), .A4(new_n641), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT30), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n500), .A2(new_n550), .ZN(new_n647));
  INV_X1    g0447(.A(new_n530), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(new_n426), .A4(new_n464), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n643), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n614), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT31), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(KEYINPUT31), .A3(new_n614), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(G330), .B1(new_n640), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT26), .B1(new_n601), .B2(new_n533), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n599), .B2(KEYINPUT26), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n592), .A2(new_n542), .A3(new_n569), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n533), .A2(new_n577), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n597), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n614), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n639), .B(new_n656), .C1(new_n663), .C2(new_n637), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n636), .B1(new_n665), .B2(G1), .ZN(G364));
  AND2_X1   g0466(.A1(new_n616), .A2(new_n617), .ZN(new_n667));
  NOR2_X1   g0467(.A1(G13), .A2(G33), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n231), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n608), .A2(G45), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n632), .A2(G1), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n249), .A2(G45), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT92), .Z(new_n675));
  NOR2_X1   g0475(.A1(new_n630), .A2(new_n276), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(G45), .B2(new_n233), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n675), .A2(new_n677), .B1(G116), .B2(new_n208), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n630), .A2(new_n457), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT91), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n678), .B1(G355), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n669), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n230), .B1(G20), .B2(new_n361), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n231), .A2(new_n293), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n338), .A2(G179), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n276), .B1(new_n689), .B2(G303), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n231), .A2(G190), .ZN(new_n691));
  NOR2_X1   g0491(.A1(G179), .A2(G200), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G329), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n426), .A2(G200), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n686), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G322), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n690), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n231), .B1(new_n692), .B2(G190), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT95), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT95), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n691), .A2(new_n687), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT94), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n705), .A2(G294), .B1(G283), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G326), .ZN(new_n709));
  NAND3_X1  g0509(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT93), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n293), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n708), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n711), .A2(G190), .ZN(new_n715));
  XNOR2_X1  g0515(.A(KEYINPUT33), .B(G317), .ZN(new_n716));
  AOI211_X1 g0516(.A(new_n700), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n691), .A2(new_n696), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G311), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n705), .A2(G97), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(G77), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT32), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n694), .B2(G159), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(G87), .B2(new_n689), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n694), .A2(new_n723), .A3(G159), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n721), .A2(new_n722), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(G50), .A2(new_n712), .B1(new_n715), .B2(G68), .ZN(new_n728));
  INV_X1    g0528(.A(G58), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n729), .B2(new_n697), .ZN(new_n730));
  INV_X1    g0530(.A(new_n707), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n380), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n727), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n717), .A2(new_n720), .B1(new_n276), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT96), .ZN(new_n735));
  INV_X1    g0535(.A(new_n683), .ZN(new_n736));
  OAI221_X1 g0536(.A(new_n673), .B1(new_n681), .B2(new_n685), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n667), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n618), .A2(new_n672), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n670), .A2(new_n737), .B1(new_n738), .B2(new_n739), .ZN(G396));
  NAND2_X1  g0540(.A1(new_n603), .A2(new_n638), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n393), .B1(new_n378), .B2(new_n638), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n430), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n580), .A2(new_n638), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n745), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n603), .A2(new_n638), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G330), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n653), .A2(new_n654), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n533), .A2(new_n572), .A3(new_n577), .ZN(new_n752));
  INV_X1    g0552(.A(new_n506), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(new_n542), .A4(new_n638), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n749), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n672), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n745), .A2(new_n668), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G137), .A2(new_n712), .B1(new_n715), .B2(G150), .ZN(new_n759));
  INV_X1    g0559(.A(G143), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n759), .B1(new_n760), .B2(new_n697), .C1(new_n307), .C2(new_n718), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT34), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n707), .A2(G68), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n688), .A2(new_n257), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n457), .B(new_n764), .C1(G132), .C2(new_n694), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n704), .A2(new_n729), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n731), .A2(new_n222), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  INV_X1    g0569(.A(new_n715), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n721), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n768), .B(new_n771), .C1(G311), .C2(new_n694), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n712), .A2(G303), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n719), .A2(new_n436), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n276), .B1(new_n689), .B2(G107), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n772), .A2(new_n773), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n697), .A2(new_n494), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n766), .A2(new_n767), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n683), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n683), .A2(new_n668), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n220), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n758), .A2(new_n673), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n757), .A2(new_n782), .ZN(G384));
  NAND2_X1  g0583(.A1(new_n751), .A2(new_n754), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n428), .B1(new_n420), .B2(new_n421), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n416), .A2(new_n614), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n428), .B(new_n786), .C1(new_n420), .C2(new_n421), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n745), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT103), .ZN(new_n792));
  NOR2_X1   g0592(.A1(KEYINPUT79), .A2(KEYINPUT17), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n325), .A2(new_n256), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n347), .B1(new_n794), .B2(new_n317), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n793), .B1(new_n795), .B2(new_n344), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n349), .A2(new_n351), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n797), .B1(new_n584), .B2(new_n585), .ZN(new_n798));
  INV_X1    g0598(.A(new_n612), .ZN(new_n799));
  AOI21_X1  g0599(.A(KEYINPUT16), .B1(new_n324), .B2(new_n314), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n348), .B1(new_n354), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n358), .A2(G169), .A3(new_n359), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n612), .B1(new_n803), .B2(new_n357), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n801), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n805), .A2(KEYINPUT37), .A3(new_n349), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT37), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n356), .A2(new_n799), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n363), .A2(new_n808), .A3(new_n349), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g0610(.A1(new_n802), .A2(KEYINPUT38), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(KEYINPUT38), .B1(new_n802), .B2(new_n810), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT103), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n784), .A2(new_n814), .A3(new_n790), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n792), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n808), .A2(new_n583), .A3(new_n349), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(KEYINPUT37), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n809), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n808), .A2(new_n349), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n823), .A2(KEYINPUT88), .A3(KEYINPUT37), .A4(new_n363), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n808), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n352), .A2(new_n586), .A3(new_n587), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT100), .B1(new_n828), .B2(KEYINPUT38), .ZN(new_n829));
  INV_X1    g0629(.A(new_n811), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT100), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n827), .A2(new_n826), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n831), .B(new_n832), .C1(new_n834), .C2(new_n825), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n829), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n836), .A2(KEYINPUT40), .A3(new_n784), .A4(new_n790), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n819), .A2(new_n837), .A3(G330), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n432), .A2(new_n755), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n819), .A2(new_n784), .A3(new_n837), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n433), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n663), .A2(new_n637), .ZN(new_n843));
  INV_X1    g0643(.A(new_n639), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n432), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n590), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n842), .B(new_n846), .Z(new_n847));
  NOR2_X1   g0647(.A1(new_n428), .A2(new_n614), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT39), .B1(new_n811), .B2(new_n812), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT99), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(KEYINPUT99), .B(KEYINPUT39), .C1(new_n811), .C2(new_n812), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT39), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n829), .A2(new_n835), .A3(new_n854), .A4(new_n830), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n853), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT101), .B1(new_n853), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n848), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n748), .A2(new_n744), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n788), .A2(new_n789), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n863), .A2(new_n813), .B1(new_n588), .B2(new_n612), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n847), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n267), .B2(new_n608), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n311), .A2(new_n234), .A3(G77), .A4(new_n312), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(G50), .B2(new_n214), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(G1), .A3(new_n269), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n514), .B(KEYINPUT97), .Z(new_n871));
  AOI21_X1  g0671(.A(new_n442), .B1(new_n871), .B2(KEYINPUT35), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n872), .B(new_n232), .C1(KEYINPUT35), .C2(new_n871), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT98), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT36), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n867), .A2(new_n870), .A3(new_n875), .ZN(G367));
  AOI21_X1  g0676(.A(new_n685), .B1(new_n244), .B2(new_n676), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n370), .A2(new_n630), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n672), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n712), .A2(G311), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n880), .B1(new_n704), .B2(new_n380), .C1(new_n770), .C2(new_n494), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT46), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n688), .A2(new_n882), .A3(new_n442), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n440), .B2(new_n688), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n884), .B(new_n457), .C1(new_n769), .C2(new_n718), .ZN(new_n885));
  INV_X1    g0685(.A(new_n706), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n883), .B(new_n885), .C1(G97), .C2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(G303), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n888), .B2(new_n697), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n881), .B(new_n889), .C1(G317), .C2(new_n694), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n457), .B1(new_n694), .B2(G137), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n891), .B1(new_n257), .B2(new_n718), .C1(new_n713), .C2(new_n760), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n705), .A2(G68), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n698), .A2(G150), .B1(new_n886), .B2(G77), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n893), .B(new_n894), .C1(new_n307), .C2(new_n770), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n892), .B(new_n895), .C1(G58), .C2(new_n689), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT47), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n879), .B1(new_n898), .B2(new_n736), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT109), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n565), .A2(new_n638), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n597), .A2(new_n569), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n597), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n900), .B1(new_n669), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n671), .A2(G1), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n522), .A2(new_n614), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n660), .A2(new_n908), .B1(new_n533), .B2(new_n638), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n628), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT45), .Z(new_n911));
  NOR2_X1   g0711(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n912));
  OR3_X1    g0712(.A1(new_n628), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n628), .B2(new_n909), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n625), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n623), .B(new_n627), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n618), .B(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(new_n664), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n911), .A2(new_n626), .A3(new_n916), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT107), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT107), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n918), .A2(new_n921), .A3(new_n925), .A4(new_n922), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n664), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n631), .B(KEYINPUT41), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n907), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n909), .B(KEYINPUT104), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n502), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n638), .B1(new_n932), .B2(new_n598), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n623), .A2(new_n909), .A3(new_n627), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT42), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(KEYINPUT105), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(KEYINPUT105), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n904), .B(KEYINPUT43), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n937), .B2(new_n939), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n941), .A2(new_n943), .B1(new_n626), .B2(new_n931), .ZN(new_n944));
  INV_X1    g0744(.A(new_n943), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n626), .A2(new_n931), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(new_n940), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT108), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n930), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n930), .B2(new_n948), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n905), .B1(new_n951), .B2(new_n952), .ZN(G387));
  AND2_X1   g0753(.A1(new_n920), .A2(new_n664), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n954), .A2(new_n921), .A3(new_n632), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G159), .A2(new_n712), .B1(new_n715), .B2(new_n345), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n257), .B2(new_n697), .C1(new_n211), .C2(new_n731), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G68), .B2(new_n719), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n705), .A2(new_n370), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n688), .A2(new_n220), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G150), .B2(new_n694), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n958), .A2(new_n276), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G311), .A2(new_n715), .B1(new_n712), .B2(G322), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n888), .B2(new_n718), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G317), .B2(new_n698), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT48), .Z(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n769), .B2(new_n704), .C1(new_n494), .C2(new_n688), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n457), .B1(new_n693), .B2(new_n709), .C1(new_n440), .C2(new_n706), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n962), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n683), .ZN(new_n972));
  AOI21_X1  g0772(.A(G45), .B1(G68), .B2(G77), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n345), .A2(new_n257), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n633), .B(new_n973), .C1(new_n974), .C2(KEYINPUT50), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(KEYINPUT50), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n676), .B1(new_n241), .B2(new_n450), .ZN(new_n977));
  INV_X1    g0777(.A(new_n633), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n680), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n208), .A2(G107), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n684), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n624), .A2(new_n682), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n972), .A2(new_n673), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n955), .B(new_n984), .C1(new_n907), .C2(new_n920), .ZN(G393));
  NAND2_X1  g0785(.A1(new_n924), .A2(new_n926), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n918), .A2(KEYINPUT111), .A3(new_n922), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(KEYINPUT111), .B2(new_n922), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n631), .C1(new_n921), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n906), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n712), .A2(G317), .B1(G311), .B2(new_n698), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT52), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n276), .B(new_n732), .C1(G322), .C2(new_n694), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n769), .B2(new_n688), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT114), .Z(new_n995));
  AOI211_X1 g0795(.A(new_n992), .B(new_n995), .C1(G294), .C2(new_n719), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n888), .B2(new_n770), .C1(new_n440), .C2(new_n704), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT115), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n712), .A2(G150), .B1(G159), .B2(new_n698), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT51), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n718), .A2(new_n260), .B1(new_n693), .B2(new_n760), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n457), .B1(new_n705), .B2(G77), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n689), .A2(new_n218), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n768), .B1(G50), .B2(new_n715), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT113), .Z(new_n1007));
  OAI21_X1  g0807(.A(new_n683), .B1(new_n998), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n676), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n684), .B1(new_n211), .B2(new_n208), .C1(new_n252), .C2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT112), .Z(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n673), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT116), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1012), .A2(new_n1013), .B1(new_n682), .B2(new_n931), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n989), .A2(new_n990), .A3(new_n1015), .ZN(G390));
  INV_X1    g0816(.A(new_n857), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n853), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n668), .A3(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n705), .A2(G159), .B1(G128), .B2(new_n712), .ZN(new_n1020));
  INV_X1    g0820(.A(G137), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n770), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n688), .A2(new_n263), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT53), .Z(new_n1024));
  AOI211_X1 g0824(.A(new_n457), .B(new_n1024), .C1(G132), .C2(new_n698), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT54), .B(G143), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1025), .B1(new_n257), .B2(new_n706), .C1(new_n718), .C2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1022), .B(new_n1028), .C1(G125), .C2(new_n694), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G87), .A2(new_n689), .B1(new_n698), .B2(G116), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n276), .B1(new_n694), .B2(G294), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n763), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n705), .A2(G77), .B1(G283), .B2(new_n712), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n380), .B2(new_n770), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(G97), .C2(new_n719), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n683), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n780), .A2(new_n260), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1019), .A2(new_n673), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n784), .A2(G330), .A3(new_n790), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n848), .B1(new_n859), .B2(new_n861), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n856), .A2(new_n857), .A3(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n638), .B(new_n743), .C1(new_n658), .C2(new_n661), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n744), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n848), .B1(new_n1044), .B2(new_n861), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n836), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1040), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1041), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1017), .A2(new_n1049), .A3(new_n1018), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(new_n1039), .A3(new_n1046), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n906), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT120), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1048), .A2(new_n1051), .A3(KEYINPUT120), .A4(new_n906), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n845), .A2(new_n839), .A3(new_n590), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT118), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n745), .B1(new_n656), .B2(KEYINPUT117), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT117), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n755), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n861), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1039), .A2(new_n1043), .A3(new_n744), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1058), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n747), .B1(new_n755), .B2(new_n1060), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n656), .A2(KEYINPUT117), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n862), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1063), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(KEYINPUT118), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n861), .B1(new_n755), .B2(new_n747), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n859), .B1(new_n1071), .B2(new_n1040), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1057), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1048), .A2(new_n1073), .A3(new_n1051), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT119), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n631), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1038), .B(new_n1056), .C1(new_n1077), .C2(new_n1078), .ZN(G378));
  NAND2_X1  g0879(.A1(new_n295), .A2(new_n369), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n274), .A2(new_n799), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1082), .B(new_n1083), .Z(new_n1084));
  NAND2_X1  g0884(.A1(new_n838), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1084), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1086), .A2(new_n819), .A3(G330), .A4(new_n837), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n865), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1085), .A2(new_n858), .A3(new_n864), .A4(new_n1087), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n906), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n672), .B1(new_n1084), .B2(new_n668), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n780), .A2(new_n257), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G125), .A2(new_n712), .B1(new_n715), .B2(G132), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G128), .A2(new_n698), .B1(new_n719), .B2(G137), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n688), .C2(new_n1027), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G150), .B2(new_n705), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT59), .ZN(new_n1099));
  OR2_X1    g0899(.A1(KEYINPUT121), .A2(G124), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(KEYINPUT121), .A2(G124), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n694), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(G33), .B1(new_n886), .B2(G159), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n448), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n371), .A2(new_n718), .B1(new_n380), .B2(new_n697), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n893), .B(new_n448), .C1(new_n442), .C2(new_n713), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G58), .C2(new_n886), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n276), .B(new_n960), .C1(G283), .C2(new_n694), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n211), .C2(new_n770), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT58), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1104), .B(new_n1111), .C1(G50), .C2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n683), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT122), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1093), .A2(new_n1094), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1092), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1057), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1074), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1089), .A2(KEYINPUT123), .A3(new_n1090), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT123), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1088), .A2(new_n865), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT57), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1074), .A2(new_n1120), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n631), .B1(new_n1127), .B2(KEYINPUT57), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1119), .B1(new_n1126), .B2(new_n1128), .ZN(G375));
  AND2_X1   g0929(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n959), .B1(new_n888), .B2(new_n693), .C1(new_n440), .C2(new_n770), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G294), .B2(new_n712), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n731), .A2(new_n220), .B1(new_n380), .B2(new_n718), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n276), .B(new_n1134), .C1(G97), .C2(new_n689), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(new_n769), .C2(new_n697), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n770), .A2(new_n1027), .B1(new_n704), .B2(new_n257), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n697), .A2(new_n1021), .B1(new_n718), .B2(new_n263), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n689), .A2(G159), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n457), .B1(new_n886), .B2(G58), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n712), .A2(G132), .B1(G128), .B2(new_n694), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n736), .B1(new_n1136), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n672), .B(new_n1144), .C1(new_n214), .C2(new_n780), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n862), .A2(new_n668), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT124), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1131), .A2(new_n906), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1130), .A2(new_n1057), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1073), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n928), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1151), .ZN(G381));
  NAND2_X1  g0952(.A1(new_n1121), .A2(new_n1091), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT57), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n632), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1118), .B1(new_n1155), .B2(new_n1125), .ZN(new_n1156));
  INV_X1    g0956(.A(G378), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1158), .A2(G384), .A3(G381), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(G387), .A2(G390), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(G393), .A2(G396), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(G407));
  OAI211_X1 g0962(.A(G407), .B(G213), .C1(G343), .C2(new_n1158), .ZN(G409));
  XOR2_X1   g0963(.A(G393), .B(G396), .Z(new_n1164));
  INV_X1    g0964(.A(G390), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n930), .A2(new_n948), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT108), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n950), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1165), .B1(new_n1168), .B2(new_n905), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1164), .B1(new_n1160), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(G387), .A2(G390), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n905), .A3(new_n1165), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1164), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1127), .A2(new_n928), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1122), .A2(new_n906), .A3(new_n1124), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1176), .A2(new_n1117), .A3(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(G378), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT125), .B1(G375), .B2(new_n1157), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1155), .A2(new_n1125), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT125), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1181), .A2(new_n1182), .A3(G378), .A4(new_n1119), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1179), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(G213), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(G343), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT60), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1149), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n1057), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1188), .A2(new_n631), .A3(new_n1150), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1148), .ZN(new_n1191));
  INV_X1    g0991(.A(G384), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(G384), .A3(new_n1148), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1184), .A2(new_n1186), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT62), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT61), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1197), .B2(new_n1196), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(G2897), .A3(new_n1186), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1186), .A2(G2897), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1193), .A2(new_n1194), .A3(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1175), .B1(new_n1199), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT61), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1196), .B2(KEYINPUT63), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1183), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1182), .B1(new_n1156), .B2(G378), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1209), .A2(new_n1210), .B1(G378), .B2(new_n1178), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1186), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1195), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(KEYINPUT63), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1173), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1208), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1204), .A2(KEYINPUT126), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT126), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n1203), .C1(new_n1184), .C2(new_n1186), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT127), .B1(new_n1219), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1175), .B1(new_n1196), .B2(KEYINPUT63), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT63), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT61), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AND4_X1   g1028(.A1(KEYINPUT127), .A2(new_n1223), .A3(new_n1225), .A4(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1206), .B1(new_n1224), .B2(new_n1229), .ZN(G405));
  OAI22_X1  g1030(.A1(new_n1209), .A2(new_n1210), .B1(G378), .B2(new_n1156), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1175), .B(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(new_n1213), .ZN(G402));
endmodule


