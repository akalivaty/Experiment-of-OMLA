//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930;
  XOR2_X1   g000(.A(G110), .B(G140), .Z(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT87), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT0), .A4(G128), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n197), .B(KEYINPUT65), .ZN(new_n198));
  OR3_X1    g012(.A1(new_n193), .A2(KEYINPUT64), .A3(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(KEYINPUT64), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n194), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT0), .B(G128), .Z(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n198), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT88), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n207), .A2(new_n210), .A3(new_n214), .A4(new_n211), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(G101), .A3(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n216), .A2(KEYINPUT4), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n212), .A2(G101), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n205), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n194), .A2(new_n196), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(KEYINPUT1), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n202), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n211), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n206), .A2(G107), .ZN(new_n229));
  OAI21_X1  g043(.A(G101), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n218), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n232), .A3(KEYINPUT10), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n220), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT11), .ZN(new_n236));
  INV_X1    g050(.A(G134), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n240), .B(new_n236), .C1(new_n237), .C2(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G134), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n237), .A2(KEYINPUT67), .A3(G137), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n237), .A2(G137), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n246), .A2(new_n247), .B1(new_n248), .B2(KEYINPUT11), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n242), .A2(new_n249), .A3(new_n252), .A4(new_n243), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n242), .A2(new_n249), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n251), .A2(new_n253), .B1(G131), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT10), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n223), .B1(new_n225), .B2(new_n221), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n231), .B2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n234), .A2(new_n235), .A3(new_n255), .A4(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n220), .A2(new_n255), .A3(new_n258), .A4(new_n233), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT89), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT90), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n226), .A2(new_n231), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n231), .B2(new_n257), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n251), .A2(new_n253), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n254), .A2(G131), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n264), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n263), .A2(KEYINPUT90), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n266), .A2(new_n269), .A3(KEYINPUT90), .A4(new_n263), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n192), .B1(new_n262), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n220), .A2(new_n258), .A3(new_n233), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n269), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n260), .A2(KEYINPUT89), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n260), .A2(KEYINPUT89), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n192), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT91), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n191), .B1(new_n259), .B2(new_n261), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT91), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n276), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G469), .B1(new_n287), .B2(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT92), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT92), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n290), .B(G469), .C1(new_n287), .C2(G902), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n260), .B(new_n235), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n191), .B1(new_n292), .B2(new_n279), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n262), .A2(new_n275), .A3(new_n192), .ZN(new_n294));
  AOI211_X1 g108(.A(G469), .B(G902), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n289), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT9), .B(G234), .Z(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n300), .A2(G221), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n226), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n198), .B2(new_n204), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT95), .ZN(new_n308));
  INV_X1    g122(.A(G224), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G953), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n306), .A2(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT7), .B1(new_n309), .B2(G953), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n311), .B(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G116), .B(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G116), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n315), .B(G113), .C1(KEYINPUT5), .C2(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT2), .B(G113), .Z(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n314), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n321), .A2(new_n231), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT94), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(new_n321), .B2(new_n231), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G122), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n326), .B(KEYINPUT93), .Z(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT8), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n232), .A2(new_n323), .A3(new_n320), .A4(new_n318), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n319), .A2(new_n314), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n320), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n217), .A2(new_n332), .A3(new_n219), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n322), .A3(new_n327), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(G902), .B1(new_n313), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n322), .ZN(new_n337));
  INV_X1    g151(.A(new_n327), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT6), .A3(new_n334), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n305), .B1(new_n205), .B2(new_n304), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(new_n310), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n337), .A2(new_n343), .A3(new_n338), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G210), .B1(G237), .B2(G902), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n336), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n336), .B2(new_n345), .ZN(new_n348));
  OR3_X1    g162(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT96), .ZN(new_n349));
  OAI21_X1  g163(.A(G214), .B1(G237), .B2(G902), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(KEYINPUT96), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT97), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(G237), .A2(G953), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G214), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT98), .A3(G143), .ZN(new_n357));
  OR2_X1    g171(.A1(KEYINPUT98), .A2(G143), .ZN(new_n358));
  NAND2_X1  g172(.A1(KEYINPUT98), .A2(G143), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n358), .A2(G214), .A3(new_n355), .A4(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n360), .A3(G131), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT99), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n360), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n243), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n362), .B(new_n364), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n304), .A2(KEYINPUT16), .A3(G140), .ZN(new_n366));
  XNOR2_X1  g180(.A(G125), .B(G140), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(KEYINPUT16), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G146), .ZN(new_n369));
  NOR2_X1   g183(.A1(KEYINPUT100), .A2(KEYINPUT19), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT100), .A2(KEYINPUT19), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n193), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n365), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n361), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT18), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT18), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n363), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n367), .B(new_n193), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n377), .A2(new_n379), .A3(new_n380), .A4(new_n364), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n206), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n368), .B(G146), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n376), .A2(KEYINPUT17), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n388), .B(new_n389), .C1(new_n365), .C2(KEYINPUT17), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n384), .A3(new_n381), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G475), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n299), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n391), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n384), .B1(new_n390), .B2(new_n381), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n299), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G475), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n392), .A2(KEYINPUT20), .A3(new_n393), .A4(new_n299), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT81), .B(G217), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n298), .A2(new_n189), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G122), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G116), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT101), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n406), .A2(G116), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G107), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n209), .B1(new_n408), .B2(new_n409), .ZN(new_n412));
  XNOR2_X1  g226(.A(G128), .B(G143), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT102), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n414), .A2(KEYINPUT13), .B1(new_n222), .B2(G143), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n414), .B2(KEYINPUT13), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n416), .B2(G134), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n416), .A2(G134), .A3(new_n413), .ZN(new_n418));
  OAI22_X1  g232(.A1(new_n411), .A2(new_n412), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n408), .A2(KEYINPUT14), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n410), .A2(new_n420), .A3(G107), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n413), .B(new_n237), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n408), .B(new_n409), .C1(KEYINPUT14), .C2(new_n209), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n424), .A3(KEYINPUT103), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT103), .B1(new_n419), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n405), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n404), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT15), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G478), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n430), .B(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n402), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G952), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(G953), .ZN(new_n436));
  NAND2_X1  g250(.A1(G234), .A2(G237), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT21), .B(G898), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(G902), .A3(G953), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n439), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n446), .B(KEYINPUT104), .Z(new_n447));
  NAND3_X1  g261(.A1(new_n303), .A2(new_n354), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n245), .A2(G134), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(KEYINPUT70), .B2(new_n248), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n243), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n267), .A2(new_n454), .A3(new_n227), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n198), .A2(new_n204), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n255), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT30), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT71), .B1(new_n267), .B2(new_n454), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT71), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n461), .B(new_n453), .C1(new_n251), .C2(new_n253), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n205), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT69), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n255), .B2(new_n456), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n463), .A2(new_n227), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n332), .B(new_n459), .C1(new_n467), .C2(KEYINPUT30), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n332), .B(KEYINPUT72), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n457), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n472));
  NAND2_X1  g286(.A1(new_n355), .A2(G210), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT26), .B(G101), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n468), .A2(KEYINPUT74), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT74), .B1(new_n468), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT31), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT31), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n468), .A2(new_n482), .A3(new_n478), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n485));
  INV_X1    g299(.A(new_n332), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n467), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n471), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n464), .A2(new_n466), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n460), .A2(new_n462), .A3(new_n226), .ZN(new_n490));
  OAI211_X1 g304(.A(KEYINPUT76), .B(new_n332), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(KEYINPUT75), .B(KEYINPUT28), .Z(new_n493));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n458), .A2(KEYINPUT77), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n458), .A2(KEYINPUT77), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n469), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(new_n476), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT78), .B1(new_n484), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(G472), .A2(G902), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(new_n493), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n494), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n477), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT78), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n481), .A4(new_n483), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT32), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT32), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n500), .A2(new_n510), .A3(new_n507), .A4(new_n501), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT80), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT29), .B1(new_n498), .B2(new_n476), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n476), .B1(new_n468), .B2(new_n488), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n457), .A2(new_n470), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n488), .A2(KEYINPUT79), .A3(new_n518), .ZN(new_n519));
  OR3_X1    g333(.A1(new_n458), .A2(KEYINPUT79), .A3(new_n469), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT28), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n503), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n476), .A2(KEYINPUT29), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n299), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n513), .B(G472), .C1(new_n517), .C2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n514), .B2(new_n516), .ZN(new_n526));
  INV_X1    g340(.A(G472), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT80), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n512), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n316), .A2(G128), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT82), .B1(new_n531), .B2(KEYINPUT23), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n222), .A2(G119), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G110), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n533), .A2(new_n531), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT24), .B(G110), .Z(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n387), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT83), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n534), .A2(G110), .B1(new_n536), .B2(new_n537), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n367), .A2(new_n193), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n369), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT84), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT22), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(G137), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n544), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n299), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT85), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT25), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n403), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(G234), .B2(new_n299), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(KEYINPUT85), .A3(KEYINPUT25), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(G902), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n549), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT86), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT86), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n449), .A2(new_n530), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(G101), .ZN(G3));
  NAND3_X1  g380(.A1(new_n500), .A2(new_n299), .A3(new_n507), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G472), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n564), .A3(new_n508), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n297), .A2(new_n302), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n350), .B1(new_n347), .B2(new_n348), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT105), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT105), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n574), .B(new_n350), .C1(new_n347), .C2(new_n348), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n445), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n428), .A2(new_n579), .A3(new_n429), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT106), .B1(new_n419), .B2(new_n424), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n404), .ZN(new_n582));
  AOI211_X1 g396(.A(KEYINPUT106), .B(new_n405), .C1(new_n419), .C2(new_n424), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT33), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(G478), .A3(new_n299), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n430), .A2(G478), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n402), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n578), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n571), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT34), .B(G104), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G6));
  INV_X1    g407(.A(new_n402), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n433), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n578), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n571), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G107), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G9));
  NAND2_X1  g413(.A1(new_n568), .A2(new_n508), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n548), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n544), .B(new_n602), .Z(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n558), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(KEYINPUT107), .Z(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n557), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n448), .A2(new_n600), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT37), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G110), .ZN(G12));
  AOI21_X1  g424(.A(new_n607), .B1(new_n512), .B2(new_n529), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n442), .A2(G900), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n595), .B1(new_n438), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n570), .A2(new_n576), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G128), .ZN(G30));
  NOR2_X1   g430(.A1(new_n479), .A2(new_n480), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n519), .A2(new_n520), .A3(new_n477), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n299), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n509), .A2(new_n511), .B1(new_n619), .B2(G472), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n402), .A2(new_n433), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n349), .A2(new_n351), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT38), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n612), .A2(new_n438), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n625), .B(KEYINPUT39), .Z(new_n626));
  NOR2_X1   g440(.A1(new_n570), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n606), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT40), .B1(new_n570), .B2(new_n626), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n624), .A2(new_n350), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G143), .ZN(G45));
  NAND3_X1  g446(.A1(new_n402), .A2(new_n588), .A3(new_n625), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n530), .A2(new_n606), .A3(new_n614), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G146), .ZN(G48));
  INV_X1    g450(.A(G469), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n293), .A2(new_n294), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(new_n299), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n295), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n301), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n530), .A2(new_n590), .A3(new_n564), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT108), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT41), .B(G113), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G15));
  NAND4_X1  g460(.A1(new_n530), .A2(new_n596), .A3(new_n564), .A4(new_n642), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G116), .ZN(G18));
  NAND4_X1  g462(.A1(new_n640), .A2(new_n573), .A3(new_n302), .A4(new_n575), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n530), .A2(new_n447), .A3(new_n606), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G119), .ZN(G21));
  INV_X1    g466(.A(new_n560), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n522), .A2(new_n477), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n481), .A2(new_n483), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n501), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n568), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n658));
  OR3_X1    g472(.A1(new_n576), .A2(new_n658), .A3(new_n621), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n658), .B1(new_n576), .B2(new_n621), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n657), .A2(new_n445), .A3(new_n642), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G122), .ZN(G24));
  INV_X1    g477(.A(KEYINPUT110), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n633), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n649), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n568), .A2(new_n606), .A3(new_n666), .A4(new_n656), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT111), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n567), .A2(G472), .B1(new_n501), .B2(new_n655), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n606), .A4(new_n666), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G125), .ZN(G27));
  AOI22_X1  g487(.A1(new_n509), .A2(new_n511), .B1(new_n528), .B2(new_n525), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n276), .A2(KEYINPUT112), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n191), .B1(new_n292), .B2(new_n274), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT112), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n284), .A2(new_n286), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(G469), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT113), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n679), .A2(KEYINPUT113), .A3(G469), .A4(new_n680), .ZN(new_n684));
  NAND2_X1  g498(.A1(G469), .A2(G902), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n296), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n665), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n302), .A2(new_n350), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n622), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT42), .A4(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n674), .A2(new_n560), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n686), .A2(new_n690), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n530), .A2(new_n694), .A3(new_n564), .A4(new_n687), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n243), .ZN(G33));
  INV_X1    g512(.A(new_n564), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n674), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n613), .A3(new_n694), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT114), .B(G134), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G36));
  INV_X1    g517(.A(new_n588), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n402), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT43), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n600), .A2(new_n606), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n278), .B1(new_n285), .B2(KEYINPUT91), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n282), .A2(new_n283), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n676), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n680), .A2(new_n678), .A3(new_n675), .A4(KEYINPUT45), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n714), .A3(G469), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n685), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT46), .B1(new_n715), .B2(new_n685), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n717), .A3(new_n295), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n718), .A2(new_n301), .A3(new_n626), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n708), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n622), .A2(new_n350), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n707), .B2(KEYINPUT44), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G137), .ZN(G39));
  NOR3_X1   g539(.A1(new_n530), .A2(new_n564), .A3(new_n721), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n718), .B2(new_n301), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n715), .A2(new_n685), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n685), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n296), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n302), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n726), .A2(new_n634), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G140), .ZN(G42));
  NAND2_X1  g551(.A1(new_n619), .A2(G472), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n512), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n301), .B1(new_n659), .B2(new_n660), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n686), .A2(new_n607), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n625), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n615), .A2(new_n635), .A3(new_n672), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n611), .B(new_n614), .C1(new_n613), .C2(new_n634), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(KEYINPUT52), .A3(new_n672), .A4(new_n742), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  OR3_X1    g562(.A1(new_n448), .A2(new_n600), .A3(new_n607), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n595), .A2(new_n589), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n303), .A2(new_n354), .A3(new_n445), .A4(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n749), .B(new_n565), .C1(new_n569), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n669), .A2(new_n606), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n753), .A2(new_n665), .A3(new_n693), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n752), .A2(new_n697), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n643), .A2(new_n647), .A3(new_n651), .A4(new_n662), .ZN(new_n756));
  INV_X1    g570(.A(new_n701), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n434), .A2(new_n625), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT116), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n611), .A2(new_n303), .A3(new_n722), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n756), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n748), .A2(new_n755), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n647), .A2(new_n651), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n643), .A2(new_n662), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n701), .A4(new_n760), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n674), .A2(new_n699), .A3(new_n665), .A4(new_n693), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n530), .A2(new_n653), .ZN(new_n770));
  OAI22_X1  g584(.A1(new_n769), .A2(KEYINPUT42), .B1(new_n770), .B2(new_n691), .ZN(new_n771));
  INV_X1    g585(.A(new_n754), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n674), .A2(new_n448), .A3(new_n699), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n751), .A2(new_n569), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n608), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n768), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n748), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n765), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n765), .B2(new_n778), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n706), .A2(new_n439), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n657), .A2(new_n650), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n295), .B1(new_n729), .B2(new_n730), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n727), .B(new_n301), .C1(new_n788), .C2(new_n732), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT47), .B1(new_n733), .B2(new_n302), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n728), .A2(KEYINPUT119), .A3(new_n734), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n640), .B(KEYINPUT115), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(KEYINPUT120), .A3(new_n302), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n793), .B2(new_n301), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n657), .A2(new_n722), .A3(new_n785), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n657), .A2(new_n623), .A3(new_n642), .A4(new_n785), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n350), .B1(KEYINPUT121), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  OAI22_X1  g619(.A1(new_n802), .A2(new_n805), .B1(KEYINPUT121), .B2(new_n803), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n653), .A2(new_n669), .A3(new_n785), .A4(new_n642), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n803), .A2(KEYINPUT121), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n623), .A3(new_n808), .A4(new_n804), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n785), .A2(new_n640), .A3(new_n690), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n753), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n641), .B(new_n689), .C1(new_n561), .C2(new_n563), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n439), .A2(new_n620), .A3(new_n704), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n814), .B2(new_n594), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n801), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n589), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n620), .A2(new_n439), .A3(new_n819), .A4(new_n813), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n794), .A2(new_n302), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n800), .B1(new_n735), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n810), .A2(new_n815), .A3(KEYINPUT51), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n818), .A2(new_n436), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n770), .A2(new_n811), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT48), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n784), .A2(KEYINPUT122), .A3(new_n786), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n435), .A2(new_n189), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n763), .A2(new_n764), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n777), .B2(new_n748), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n765), .A2(new_n778), .A3(new_n780), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n827), .A3(new_n786), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n828), .A2(new_n829), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n793), .B(KEYINPUT49), .Z(new_n838));
  NAND2_X1  g652(.A1(new_n623), .A2(new_n653), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n838), .A2(new_n739), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n688), .A3(new_n705), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n837), .A2(new_n841), .ZN(G75));
  AOI21_X1  g656(.A(new_n299), .B1(new_n765), .B2(new_n778), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(G210), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n340), .A2(new_n344), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(new_n342), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT55), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n844), .B2(new_n845), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n189), .A2(G952), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G51));
  NAND2_X1  g666(.A1(new_n765), .A2(new_n778), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n779), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n833), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n685), .A2(KEYINPUT57), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n685), .A2(KEYINPUT57), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n638), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n843), .A2(G469), .A3(new_n713), .A4(new_n714), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(G54));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n863), .B2(new_n393), .ZN(new_n864));
  NAND3_X1  g678(.A1(KEYINPUT123), .A2(KEYINPUT58), .A3(G475), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n843), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n866), .A2(new_n391), .A3(new_n386), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n866), .B1(new_n391), .B2(new_n386), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n867), .A2(new_n868), .A3(new_n851), .ZN(G60));
  NAND2_X1  g683(.A1(new_n855), .A2(new_n585), .ZN(new_n870));
  NAND2_X1  g684(.A1(G478), .A2(G902), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT59), .Z(new_n872));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n851), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n832), .B2(new_n833), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n875), .B2(new_n585), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n873), .A2(new_n876), .ZN(G63));
  NAND2_X1  g691(.A1(G217), .A2(G902), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT60), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n765), .B2(new_n778), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n603), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n881), .B(new_n874), .C1(new_n549), .C2(new_n880), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT61), .B1(new_n881), .B2(KEYINPUT124), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(G66));
  OAI21_X1  g698(.A(G953), .B1(new_n441), .B2(new_n309), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n752), .A2(new_n756), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n846), .B1(G898), .B2(new_n189), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(G69));
  AOI21_X1  g703(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  MUX2_X1   g705(.A(new_n467), .B(new_n457), .S(KEYINPUT30), .Z(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n373), .ZN(new_n893));
  NAND2_X1  g707(.A1(G900), .A2(G953), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n771), .A2(new_n701), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT126), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n719), .A2(new_n653), .A3(new_n530), .A4(new_n661), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT125), .Z(new_n898));
  OAI21_X1  g712(.A(new_n736), .B1(new_n720), .B2(new_n723), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n746), .A2(new_n672), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n896), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n893), .B(new_n894), .C1(new_n902), .C2(G953), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n904));
  INV_X1    g718(.A(new_n893), .ZN(new_n905));
  AND4_X1   g719(.A1(new_n700), .A2(new_n627), .A3(new_n722), .A4(new_n750), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n901), .A2(new_n631), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n901), .A2(KEYINPUT62), .A3(new_n631), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n906), .B(new_n899), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n905), .B1(new_n911), .B2(G953), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n903), .A2(new_n904), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n904), .B1(new_n903), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n891), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n903), .A2(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT127), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n903), .A2(new_n904), .A3(new_n912), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n890), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(G72));
  NAND2_X1  g734(.A1(new_n911), .A2(new_n886), .ZN(new_n921));
  NAND2_X1  g735(.A1(G472), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT63), .Z(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n468), .A2(new_n488), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n476), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n886), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n923), .B1(new_n902), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(new_n488), .A3(new_n477), .A4(new_n468), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n853), .B(new_n923), .C1(new_n617), .C2(new_n515), .ZN(new_n930));
  AND4_X1   g744(.A1(new_n874), .A2(new_n926), .A3(new_n929), .A4(new_n930), .ZN(G57));
endmodule


