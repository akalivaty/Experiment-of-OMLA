//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G131), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G131), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n192), .A2(new_n194), .A3(new_n199), .A4(new_n195), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT78), .A2(G104), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT78), .A2(G104), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(G101), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n202), .B2(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n206), .A3(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT79), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n212), .A2(new_n209), .A3(new_n206), .A4(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n205), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G128), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n218), .B1(new_n222), .B2(new_n216), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n207), .B1(G104), .B2(new_n206), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  AND4_X1   g039(.A1(KEYINPUT10), .A2(new_n215), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(KEYINPUT81), .B(KEYINPUT1), .C1(new_n228), .C2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G128), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT81), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n218), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n215), .A3(new_n225), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT10), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n227), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n204), .A2(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n208), .A2(new_n214), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G101), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n216), .B2(KEYINPUT64), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n230), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(new_n251), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT69), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n245), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n257));
  INV_X1    g071(.A(G101), .ZN(new_n258));
  AOI22_X1  g072(.A1(KEYINPUT3), .A2(new_n207), .B1(new_n211), .B2(new_n213), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n242), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n244), .B1(new_n259), .B2(new_n205), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n243), .A2(G101), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT80), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n256), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n201), .B1(new_n241), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n255), .A2(new_n253), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT80), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT80), .B1(new_n263), .B2(new_n264), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n268), .B(new_n245), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n236), .A2(new_n238), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT82), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n198), .A2(new_n200), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n271), .A2(new_n275), .A3(new_n276), .A4(new_n227), .ZN(new_n277));
  XNOR2_X1  g091(.A(G110), .B(G140), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(G227), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n278), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n267), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n223), .B1(new_n215), .B2(new_n225), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n236), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g100(.A(KEYINPUT83), .B(new_n223), .C1(new_n215), .C2(new_n225), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n201), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT12), .B(new_n201), .C1(new_n286), .C2(new_n287), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n282), .B1(new_n292), .B2(new_n277), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n189), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n267), .A2(new_n277), .A3(new_n282), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n241), .A2(new_n266), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n296), .A2(new_n276), .B1(new_n291), .B2(new_n290), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT84), .B(new_n295), .C1(new_n297), .C2(new_n282), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n294), .A2(G469), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n292), .A2(new_n277), .A3(new_n282), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n282), .B1(new_n267), .B2(new_n277), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n300), .B(new_n301), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n300), .A2(new_n301), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n188), .B1(new_n299), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT85), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n241), .A2(new_n201), .A3(new_n266), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n226), .B1(new_n273), .B2(new_n274), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n276), .B1(new_n312), .B2(new_n271), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n281), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n314), .B2(new_n302), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n306), .B1(new_n315), .B2(new_n300), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n294), .A2(new_n298), .A3(G469), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(new_n188), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G214), .B1(G237), .B2(G902), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n230), .A2(KEYINPUT1), .A3(new_n219), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n222), .A2(new_n216), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n254), .A2(G125), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n324), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n324), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G224), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G953), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n334), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT2), .ZN(new_n342));
  INV_X1    g156(.A(G113), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT2), .A2(G113), .ZN(new_n347));
  XNOR2_X1  g161(.A(G116), .B(G119), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n346), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n345), .ZN(new_n352));
  NOR3_X1   g166(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n348), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT68), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n244), .A2(new_n260), .B1(new_n351), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n269), .B2(new_n270), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n215), .A2(new_n225), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n348), .A2(KEYINPUT5), .ZN(new_n362));
  INV_X1    g176(.A(G116), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n363), .A2(KEYINPUT5), .A3(G119), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n343), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n349), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G122), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n262), .A2(new_n265), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n367), .B1(new_n373), .B2(new_n359), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT87), .A3(new_n369), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n372), .A2(new_n375), .A3(KEYINPUT6), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT86), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n374), .B2(new_n369), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n360), .A2(new_n368), .ZN(new_n382));
  INV_X1    g196(.A(new_n369), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n379), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n339), .B1(new_n376), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n372), .A2(new_n375), .ZN(new_n387));
  INV_X1    g201(.A(new_n333), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n336), .B1(new_n331), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT7), .B1(new_n337), .B2(KEYINPUT89), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(KEYINPUT89), .B2(new_n337), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n332), .A2(new_n333), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n369), .B(KEYINPUT8), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n361), .A2(new_n366), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n367), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT7), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n331), .B2(new_n388), .ZN(new_n397));
  AND4_X1   g211(.A1(new_n389), .A2(new_n392), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(G902), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G210), .B1(G237), .B2(G902), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n386), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n400), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n403));
  AOI211_X1 g217(.A(new_n369), .B(new_n380), .C1(new_n360), .C2(new_n368), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n372), .A2(new_n375), .A3(KEYINPUT6), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n338), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT87), .B1(new_n374), .B2(new_n369), .ZN(new_n408));
  AND4_X1   g222(.A1(KEYINPUT87), .A2(new_n360), .A3(new_n368), .A4(new_n369), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n398), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n301), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n402), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n323), .B1(new_n401), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G952), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n414), .A2(KEYINPUT93), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(KEYINPUT93), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n279), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(G234), .B2(G237), .ZN(new_n418));
  NAND2_X1  g232(.A1(G234), .A2(G237), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(G902), .A3(G953), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT94), .Z(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(G898), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n418), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n424), .B(KEYINPUT95), .Z(new_n425));
  NAND2_X1  g239(.A1(new_n228), .A2(G128), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n219), .A2(G143), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G134), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n427), .A3(new_n191), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT92), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G122), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G116), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n206), .B1(new_n435), .B2(KEYINPUT14), .ZN(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n429), .A2(KEYINPUT92), .A3(new_n430), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT13), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n426), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n427), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n426), .A2(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(G134), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n437), .A2(G107), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n437), .A2(G107), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .A4(new_n430), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G217), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n187), .A2(new_n450), .A3(G953), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n440), .A2(new_n448), .A3(new_n451), .ZN(new_n454));
  AOI21_X1  g268(.A(G902), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n455), .B(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(G104), .Z(new_n462));
  INV_X1    g276(.A(G237), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n279), .A3(G214), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n228), .ZN(new_n465));
  NOR2_X1   g279(.A1(G237), .A2(G953), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(G143), .A3(G214), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT18), .A3(G131), .ZN(new_n469));
  XNOR2_X1  g283(.A(G125), .B(G140), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n220), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT18), .A2(G131), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n464), .A2(new_n228), .ZN(new_n475));
  AOI21_X1  g289(.A(G143), .B1(new_n466), .B2(G214), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT17), .B(G131), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT91), .ZN(new_n478));
  INV_X1    g292(.A(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G125), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n328), .A2(G140), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT16), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(G146), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(G146), .B1(new_n482), .B2(new_n483), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n475), .B2(new_n476), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n489));
  INV_X1    g303(.A(G131), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n465), .A2(new_n490), .A3(new_n467), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n462), .B(new_n474), .C1(new_n478), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n470), .A2(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n498));
  OAI211_X1 g312(.A(new_n497), .B(new_n220), .C1(new_n470), .C2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n484), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n474), .ZN(new_n501));
  INV_X1    g315(.A(new_n462), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(G475), .A2(G902), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n460), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n505), .ZN(new_n507));
  AOI211_X1 g321(.A(KEYINPUT20), .B(new_n507), .C1(new_n494), .C2(new_n503), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n474), .B1(new_n478), .B2(new_n493), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n502), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n510), .B2(new_n494), .ZN(new_n511));
  INV_X1    g325(.A(G475), .ZN(new_n512));
  OAI22_X1  g326(.A1(new_n506), .A2(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n459), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n413), .A2(new_n425), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n517));
  INV_X1    g331(.A(G119), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G128), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(G128), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n517), .B(new_n519), .C1(new_n520), .C2(KEYINPUT23), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G110), .Z(new_n522));
  XNOR2_X1  g336(.A(G119), .B(G128), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n521), .A2(G110), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n470), .A2(new_n220), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n484), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(G110), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n522), .A2(new_n528), .A3(new_n523), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n526), .B1(new_n531), .B2(new_n487), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT22), .B(G137), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n526), .B(new_n535), .C1(new_n531), .C2(new_n487), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n450), .B1(G234), .B2(new_n301), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n301), .A3(new_n538), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n537), .A2(KEYINPUT25), .A3(new_n301), .A4(new_n538), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n545), .A2(KEYINPUT76), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n540), .B1(new_n545), .B2(KEYINPUT76), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT77), .Z(new_n550));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n551));
  NOR2_X1   g365(.A1(G472), .A2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n254), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n192), .A2(new_n194), .A3(new_n490), .A4(new_n195), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n191), .A2(G137), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n193), .A2(G134), .ZN(new_n557));
  OAI21_X1  g371(.A(G131), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n554), .A2(new_n201), .B1(new_n223), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT66), .B1(new_n560), .B2(KEYINPUT30), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n223), .A2(new_n559), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n276), .B2(new_n254), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT66), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n255), .A2(new_n201), .A3(new_n253), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT30), .A3(new_n562), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n351), .A2(new_n358), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n561), .A2(new_n566), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT70), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n349), .A2(new_n350), .A3(new_n340), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT68), .B1(new_n356), .B2(new_n357), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n351), .A2(new_n358), .A3(KEYINPUT70), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n574), .A2(new_n567), .A3(new_n562), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n466), .A2(G210), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT27), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT26), .B(G101), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n570), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT31), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n570), .A2(KEYINPUT31), .A3(new_n576), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT28), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n563), .A2(new_n569), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n576), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n589), .B2(new_n586), .ZN(new_n590));
  INV_X1    g404(.A(new_n580), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n553), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n551), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n583), .A2(new_n584), .B1(new_n590), .B2(new_n591), .ZN(new_n597));
  OAI211_X1 g411(.A(KEYINPUT72), .B(new_n596), .C1(new_n597), .C2(new_n553), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n570), .A2(new_n576), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n591), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT73), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT29), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(KEYINPUT73), .A3(new_n591), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n587), .B(new_n580), .C1(new_n589), .C2(new_n586), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n576), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n574), .A2(new_n575), .B1(new_n567), .B2(new_n562), .ZN(new_n609));
  OAI211_X1 g423(.A(KEYINPUT74), .B(KEYINPUT28), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT74), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n587), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n574), .A2(new_n575), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n567), .A2(new_n562), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n586), .B1(new_n615), .B2(new_n576), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n610), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n591), .A2(new_n604), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n607), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n620), .A2(G472), .B1(KEYINPUT32), .B2(new_n593), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n550), .B1(new_n599), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n321), .A2(new_n516), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  XNOR2_X1  g438(.A(new_n549), .B(KEYINPUT77), .ZN(new_n625));
  INV_X1    g439(.A(new_n593), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n597), .B2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n310), .B2(new_n320), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n401), .A2(new_n412), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n322), .ZN(new_n631));
  INV_X1    g445(.A(new_n425), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n453), .A2(new_n454), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT33), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n453), .A2(new_n635), .A3(new_n454), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n636), .A3(G478), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n456), .A2(new_n301), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n455), .B2(new_n456), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n637), .A2(KEYINPUT96), .A3(new_n639), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n513), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n631), .A2(new_n632), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n629), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NOR2_X1   g466(.A1(new_n511), .A2(new_n512), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n504), .A2(new_n505), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT20), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n504), .A2(new_n460), .A3(new_n505), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT97), .B1(new_n506), .B2(new_n508), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n653), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n458), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n413), .A2(new_n425), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n629), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NAND2_X1  g480(.A1(new_n627), .A2(new_n626), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n536), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n532), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n541), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n547), .B2(new_n548), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n321), .A2(new_n516), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n418), .B1(new_n422), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n660), .A2(new_n459), .A3(new_n671), .A4(new_n679), .ZN(new_n680));
  AOI211_X1 g494(.A(new_n323), .B(new_n680), .C1(new_n412), .C2(new_n401), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n599), .A2(new_n621), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n319), .B1(new_n318), .B2(new_n188), .ZN(new_n683));
  INV_X1    g497(.A(new_n188), .ZN(new_n684));
  AOI211_X1 g498(.A(KEYINPUT85), .B(new_n684), .C1(new_n316), .C2(new_n317), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n681), .B(new_n682), .C1(new_n683), .C2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT98), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n321), .A2(KEYINPUT98), .A3(new_n682), .A4(new_n681), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  INV_X1    g505(.A(KEYINPUT38), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n630), .B(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(G472), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n608), .A2(new_n609), .ZN(new_n695));
  AOI21_X1  g509(.A(G902), .B1(new_n695), .B2(new_n591), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n600), .A2(new_n580), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n593), .B2(KEYINPUT32), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n599), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n672), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n646), .A2(new_n458), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n322), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n693), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n678), .B(KEYINPUT39), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n321), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT99), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT99), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n709), .B(new_n706), .C1(new_n683), .C2(new_n685), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(KEYINPUT40), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT40), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n709), .B1(new_n321), .B2(new_n706), .ZN(new_n713));
  INV_X1    g527(.A(new_n710), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n705), .B1(new_n711), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n228), .ZN(G45));
  AOI22_X1  g531(.A1(new_n310), .A2(new_n320), .B1(new_n599), .B2(new_n621), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n644), .A2(new_n513), .A3(new_n679), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n631), .A2(new_n672), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT100), .B(G146), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G48));
  NOR2_X1   g537(.A1(new_n631), .A2(new_n632), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n314), .A2(new_n302), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n301), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n188), .A3(new_n305), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n622), .A3(new_n647), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n663), .A2(new_n622), .A3(new_n728), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NOR3_X1   g547(.A1(new_n459), .A2(new_n513), .A3(new_n632), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n727), .A2(new_n734), .A3(new_n188), .A4(new_n305), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n599), .B2(new_n621), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n631), .A2(new_n672), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  OAI211_X1 g553(.A(new_n610), .B(new_n591), .C1(new_n612), .C2(new_n616), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n553), .B1(new_n585), .B2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n549), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n627), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT101), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n727), .A2(new_n188), .A3(new_n305), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n631), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n747), .A3(new_n425), .A4(new_n702), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n750));
  INV_X1    g564(.A(new_n719), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT102), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n585), .A2(new_n592), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n301), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n741), .B1(new_n754), .B2(G472), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n752), .B1(new_n755), .B2(new_n671), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n752), .A2(new_n627), .A3(new_n742), .A4(new_n671), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n751), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n728), .A2(new_n413), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n750), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n755), .A2(new_n752), .A3(new_n671), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n627), .A2(new_n742), .A3(new_n671), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT102), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n719), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n747), .A3(KEYINPUT103), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  NAND3_X1  g581(.A1(new_n401), .A2(new_n412), .A3(new_n322), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n401), .A2(new_n412), .A3(KEYINPUT104), .A4(new_n322), .ZN(new_n771));
  INV_X1    g585(.A(new_n293), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(G469), .A3(new_n295), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n684), .B1(new_n316), .B2(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n770), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n622), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n770), .A2(new_n751), .A3(new_n771), .A4(new_n774), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n593), .B2(KEYINPUT32), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT32), .ZN(new_n781));
  OAI211_X1 g595(.A(KEYINPUT106), .B(new_n781), .C1(new_n597), .C2(new_n553), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n593), .A2(KEYINPUT32), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n780), .B(new_n782), .C1(KEYINPUT105), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT105), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n620), .A2(G472), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n743), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT42), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n777), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n490), .ZN(G33));
  NAND4_X1  g605(.A1(new_n622), .A2(new_n770), .A3(new_n771), .A4(new_n774), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n662), .A2(new_n679), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n191), .ZN(G36));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n294), .B2(new_n298), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n772), .A2(KEYINPUT45), .A3(new_n295), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(G469), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n307), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n799), .A2(new_n800), .B1(new_n300), .B2(new_n315), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n800), .B2(new_n799), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n802), .A2(new_n188), .A3(new_n706), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n513), .B1(new_n642), .B2(new_n643), .ZN(new_n804));
  NOR2_X1   g618(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n805));
  AND2_X1   g619(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n804), .B2(new_n806), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n667), .A3(new_n671), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n770), .A2(new_n771), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT108), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n808), .A2(KEYINPUT44), .A3(new_n667), .A4(new_n671), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n814), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n803), .B(new_n811), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  AND2_X1   g633(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n820));
  NOR2_X1   g634(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n802), .B(new_n188), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n812), .A2(new_n682), .A3(new_n625), .A4(new_n719), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n802), .A2(new_n188), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n822), .B(new_n823), .C1(new_n825), .C2(new_n821), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  NAND2_X1  g641(.A1(new_n727), .A2(new_n305), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT49), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n549), .A2(new_n684), .A3(new_n323), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n829), .A2(new_n804), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n700), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n828), .A2(KEYINPUT49), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n693), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n661), .A2(new_n672), .A3(new_n459), .A4(new_n678), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n682), .B(new_n836), .C1(new_n683), .C2(new_n685), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n751), .B(new_n774), .C1(new_n756), .C2(new_n757), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n812), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n790), .A2(new_n794), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n701), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n413), .A2(new_n774), .A3(new_n679), .A4(new_n702), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n718), .A2(new_n720), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n690), .A2(new_n766), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n514), .B1(new_n645), .B2(new_n513), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n425), .A2(new_n630), .A3(new_n322), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n628), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n847), .B(new_n848), .C1(new_n685), .C2(new_n683), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n674), .A2(new_n849), .A3(new_n729), .A4(new_n732), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n623), .A2(new_n748), .A3(new_n738), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n840), .A2(new_n845), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n690), .A2(new_n766), .A3(new_n843), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n835), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n837), .A2(new_n838), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n813), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n792), .A2(new_n793), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n789), .A3(new_n777), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n515), .B1(new_n310), .B2(new_n320), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n682), .A2(new_n625), .A3(new_n728), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n862), .A2(new_n673), .B1(new_n863), .B2(new_n649), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n629), .A2(new_n847), .B1(new_n863), .B2(new_n663), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n702), .A2(new_n425), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n759), .A2(new_n866), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n867), .A2(new_n745), .B1(new_n737), .B2(new_n736), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n864), .A2(new_n865), .A3(new_n623), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(KEYINPUT53), .A3(new_n845), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n857), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT54), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n688), .A2(new_n689), .B1(new_n760), .B2(new_n765), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n844), .B1(new_n876), .B2(new_n843), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n835), .B1(new_n853), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n854), .A2(new_n855), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n870), .A2(KEYINPUT53), .A3(new_n845), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n874), .B1(new_n873), .B2(KEYINPUT54), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n418), .A2(new_n770), .A3(new_n728), .A4(new_n771), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n808), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n788), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT48), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n745), .A2(new_n418), .A3(new_n808), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n417), .B1(new_n890), .B2(new_n747), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n885), .A2(new_n625), .A3(new_n832), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n648), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n746), .A2(new_n322), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n693), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT112), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n693), .A2(KEYINPUT112), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT50), .B1(new_n900), .B2(new_n890), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT50), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n903), .B(new_n889), .C1(new_n898), .C2(new_n899), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n905), .A3(KEYINPUT113), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n644), .A2(new_n513), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n756), .A2(new_n757), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n892), .A2(new_n908), .B1(new_n886), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT113), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n901), .B2(new_n904), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n727), .A2(new_n684), .A3(new_n305), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n820), .A2(new_n821), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n824), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n821), .B1(new_n802), .B2(new_n188), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n889), .A2(new_n812), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n906), .A2(new_n911), .A3(new_n914), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(KEYINPUT114), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT114), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n924), .B(new_n915), .C1(new_n917), .C2(new_n918), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n910), .B1(new_n902), .B2(new_n905), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n912), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n894), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n883), .A2(new_n884), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(G952), .A2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n834), .B1(new_n930), .B2(new_n931), .ZN(G75));
  NOR2_X1   g746(.A1(new_n279), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n301), .B1(new_n878), .B2(new_n881), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(G210), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n376), .A2(new_n385), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n338), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n386), .ZN(new_n939));
  XOR2_X1   g753(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n934), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n936), .A2(new_n941), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT116), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n936), .A2(KEYINPUT116), .A3(new_n941), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(G51));
  INV_X1    g761(.A(new_n882), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n879), .B1(new_n878), .B2(new_n881), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n306), .B(KEYINPUT57), .Z(new_n951));
  OAI21_X1  g765(.A(new_n725), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n796), .A2(new_n798), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT117), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n935), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n933), .B1(new_n952), .B2(new_n955), .ZN(G54));
  AND3_X1   g770(.A1(new_n935), .A2(KEYINPUT58), .A3(G475), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n934), .B1(new_n957), .B2(new_n504), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n504), .B2(new_n957), .ZN(G60));
  NAND2_X1  g773(.A1(new_n634), .A2(new_n636), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n638), .B(KEYINPUT59), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n934), .B1(new_n950), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n883), .B2(new_n884), .ZN(new_n965));
  INV_X1    g779(.A(new_n960), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n878), .B2(new_n881), .ZN(new_n970));
  OR3_X1    g784(.A1(new_n970), .A2(KEYINPUT119), .A3(new_n539), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT119), .B1(new_n970), .B2(new_n539), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n669), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n934), .A2(KEYINPUT61), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT118), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n970), .A2(new_n976), .A3(new_n669), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n934), .B1(new_n970), .B2(new_n539), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n970), .B2(new_n669), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n975), .B1(new_n980), .B2(KEYINPUT61), .ZN(G66));
  NAND2_X1  g795(.A1(new_n869), .A2(new_n279), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT120), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n423), .B2(new_n335), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT121), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n937), .B1(G898), .B2(new_n279), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  NAND3_X1  g802(.A1(new_n561), .A2(new_n566), .A3(new_n568), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n497), .B1(new_n470), .B2(new_n498), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n279), .B1(G227), .B2(G900), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n826), .A2(new_n818), .ZN(new_n996));
  INV_X1    g810(.A(new_n788), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n803), .A2(new_n413), .A3(new_n702), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n860), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n876), .A2(new_n721), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n996), .A2(new_n999), .A3(new_n790), .A4(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1001), .A2(new_n279), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n991), .B1(new_n677), .B2(new_n279), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT62), .B1(new_n716), .B2(new_n1000), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n713), .A2(new_n714), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n846), .B(KEYINPUT123), .Z(new_n1006));
  NAND4_X1  g820(.A1(new_n1005), .A2(new_n622), .A3(new_n813), .A4(new_n1006), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1007), .A2(new_n826), .A3(new_n818), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n711), .A2(new_n715), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n704), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT62), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n876), .A2(new_n721), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT122), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n716), .A2(new_n1000), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT122), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1016), .A2(new_n1017), .A3(new_n1012), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1009), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1019), .A2(G953), .ZN(new_n1020));
  OAI221_X1 g834(.A(new_n995), .B1(new_n1002), .B2(new_n1003), .C1(new_n1020), .C2(new_n991), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1014), .A2(KEYINPUT122), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1017), .B1(new_n1016), .B2(new_n1012), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n991), .B1(new_n1025), .B2(new_n279), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n993), .B(new_n994), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1021), .A2(new_n1028), .ZN(G72));
  XNOR2_X1  g843(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n694), .A2(new_n301), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1030), .B(new_n1031), .Z(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n603), .A2(new_n581), .A3(new_n605), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n873), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1032), .B1(new_n1001), .B2(new_n852), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n570), .A2(new_n576), .A3(new_n591), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n1035), .B(new_n934), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1032), .B1(new_n1019), .B2(new_n852), .ZN(new_n1039));
  OAI21_X1  g853(.A(KEYINPUT126), .B1(new_n1039), .B2(new_n697), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1033), .B1(new_n1025), .B2(new_n869), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT126), .ZN(new_n1042));
  INV_X1    g856(.A(new_n697), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1038), .B1(new_n1040), .B2(new_n1044), .ZN(G57));
endmodule


