//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1248, new_n1249, new_n1250, new_n1251;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G116), .ZN(new_n210));
  INV_X1    g0010(.A(G270), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n213), .A2(new_n214), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n206), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  AND2_X1   g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n226), .B(new_n229), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n216), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n211), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  INV_X1    g0045(.A(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n210), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n208), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G33), .A3(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n256), .A3(new_n230), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT69), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(new_n262), .A3(new_n259), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(G238), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G226), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n230), .A2(new_n253), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT67), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n230), .A2(KEYINPUT67), .A3(new_n253), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n259), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n264), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n264), .A2(new_n276), .A3(new_n282), .A4(new_n279), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G169), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT14), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n281), .A2(G179), .A3(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n284), .A2(new_n289), .A3(G169), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n286), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT72), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n289), .B1(new_n284), .B2(G169), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI211_X1 g0094(.A(KEYINPUT14), .B(new_n294), .C1(new_n281), .C2(new_n283), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT72), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(new_n288), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G1), .A2(G13), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT68), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  INV_X1    g0105(.A(G20), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(G20), .A2(G33), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n305), .B1(new_n307), .B2(new_n208), .C1(new_n309), .C2(new_n202), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT70), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT11), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n311), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n317));
  INV_X1    g0117(.A(G13), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n305), .A2(G1), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(KEYINPUT71), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT12), .ZN(new_n321));
  INV_X1    g0121(.A(new_n301), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n258), .A2(G20), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G68), .A3(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n314), .A2(new_n317), .A3(new_n321), .A4(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n325), .B(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n292), .A2(new_n298), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n258), .B2(G20), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n318), .A2(new_n306), .A3(G1), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n322), .A2(new_n302), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n330), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(new_n331), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n335), .A2(KEYINPUT75), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT75), .B1(new_n335), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n265), .A2(G226), .A3(G1698), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n265), .A2(G223), .A3(new_n266), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G87), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n278), .B1(new_n343), .B2(new_n275), .ZN(new_n344));
  INV_X1    g0144(.A(new_n260), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G232), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(G190), .A3(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(KEYINPUT3), .A2(G33), .ZN(new_n348));
  NAND2_X1  g0148(.A1(KEYINPUT3), .A2(G33), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n306), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n348), .A2(KEYINPUT7), .A3(new_n306), .A4(new_n349), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT74), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT74), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n350), .B2(new_n351), .ZN(new_n356));
  OAI21_X1  g0156(.A(G68), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n215), .A2(new_n304), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n358), .B2(new_n201), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n308), .A2(G159), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT16), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n304), .B1(new_n352), .B2(new_n353), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT16), .ZN(new_n365));
  OR3_X1    g0165(.A1(new_n364), .A2(new_n365), .A3(new_n361), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n301), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n339), .B(new_n347), .C1(new_n363), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT77), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n343), .A2(new_n275), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(new_n279), .A3(new_n346), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G200), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT17), .A4(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n370), .A2(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n370), .A2(KEYINPUT17), .ZN(new_n376));
  INV_X1    g0176(.A(new_n373), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n375), .B(new_n376), .C1(new_n368), .C2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G179), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n344), .A2(new_n379), .A3(new_n346), .ZN(new_n380));
  AOI21_X1  g0180(.A(G169), .B1(new_n344), .B2(new_n346), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT76), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n372), .A2(new_n294), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT76), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n344), .A2(new_n379), .A3(new_n346), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n339), .B1(new_n363), .B2(new_n367), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n387), .A2(KEYINPUT18), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT18), .B1(new_n387), .B2(new_n388), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n374), .B(new_n378), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n265), .A2(G223), .A3(G1698), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n265), .A2(new_n266), .ZN(new_n393));
  INV_X1    g0193(.A(G222), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n392), .B1(new_n208), .B2(new_n265), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n275), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n345), .A2(G226), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n279), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G200), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n396), .A2(G190), .A3(new_n279), .A4(new_n397), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n203), .A2(G20), .ZN(new_n401));
  INV_X1    g0201(.A(G150), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n401), .B1(new_n402), .B2(new_n309), .C1(new_n307), .C2(new_n329), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n303), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n301), .B(KEYINPUT68), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n405), .A2(G50), .A3(new_n323), .A4(new_n332), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n331), .A2(new_n202), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT9), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n404), .A2(new_n406), .A3(KEYINPUT9), .A4(new_n407), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n399), .A2(new_n400), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT10), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n398), .A2(G200), .B1(new_n408), .B2(new_n409), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT10), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(new_n400), .A4(new_n411), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n398), .A2(new_n294), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n408), .B1(new_n398), .B2(G179), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n265), .A2(G1698), .ZN(new_n422));
  INV_X1    g0222(.A(G238), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n421), .B1(new_n246), .B2(new_n265), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n278), .B1(new_n424), .B2(new_n275), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n209), .B2(new_n260), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n294), .ZN(new_n427));
  INV_X1    g0227(.A(new_n329), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n308), .B1(G20), .B2(G77), .ZN(new_n429));
  XOR2_X1   g0229(.A(KEYINPUT15), .B(G87), .Z(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n307), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(new_n301), .B1(new_n208), .B2(new_n331), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n322), .A2(G77), .A3(new_n323), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n427), .B(new_n435), .C1(G179), .C2(new_n426), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n417), .A2(new_n420), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n391), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n325), .B1(G200), .B2(new_n284), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n281), .A2(G190), .A3(new_n283), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n435), .B1(G200), .B2(new_n426), .ZN(new_n442));
  INV_X1    g0242(.A(G190), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(new_n426), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n328), .A2(new_n438), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n258), .A2(G33), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT78), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(new_n322), .A3(G116), .A4(new_n332), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n299), .A2(new_n300), .B1(G20), .B2(new_n210), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(new_n306), .C1(G33), .C2(new_n222), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT20), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n448), .B1(G116), .B2(new_n332), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  INV_X1    g0255(.A(G41), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT5), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(KEYINPUT80), .B2(G41), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G1), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(new_n257), .A3(G270), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n457), .A2(new_n459), .A3(new_n461), .A4(G274), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT3), .A2(G33), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT3), .A2(G33), .ZN(new_n467));
  OAI211_X1 g0267(.A(G257), .B(new_n266), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G264), .B(G1698), .C1(new_n466), .C2(new_n467), .ZN(new_n469));
  INV_X1    g0269(.A(G303), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n468), .B(new_n469), .C1(new_n470), .C2(new_n265), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n275), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n294), .B1(new_n465), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT21), .B1(new_n454), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT85), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n463), .A2(new_n464), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n275), .B2(new_n471), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n473), .A2(KEYINPUT21), .B1(new_n477), .B2(G179), .ZN(new_n478));
  INV_X1    g0278(.A(new_n454), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n465), .A2(new_n472), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(KEYINPUT21), .A3(G169), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n465), .A2(G179), .A3(new_n472), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(KEYINPUT85), .A3(new_n454), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n474), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n454), .B1(new_n481), .B2(G200), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n443), .B2(new_n481), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n306), .B(G87), .C1(new_n466), .C2(new_n467), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT22), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT22), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n265), .A2(new_n492), .A3(new_n306), .A4(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G20), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n306), .A2(G107), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT23), .ZN(new_n499));
  AND4_X1   g0299(.A1(new_n489), .A2(new_n494), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n491), .B2(new_n493), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n489), .B1(new_n501), .B2(new_n499), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n301), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n405), .A2(new_n332), .A3(new_n447), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n331), .A2(new_n246), .ZN(new_n507));
  XOR2_X1   g0307(.A(new_n507), .B(KEYINPUT25), .Z(new_n508));
  NAND3_X1  g0308(.A1(new_n503), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n218), .A2(new_n393), .B1(new_n422), .B2(new_n223), .ZN(new_n510));
  AND2_X1   g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n275), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n462), .A2(new_n257), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G264), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n464), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n294), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n512), .A2(new_n514), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n379), .A3(new_n464), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n503), .A2(new_n506), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n515), .A2(G200), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(G190), .A3(new_n464), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n520), .A2(new_n508), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n486), .A2(new_n488), .A3(new_n519), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n331), .A2(new_n222), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n504), .B2(new_n222), .ZN(new_n526));
  OAI21_X1  g0326(.A(G107), .B1(new_n354), .B2(new_n356), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n246), .A2(KEYINPUT6), .A3(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n222), .A2(new_n246), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n528), .B1(new_n531), .B2(KEYINPUT6), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(G20), .B1(G77), .B2(new_n308), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n526), .B1(new_n534), .B2(new_n301), .ZN(new_n535));
  OAI211_X1 g0335(.A(G250), .B(G1698), .C1(new_n466), .C2(new_n467), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n265), .A2(KEYINPUT79), .A3(G250), .A4(G1698), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n450), .ZN(new_n540));
  OAI211_X1 g0340(.A(G244), .B(new_n266), .C1(new_n466), .C2(new_n467), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n275), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n464), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n513), .B2(G257), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n548), .A3(G190), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT81), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n548), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n546), .A2(new_n548), .A3(KEYINPUT81), .A4(G190), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n535), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n294), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n546), .A2(new_n548), .A3(new_n379), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n322), .B1(new_n527), .B2(new_n533), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n556), .B(new_n557), .C1(new_n558), .C2(new_n526), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n265), .A2(new_n306), .A3(G68), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n306), .B1(new_n269), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n530), .A2(new_n217), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n561), .B1(new_n269), .B2(G20), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n301), .B1(new_n431), .B2(new_n331), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n405), .A2(G87), .A3(new_n332), .A4(new_n447), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(G1698), .C1(new_n466), .C2(new_n467), .ZN(new_n570));
  OAI211_X1 g0370(.A(G238), .B(new_n266), .C1(new_n466), .C2(new_n467), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n495), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n275), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n461), .A2(G274), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n257), .B(G250), .C1(G1), .C2(new_n460), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n573), .A2(G190), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT83), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n572), .A2(new_n275), .B1(G274), .B2(new_n461), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT83), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n578), .A2(new_n579), .A3(G190), .A4(new_n575), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n569), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n505), .A2(new_n430), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(new_n567), .B1(new_n582), .B2(new_n294), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT82), .B1(new_n582), .B2(G179), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT82), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n578), .A2(new_n588), .A3(new_n379), .A4(new_n575), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n555), .A2(new_n559), .A3(new_n584), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT84), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n583), .A2(new_n581), .B1(new_n586), .B2(new_n590), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT84), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n559), .A4(new_n555), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n524), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n445), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g0398(.A(new_n598), .B(KEYINPUT86), .Z(G372));
  INV_X1    g0399(.A(new_n420), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n389), .A2(new_n390), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n297), .B1(new_n296), .B2(new_n288), .ZN(new_n603));
  NOR4_X1   g0403(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT72), .A4(new_n287), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n605), .B2(new_n327), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n374), .A2(new_n378), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n600), .B1(new_n608), .B2(new_n417), .ZN(new_n609));
  INV_X1    g0409(.A(new_n582), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n379), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n586), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n577), .A2(new_n580), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT87), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n583), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n569), .A2(KEYINPUT88), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT88), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n567), .A2(new_n618), .A3(new_n568), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n582), .A2(KEYINPUT87), .A3(G200), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n616), .A2(new_n617), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT89), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n619), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n618), .B1(new_n567), .B2(new_n568), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(KEYINPUT89), .A3(new_n616), .A4(new_n620), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n613), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n555), .A2(new_n559), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n474), .B1(new_n484), .B2(new_n454), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n519), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n628), .A2(new_n629), .A3(new_n523), .A4(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n594), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT26), .B1(new_n633), .B2(new_n559), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n623), .A2(new_n627), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  INV_X1    g0436(.A(new_n559), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .A4(new_n612), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n632), .A2(new_n634), .A3(new_n612), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n445), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n609), .A2(new_n640), .ZN(G369));
  NOR2_X1   g0441(.A1(new_n318), .A2(G20), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n258), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n519), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n509), .A2(new_n648), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n523), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n653), .B2(new_n519), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n486), .A2(new_n648), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT91), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n649), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n630), .A2(new_n454), .A3(new_n648), .ZN(new_n659));
  INV_X1    g0459(.A(new_n648), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n479), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n488), .B(new_n659), .C1(new_n486), .C2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G330), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g0466(.A(new_n666), .B(KEYINPUT92), .Z(G399));
  INV_X1    g0467(.A(new_n227), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n563), .A2(G116), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n233), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n552), .A2(new_n582), .ZN(new_n675));
  INV_X1    g0475(.A(new_n483), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n517), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT93), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n677), .B(new_n679), .Z(new_n680));
  NOR3_X1   g0480(.A1(new_n610), .A2(new_n477), .A3(G179), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n681), .A2(new_n552), .A3(new_n515), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n648), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(KEYINPUT31), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT31), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n597), .B2(new_n660), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n686), .B2(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n639), .A2(new_n660), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n628), .A2(new_n637), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT26), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n486), .A2(new_n519), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n628), .A3(new_n629), .A4(new_n523), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n594), .A2(new_n637), .A3(new_n636), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n693), .A2(new_n612), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .A3(new_n660), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n688), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n674), .B1(new_n701), .B2(G1), .ZN(G364));
  INV_X1    g0502(.A(new_n664), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n258), .B1(new_n642), .B2(G45), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n669), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n662), .A2(new_n663), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n668), .A2(new_n265), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n232), .A2(new_n460), .A3(G50), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n710), .B(new_n711), .C1(new_n251), .C2(new_n460), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(G116), .B2(new_n227), .ZN(new_n713));
  INV_X1    g0513(.A(new_n265), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n668), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n713), .B1(G355), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT95), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G13), .A2(G33), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n300), .B1(G20), .B2(new_n294), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n662), .A2(new_n720), .ZN(new_n724));
  NAND3_X1  g0524(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n443), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n265), .B1(new_n726), .B2(G326), .ZN(new_n727));
  INV_X1    g0527(.A(G311), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n306), .A2(G190), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n379), .A2(G200), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n725), .A2(G190), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(KEYINPUT33), .B(G317), .Z(new_n734));
  OAI221_X1 g0534(.A(new_n727), .B1(new_n728), .B2(new_n731), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n306), .A2(new_n443), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n730), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n729), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(G322), .A2(new_n738), .B1(new_n741), .B2(G329), .ZN(new_n742));
  INV_X1    g0542(.A(G283), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n379), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n729), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n736), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n742), .B1(new_n743), .B2(new_n745), .C1(new_n470), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n739), .A2(G190), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n735), .B(new_n747), .C1(G294), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT32), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n741), .B2(G159), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(G68), .B2(new_n732), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n749), .A2(G97), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n726), .A2(G50), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n741), .A2(new_n751), .A3(G159), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n746), .A2(new_n217), .ZN(new_n758));
  INV_X1    g0558(.A(new_n745), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G107), .A2(new_n759), .B1(new_n738), .B2(G58), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n208), .B2(new_n731), .ZN(new_n761));
  NOR4_X1   g0561(.A1(new_n757), .A2(new_n714), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n721), .B1(new_n750), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n723), .A2(new_n724), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n706), .B(KEYINPUT94), .Z(new_n765));
  OAI21_X1  g0565(.A(new_n709), .B1(new_n764), .B2(new_n765), .ZN(G396));
  NAND2_X1  g0566(.A1(new_n435), .A2(new_n648), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n444), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n436), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n436), .A2(new_n648), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n689), .B(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(new_n688), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n707), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n714), .B1(new_n741), .B2(G132), .ZN(new_n775));
  INV_X1    g0575(.A(new_n749), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n775), .B1(new_n202), .B2(new_n746), .C1(new_n215), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n731), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G159), .B1(G137), .B2(new_n726), .ZN(new_n779));
  INV_X1    g0579(.A(G143), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n779), .B1(new_n780), .B2(new_n737), .C1(new_n402), .C2(new_n733), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT34), .Z(new_n782));
  AOI211_X1 g0582(.A(new_n777), .B(new_n782), .C1(G68), .C2(new_n759), .ZN(new_n783));
  INV_X1    g0583(.A(new_n746), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G107), .A2(new_n784), .B1(new_n778), .B2(G116), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n728), .B2(new_n740), .ZN(new_n786));
  INV_X1    g0586(.A(new_n726), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n754), .B1(new_n787), .B2(new_n470), .C1(new_n743), .C2(new_n733), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n745), .A2(new_n217), .ZN(new_n789));
  INV_X1    g0589(.A(G294), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n714), .B1(new_n737), .B2(new_n790), .ZN(new_n791));
  NOR4_X1   g0591(.A1(new_n786), .A2(new_n788), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n721), .B1(new_n783), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n765), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n721), .A2(new_n718), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(G77), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n793), .B(new_n798), .C1(new_n771), .C2(new_n719), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n774), .A2(new_n799), .ZN(G384));
  NAND2_X1  g0600(.A1(new_n593), .A2(new_n596), .ZN(new_n801));
  AND3_X1   g0601(.A1(new_n486), .A2(new_n519), .A3(new_n523), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n801), .A2(new_n802), .A3(new_n488), .A4(new_n660), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n803), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n683), .A2(KEYINPUT31), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(new_n805), .A3(new_n771), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n327), .A2(new_n648), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n328), .A2(new_n441), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n328), .B2(new_n441), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n646), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n365), .B1(new_n364), .B2(new_n361), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n366), .A2(new_n303), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT98), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n339), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n339), .A2(new_n814), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT98), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n391), .A2(new_n812), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n369), .A2(new_n373), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT37), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n387), .A2(new_n388), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n388), .A2(new_n812), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n387), .A2(new_n818), .A3(new_n816), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n818), .A2(new_n812), .A3(new_n816), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n820), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n827), .B2(new_n821), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n819), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT99), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n819), .A2(new_n828), .A3(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n819), .A2(new_n828), .A3(KEYINPUT99), .A4(KEYINPUT38), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n811), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n824), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT100), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n839), .A2(KEYINPUT100), .A3(new_n824), .ZN(new_n843));
  INV_X1    g0643(.A(new_n391), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n823), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n830), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n832), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(KEYINPUT40), .A3(new_n811), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n837), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n687), .A2(new_n445), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(G330), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT39), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n833), .B2(new_n834), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT39), .B1(new_n846), .B2(new_n832), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n328), .A2(new_n648), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n601), .A2(new_n812), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n639), .A2(new_n771), .A3(new_n660), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n770), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n810), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n834), .A3(new_n833), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n860), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n691), .A2(new_n445), .A3(new_n698), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n609), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n867), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n854), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n258), .B2(new_n642), .ZN(new_n872));
  OAI211_X1 g0672(.A(G20), .B(new_n230), .C1(new_n532), .C2(KEYINPUT35), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n210), .B(new_n873), .C1(KEYINPUT35), .C2(new_n532), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT97), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT36), .Z(new_n876));
  OAI21_X1  g0676(.A(G77), .B1(new_n215), .B2(new_n304), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n233), .A2(new_n877), .B1(G50), .B2(new_n304), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(G1), .A3(new_n318), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n872), .A2(new_n876), .A3(new_n879), .ZN(G367));
  OAI21_X1  g0680(.A(new_n629), .B1(new_n535), .B2(new_n660), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n559), .B2(new_n660), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n657), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT42), .Z(new_n885));
  INV_X1    g0685(.A(KEYINPUT105), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n883), .B(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n519), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n637), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n885), .B1(new_n889), .B2(new_n648), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n648), .B1(new_n624), .B2(new_n625), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n628), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n612), .B2(new_n891), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(KEYINPUT43), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(KEYINPUT43), .B2(new_n893), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(KEYINPUT106), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  INV_X1    g0698(.A(new_n665), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n887), .A2(new_n899), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n900), .B1(new_n897), .B2(new_n898), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n669), .B(KEYINPUT41), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n658), .A2(new_n883), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT44), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n658), .A2(new_n883), .ZN(new_n907));
  XOR2_X1   g0707(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n908));
  XNOR2_X1  g0708(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n899), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n899), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n664), .A2(KEYINPUT108), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n664), .B(KEYINPUT108), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n654), .A2(new_n656), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n657), .A2(new_n916), .ZN(new_n917));
  MUX2_X1   g0717(.A(new_n914), .B(new_n915), .S(new_n917), .Z(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n700), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n912), .A2(new_n913), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n904), .B1(new_n920), .B2(new_n701), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n901), .B(new_n902), .C1(new_n705), .C2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n710), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n722), .B1(new_n227), .B2(new_n431), .C1(new_n242), .C2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n784), .A2(KEYINPUT46), .A3(G116), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT46), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n746), .B2(new_n210), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n925), .B(new_n927), .C1(new_n246), .C2(new_n776), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(G311), .B2(new_n726), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n714), .B1(new_n733), .B2(new_n790), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n745), .A2(new_n222), .B1(new_n731), .B2(new_n743), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n930), .B(new_n931), .C1(G317), .C2(new_n741), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n929), .B(new_n932), .C1(new_n470), .C2(new_n737), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n745), .A2(new_n208), .ZN(new_n934));
  INV_X1    g0734(.A(G137), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n737), .A2(new_n402), .B1(new_n740), .B2(new_n935), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n934), .B(new_n936), .C1(G50), .C2(new_n778), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n749), .A2(G68), .ZN(new_n938));
  INV_X1    g0738(.A(G159), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n733), .A2(new_n939), .B1(new_n787), .B2(new_n780), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G58), .B2(new_n784), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n937), .A2(new_n265), .A3(new_n938), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT47), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n765), .B1(new_n944), .B2(new_n721), .ZN(new_n945));
  INV_X1    g0745(.A(new_n720), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n924), .B(new_n945), .C1(new_n893), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n922), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(KEYINPUT109), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT109), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n922), .B2(new_n947), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n949), .A2(new_n951), .ZN(G387));
  INV_X1    g0752(.A(new_n919), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n670), .B1(new_n918), .B2(new_n700), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n239), .A2(new_n460), .ZN(new_n956));
  INV_X1    g0756(.A(new_n671), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n956), .A2(new_n710), .B1(new_n957), .B2(new_n715), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n329), .A2(G50), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT50), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n671), .B1(new_n304), .B2(new_n208), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  AOI211_X1 g0761(.A(G45), .B(new_n961), .C1(new_n960), .C2(new_n959), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n958), .A2(new_n962), .B1(G107), .B2(new_n227), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n765), .B1(new_n963), .B2(new_n722), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n778), .A2(G303), .B1(G322), .B2(new_n726), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n728), .B2(new_n733), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G317), .B2(new_n738), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT48), .Z(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n743), .B2(new_n776), .C1(new_n790), .C2(new_n746), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT49), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n741), .A2(G326), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n970), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n265), .B1(new_n759), .B2(G116), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n776), .A2(new_n431), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n428), .B2(new_n732), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n939), .B2(new_n787), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n746), .A2(new_n208), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G150), .B2(new_n741), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n202), .B2(new_n737), .C1(new_n304), .C2(new_n731), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n745), .A2(new_n222), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n978), .A2(new_n981), .A3(new_n714), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT110), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n975), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT111), .ZN(new_n986));
  INV_X1    g0786(.A(new_n721), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n964), .B1(new_n654), .B2(new_n946), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n955), .B(new_n988), .C1(new_n704), .C2(new_n918), .ZN(G393));
  INV_X1    g0789(.A(new_n913), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n953), .B1(new_n990), .B2(new_n911), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n920), .A3(new_n669), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n746), .A2(new_n304), .B1(new_n740), .B2(new_n780), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n776), .A2(new_n208), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n428), .C2(new_n778), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n714), .B(new_n789), .C1(G50), .C2(new_n732), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n787), .A2(new_n402), .B1(new_n737), .B2(new_n939), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT51), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n738), .A2(G311), .B1(G317), .B2(new_n726), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT52), .Z(new_n1001));
  AOI22_X1  g0801(.A1(new_n784), .A2(G283), .B1(new_n741), .B2(G322), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n733), .A2(new_n470), .B1(new_n745), .B2(new_n246), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n265), .B(new_n1003), .C1(G116), .C2(new_n749), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n731), .A2(new_n790), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n999), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n765), .B1(new_n1007), .B2(new_n721), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n887), .B2(new_n946), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n248), .A2(new_n710), .B1(G97), .B2(new_n668), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(new_n722), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n990), .A2(new_n911), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n705), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT112), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n992), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1014), .B1(new_n992), .B2(new_n1013), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(G390));
  NAND4_X1  g0818(.A1(new_n445), .A2(G330), .A3(new_n804), .A4(new_n805), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n609), .A2(new_n868), .A3(new_n1019), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n806), .A2(new_n810), .A3(new_n663), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n804), .A2(new_n805), .A3(G330), .A4(new_n771), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1022), .A2(new_n810), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n863), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n441), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n327), .B(new_n648), .C1(new_n605), .C2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n328), .A2(new_n441), .A3(new_n807), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n687), .A2(G330), .A3(new_n771), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1022), .A2(new_n810), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n697), .A2(new_n660), .A3(new_n769), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n770), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1020), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n856), .A2(new_n857), .B1(new_n865), .B2(new_n859), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n859), .B(KEYINPUT113), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n847), .B(new_n1037), .C1(new_n810), .C2(new_n1033), .ZN(new_n1038));
  AOI211_X1 g0838(.A(KEYINPUT114), .B(new_n1021), .C1(new_n1036), .C2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1029), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1021), .A2(KEYINPUT114), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1036), .A2(new_n1041), .A3(new_n1042), .A4(new_n1038), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1035), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n1040), .A3(new_n1029), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n609), .A2(new_n868), .A3(new_n1019), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n864), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1047), .A2(new_n1051), .A3(new_n1043), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1045), .A2(new_n669), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n726), .A2(G128), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n733), .B2(new_n935), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n265), .B1(new_n776), .B2(new_n939), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G50), .C2(new_n759), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n746), .A2(new_n402), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1059));
  XNOR2_X1  g0859(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(KEYINPUT54), .B(G143), .Z(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(G125), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1062), .A2(new_n731), .B1(new_n1063), .B2(new_n740), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(G132), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1057), .B(new_n1065), .C1(new_n1066), .C2(new_n737), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n745), .A2(new_n304), .B1(new_n737), .B2(new_n210), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1068), .B(new_n994), .C1(G294), .C2(new_n741), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n265), .B(new_n758), .C1(G283), .C2(new_n726), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n778), .A2(G97), .B1(G107), .B2(new_n732), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT117), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n765), .B1(new_n1074), .B2(new_n721), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n428), .B2(new_n796), .C1(new_n858), .C2(new_n719), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT115), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1047), .A2(new_n1043), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n705), .ZN(new_n1079));
  AOI211_X1 g0879(.A(KEYINPUT115), .B(new_n704), .C1(new_n1047), .C2(new_n1043), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1053), .B(new_n1076), .C1(new_n1079), .C2(new_n1080), .ZN(G378));
  INV_X1    g0881(.A(KEYINPUT57), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n837), .A2(G330), .A3(new_n848), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n408), .A2(new_n812), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n417), .A2(new_n420), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n417), .B2(new_n420), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT55), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT56), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1085), .A2(new_n1086), .A3(KEYINPUT55), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1083), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT119), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1093), .A2(KEYINPUT119), .A3(new_n1094), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1100), .A2(G330), .A3(new_n837), .A4(new_n848), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n867), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n860), .A2(new_n861), .A3(new_n866), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n1101), .A3(new_n1096), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1024), .A2(new_n1034), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1020), .B1(new_n1078), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1082), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(KEYINPUT57), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n669), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n719), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n796), .A2(G50), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n733), .A2(new_n1066), .B1(new_n787), .B2(new_n1063), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G128), .A2(new_n738), .B1(new_n778), .B2(G137), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n746), .B2(new_n1062), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(G150), .C2(new_n749), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT59), .ZN(new_n1120));
  AOI21_X1  g0920(.A(G41), .B1(new_n741), .B2(G124), .ZN(new_n1121));
  AOI21_X1  g0921(.A(G33), .B1(new_n759), .B2(G159), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n938), .B1(new_n787), .B2(new_n210), .C1(new_n222), .C2(new_n733), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n1124), .A2(G41), .A3(new_n265), .A4(new_n979), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n737), .A2(new_n246), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n745), .A2(new_n215), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n430), .C2(new_n778), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1125), .B(new_n1128), .C1(new_n743), .C2(new_n740), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT58), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n202), .B1(new_n466), .B2(G41), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1123), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT118), .Z(new_n1133));
  OAI21_X1  g0933(.A(new_n706), .B1(new_n1133), .B2(new_n987), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1114), .A2(new_n1115), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n1111), .B2(new_n705), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1113), .A2(new_n1136), .ZN(G375));
  NAND2_X1  g0937(.A1(new_n1107), .A2(new_n705), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G137), .A2(new_n738), .B1(new_n741), .B2(G128), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n402), .B2(new_n731), .C1(new_n939), .C2(new_n746), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n749), .A2(G50), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1061), .A2(new_n732), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n726), .A2(G132), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n265), .A4(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1140), .A2(new_n1127), .A3(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G97), .A2(new_n784), .B1(new_n738), .B2(G283), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n246), .B2(new_n731), .C1(new_n470), .C2(new_n740), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n733), .A2(new_n210), .B1(new_n787), .B2(new_n790), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1147), .A2(new_n934), .A3(new_n976), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1145), .B1(new_n1149), .B2(new_n714), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n794), .B1(G68), .B2(new_n796), .C1(new_n1150), .C2(new_n987), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT120), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1028), .B2(new_n719), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1138), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1024), .A2(new_n1020), .A3(new_n1034), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1051), .A2(new_n903), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(G381));
  NOR4_X1   g0958(.A1(G387), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1159));
  INV_X1    g0959(.A(G384), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(G375), .A2(G378), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(G407));
  INV_X1    g0963(.A(G213), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1164), .A2(G343), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT121), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(G407), .A2(G213), .A3(new_n1167), .ZN(G409));
  INV_X1    g0968(.A(new_n1165), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1076), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1053), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1110), .A2(new_n903), .A3(new_n1111), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1136), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1136), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n670), .B1(new_n1176), .B2(new_n1082), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1177), .B2(new_n1112), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1169), .B(new_n1174), .C1(new_n1178), .C2(new_n1172), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1165), .A2(G2897), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT122), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1049), .A2(new_n1050), .A3(new_n1048), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n669), .B1(new_n1182), .B2(KEYINPUT60), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT60), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1051), .B2(new_n1156), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1181), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT60), .B1(new_n1182), .B2(new_n1035), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n670), .B1(new_n1156), .B2(new_n1184), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(KEYINPUT122), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G384), .B1(new_n1190), .B2(new_n1155), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1160), .B(new_n1154), .C1(new_n1186), .C2(new_n1189), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT123), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1183), .A2(new_n1185), .A3(new_n1181), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT122), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1155), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1160), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(G384), .A3(new_n1155), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT123), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1180), .B1(new_n1194), .B2(new_n1200), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1191), .A2(new_n1192), .A3(new_n1180), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT124), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1180), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1193), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1198), .A2(KEYINPUT123), .A3(new_n1199), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT124), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1208), .A2(new_n1209), .A3(new_n1202), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1179), .B1(new_n1204), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT126), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT61), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1172), .B1(new_n1113), .B2(new_n1136), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1173), .A2(new_n1136), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1216), .A2(G378), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1215), .A2(new_n1165), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1201), .A2(KEYINPUT124), .A3(new_n1203), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1209), .B1(new_n1208), .B2(new_n1202), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT126), .B1(new_n1221), .B2(KEYINPUT61), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1194), .A2(new_n1200), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1225));
  NOR3_X1   g1025(.A1(new_n1179), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT62), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(KEYINPUT127), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1226), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1214), .A2(new_n1222), .A3(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n948), .A2(new_n1161), .ZN(new_n1232));
  XOR2_X1   g1032(.A(G393), .B(G396), .Z(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n949), .A2(new_n951), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(G390), .B(KEYINPUT125), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n948), .A2(new_n1161), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1233), .B1(new_n1238), .B2(new_n1232), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1231), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT63), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1227), .B1(new_n1221), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1218), .A2(KEYINPUT63), .A3(new_n1223), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1213), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1246), .ZN(G405));
  NOR2_X1   g1047(.A1(new_n1162), .A2(new_n1215), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1224), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1248), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1242), .B(new_n1251), .ZN(G402));
endmodule


