//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  NOR2_X1   g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n188), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(new_n194), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n187), .B1(new_n197), .B2(new_n194), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(new_n195), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT66), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT64), .A2(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G137), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n207), .A2(G137), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n205), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT64), .B(G134), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT11), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT64), .A2(G134), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT64), .A2(G134), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n205), .B1(new_n221), .B2(G137), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n211), .B1(new_n221), .B2(G137), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n218), .B(new_n222), .C1(new_n223), .C2(new_n205), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(G143), .B2(new_n189), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n191), .A2(G146), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n189), .A2(G143), .ZN(new_n230));
  OAI22_X1  g044(.A1(new_n227), .A2(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n190), .A2(new_n192), .A3(new_n226), .A4(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(G137), .B1(new_n208), .B2(new_n209), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT65), .B1(new_n215), .B2(G134), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n207), .A3(G137), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n204), .A2(new_n225), .B1(new_n224), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT2), .B(G113), .Z(new_n242));
  XNOR2_X1  g056(.A(G116), .B(G119), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT28), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n248));
  NOR2_X1   g062(.A1(G237), .A2(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n248), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n240), .A2(new_n224), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n219), .A2(new_n220), .A3(new_n215), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT11), .B1(new_n256), .B2(new_n211), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n218), .B1(new_n257), .B2(new_n222), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n213), .A2(new_n216), .A3(G131), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n199), .B1(new_n196), .B2(new_n198), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT66), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n245), .B(new_n255), .C1(new_n260), .C2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n196), .A2(new_n198), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n217), .B2(new_n224), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n233), .A2(new_n239), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n244), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n247), .B(new_n254), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n204), .A2(new_n225), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT30), .A3(new_n255), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n266), .B2(new_n268), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n244), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n264), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n253), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n254), .A2(KEYINPUT29), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n241), .A2(KEYINPUT70), .A3(new_n245), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n264), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n274), .A2(new_n255), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT71), .B1(new_n289), .B2(new_n244), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n241), .A2(new_n291), .A3(new_n245), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n286), .B(new_n288), .C1(new_n290), .C2(new_n292), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n246), .B(new_n285), .C1(new_n293), .C2(KEYINPUT28), .ZN(new_n294));
  OAI21_X1  g108(.A(G472), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n272), .B1(new_n264), .B2(new_n269), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n253), .B1(new_n296), .B2(new_n246), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT31), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n278), .A2(new_n300), .A3(new_n264), .A4(new_n254), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n278), .A2(new_n264), .A3(new_n254), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT31), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT69), .B(new_n253), .C1(new_n296), .C2(new_n246), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n299), .A2(new_n301), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT32), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n295), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT22), .B(G137), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(G221), .A3(G234), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT77), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(G128), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n228), .A2(KEYINPUT73), .A3(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT24), .B(G110), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n317), .B2(G128), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n228), .A2(KEYINPUT23), .A3(G119), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n319), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n323), .B1(G110), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G125), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT74), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n331), .A2(G140), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n336), .A3(KEYINPUT16), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n189), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n189), .B1(new_n337), .B2(new_n339), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI211_X1 g157(.A(KEYINPUT75), .B(new_n189), .C1(new_n337), .C2(new_n339), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n328), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n327), .ZN(new_n346));
  INV_X1    g160(.A(G110), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n346), .A2(new_n347), .B1(new_n321), .B2(new_n322), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n329), .A2(G125), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT76), .B1(new_n334), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n330), .A2(new_n332), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n189), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n341), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n315), .B1(new_n345), .B2(new_n356), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n331), .A2(KEYINPUT74), .A3(G140), .ZN(new_n358));
  XNOR2_X1  g172(.A(G125), .B(G140), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(KEYINPUT74), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n338), .B1(new_n360), .B2(KEYINPUT16), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT75), .B1(new_n361), .B2(new_n189), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n341), .A2(new_n342), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n340), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n355), .B1(new_n364), .B2(new_n328), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n357), .A2(KEYINPUT78), .B1(new_n365), .B2(new_n314), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n365), .B2(new_n315), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT72), .B(G217), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(G234), .B2(new_n283), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G902), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT79), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT80), .ZN(new_n374));
  INV_X1    g188(.A(new_n370), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n345), .A2(new_n356), .ZN(new_n376));
  INV_X1    g190(.A(new_n315), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(KEYINPUT78), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n365), .A2(new_n314), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n368), .A2(new_n283), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n366), .A2(KEYINPUT25), .A3(new_n283), .A4(new_n368), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G469), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(G104), .ZN(new_n390));
  INV_X1    g204(.A(G104), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT81), .A3(G107), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G101), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n388), .A2(G104), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G101), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n388), .A2(KEYINPUT3), .A3(G104), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT3), .B1(new_n388), .B2(G104), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n396), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n232), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n402), .A2(G128), .B1(new_n190), .B2(new_n192), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n394), .B(new_n400), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT10), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n391), .B2(G107), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n388), .A2(KEYINPUT3), .A3(G104), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n395), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n407), .B1(new_n411), .B2(new_n397), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n407), .A3(G101), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n406), .B1(new_n417), .B2(new_n204), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n404), .A2(new_n405), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n404), .A2(KEYINPUT82), .A3(new_n405), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n423), .A3(new_n260), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n394), .A2(new_n400), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n401), .A2(new_n403), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n404), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n225), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT12), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(KEYINPUT12), .A3(new_n225), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G140), .ZN(new_n434));
  INV_X1    g248(.A(G227), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(G953), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n434), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n424), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n404), .A2(new_n405), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n415), .A2(new_n261), .A3(new_n262), .A4(new_n416), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n404), .A2(KEYINPUT82), .A3(new_n405), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT82), .B1(new_n404), .B2(new_n405), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n440), .B(new_n441), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n225), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n438), .B1(new_n445), .B2(new_n424), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n386), .B(new_n283), .C1(new_n439), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(G469), .A2(G902), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n424), .A2(new_n433), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n437), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n445), .A2(new_n424), .A3(new_n438), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(G469), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G214), .B1(G237), .B2(G902), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G210), .B1(G237), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n233), .A2(new_n331), .ZN(new_n458));
  OAI21_X1  g272(.A(G125), .B1(new_n196), .B2(new_n198), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n312), .A2(G224), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT6), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n415), .A2(new_n244), .A3(new_n416), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n317), .A2(G116), .ZN(new_n468));
  INV_X1    g282(.A(G116), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G119), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT5), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n469), .A2(KEYINPUT5), .A3(G119), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(G113), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n242), .A2(new_n243), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n425), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G122), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n467), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n467), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n466), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n467), .A2(new_n476), .ZN(new_n481));
  INV_X1    g295(.A(new_n477), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n465), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n463), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n461), .A2(KEYINPUT7), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n458), .A2(new_n459), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n460), .A2(KEYINPUT7), .A3(new_n461), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n477), .B(KEYINPUT8), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n425), .A2(new_n475), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n400), .A2(new_n394), .B1(new_n473), .B2(new_n474), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT84), .A4(new_n486), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n489), .A2(new_n490), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n283), .B1(new_n496), .B2(new_n478), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n457), .B1(new_n485), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n467), .A2(new_n476), .A3(new_n477), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n465), .B1(new_n483), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n479), .A2(new_n466), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n462), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND4_X1   g316(.A1(new_n489), .A2(new_n490), .A3(new_n494), .A4(new_n495), .ZN(new_n503));
  AOI21_X1  g317(.A(G902), .B1(new_n503), .B2(new_n499), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n456), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n455), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT9), .B(G234), .ZN(new_n507));
  OAI21_X1  g321(.A(G221), .B1(new_n507), .B2(G902), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n453), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G237), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n312), .A3(G214), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n191), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n249), .A2(G143), .A3(G214), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G131), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT17), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n514), .B(new_n218), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(KEYINPUT17), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n518), .A2(new_n363), .A3(new_n340), .A4(new_n362), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n333), .A2(new_n336), .A3(G146), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n353), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT18), .A2(G131), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AND4_X1   g337(.A1(G143), .A2(new_n510), .A3(new_n312), .A4(G214), .ZN(new_n524));
  AOI21_X1  g338(.A(G143), .B1(new_n249), .B2(G214), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n512), .A2(new_n527), .A3(new_n513), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n522), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n521), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT86), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n526), .A2(new_n527), .A3(new_n523), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n522), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT86), .A3(new_n521), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n519), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G113), .B(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n391), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n519), .A2(new_n541), .A3(new_n538), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n283), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G475), .ZN(new_n547));
  INV_X1    g361(.A(G122), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G116), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n469), .A2(G122), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n388), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n191), .A2(G128), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n228), .A2(G143), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n553), .A2(new_n554), .ZN(new_n558));
  OAI21_X1  g372(.A(G134), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n221), .A2(new_n553), .A3(new_n556), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n553), .A2(new_n556), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n214), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n551), .A2(new_n388), .ZN(new_n565));
  OR3_X1    g379(.A1(new_n548), .A2(KEYINPUT14), .A3(G116), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n566), .A2(new_n549), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n564), .B(new_n565), .C1(new_n388), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  OR3_X1    g384(.A1(new_n369), .A2(new_n507), .A3(G953), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n283), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n312), .A2(G952), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(G234), .B2(G237), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n283), .B(new_n312), .C1(G234), .C2(G237), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT21), .B(G898), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n572), .B(new_n283), .C1(KEYINPUT15), .C2(new_n574), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n576), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n360), .A2(KEYINPUT19), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n350), .A2(new_n352), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n585), .B(new_n189), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n526), .A2(new_n218), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n341), .B1(new_n515), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n533), .A2(new_n537), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT88), .B1(new_n591), .B2(new_n541), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n588), .ZN(new_n593));
  INV_X1    g407(.A(new_n537), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT86), .B1(new_n536), .B2(new_n521), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT88), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n542), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n598), .A3(new_n544), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT20), .ZN(new_n600));
  NOR2_X1   g414(.A1(G475), .A2(G902), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n600), .B1(new_n599), .B2(new_n601), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n547), .B(new_n584), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n509), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n310), .A2(new_n385), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(new_n305), .A2(new_n283), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n608), .A2(G472), .B1(new_n307), .B2(new_n305), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n453), .A2(new_n508), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n385), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G475), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n545), .B2(new_n283), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n599), .A2(new_n601), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT20), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n485), .A2(new_n457), .A3(new_n497), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n456), .B1(new_n502), .B2(new_n504), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n454), .B(new_n582), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n573), .A2(new_n574), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n572), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n570), .A2(KEYINPUT89), .A3(new_n571), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n571), .A2(KEYINPUT89), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n561), .A2(new_n569), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(KEYINPUT33), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT90), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n626), .A2(KEYINPUT90), .A3(KEYINPUT33), .A4(new_n628), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n625), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n574), .A2(G902), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n623), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n619), .A2(new_n622), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n613), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n506), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT91), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n617), .A2(new_n643), .A3(new_n618), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n615), .B1(new_n576), .B2(new_n583), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n603), .A2(KEYINPUT91), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n644), .A2(new_n645), .A3(new_n582), .A4(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n642), .B1(new_n648), .B2(KEYINPUT92), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT92), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n613), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n382), .A2(new_n383), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n370), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n377), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n376), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n372), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n605), .A2(new_n609), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT93), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n578), .B1(new_n579), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AND4_X1   g481(.A1(new_n646), .A2(new_n644), .A3(new_n645), .A4(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n509), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n310), .A2(new_n668), .A3(new_n669), .A4(new_n660), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  INV_X1    g485(.A(KEYINPUT96), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n666), .B(KEYINPUT39), .Z(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT40), .B1(new_n610), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n610), .A2(KEYINPUT40), .A3(new_n674), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(KEYINPUT96), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n498), .A2(new_n505), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n547), .B1(new_n602), .B2(new_n603), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n576), .A2(new_n583), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n683), .A2(new_n686), .A3(new_n455), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n305), .A2(new_n307), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT32), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n293), .A2(new_n253), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT95), .B1(new_n692), .B2(new_n302), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(KEYINPUT95), .A3(new_n302), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n283), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n660), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n678), .A2(new_n680), .A3(new_n687), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NOR3_X1   g513(.A1(new_n619), .A2(new_n637), .A3(new_n666), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n310), .A2(new_n669), .A3(new_n700), .A4(new_n660), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NAND3_X1  g516(.A1(new_n424), .A2(new_n433), .A3(new_n438), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n445), .A2(new_n424), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n703), .B1(new_n704), .B2(new_n438), .ZN(new_n705));
  NAND2_X1  g519(.A1(KEYINPUT97), .A2(G469), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n283), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n283), .B1(new_n439), .B2(new_n446), .ZN(new_n708));
  INV_X1    g522(.A(new_n706), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n707), .A2(new_n710), .A3(new_n508), .ZN(new_n711));
  AND4_X1   g525(.A1(new_n310), .A2(new_n385), .A3(new_n638), .A4(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT41), .B(G113), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  OR2_X1    g528(.A1(new_n374), .A2(new_n384), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n691), .B2(new_n295), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n649), .A2(new_n716), .A3(new_n651), .A4(new_n711), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  INV_X1    g532(.A(new_n604), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n660), .A3(new_n711), .A4(new_n506), .ZN(new_n720));
  INV_X1    g534(.A(G472), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n296), .A2(new_n246), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT29), .B1(new_n722), .B2(new_n254), .ZN(new_n723));
  AOI21_X1  g537(.A(G902), .B1(new_n723), .B2(new_n280), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n293), .A2(KEYINPUT28), .ZN(new_n725));
  INV_X1    g539(.A(new_n285), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n247), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n721), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n689), .B2(new_n690), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT98), .B1(new_n720), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n506), .A2(new_n508), .A3(new_n707), .A4(new_n710), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n604), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT98), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n310), .A2(new_n732), .A3(new_n733), .A4(new_n660), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT99), .B(G119), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G21));
  INV_X1    g551(.A(new_n622), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n711), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT101), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n686), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n684), .A2(KEYINPUT101), .A3(new_n685), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n246), .B1(new_n293), .B2(KEYINPUT28), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n303), .B1(new_n744), .B2(new_n254), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT100), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(KEYINPUT100), .B(new_n303), .C1(new_n744), .C2(new_n254), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n301), .A3(new_n748), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n749), .A2(new_n307), .B1(G472), .B2(new_n608), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n743), .A2(new_n750), .A3(new_n385), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n307), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n608), .A2(G472), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n684), .A2(new_n636), .A3(new_n667), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n731), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n753), .A2(new_n754), .A3(new_n756), .A4(new_n660), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT103), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n310), .A2(new_n385), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n498), .A2(new_n505), .A3(new_n454), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT102), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n498), .A2(new_n505), .A3(KEYINPUT102), .A4(new_n454), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n700), .A2(new_n765), .A3(new_n611), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n760), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n763), .A2(new_n508), .A3(new_n453), .A4(new_n764), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n755), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT42), .B1(new_n716), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n759), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n767), .B1(new_n760), .B2(new_n766), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n716), .A2(KEYINPUT42), .A3(new_n770), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(KEYINPUT103), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n218), .ZN(G33));
  NAND2_X1  g591(.A1(new_n668), .A2(KEYINPUT104), .ZN(new_n778));
  INV_X1    g592(.A(new_n769), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n644), .A2(new_n645), .A3(new_n646), .A4(new_n667), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT104), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n716), .A2(new_n778), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  INV_X1    g598(.A(new_n660), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n609), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT43), .B1(new_n684), .B2(new_n637), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n684), .A2(KEYINPUT43), .A3(new_n637), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n508), .ZN(new_n792));
  INV_X1    g606(.A(new_n447), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n450), .A2(new_n451), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n450), .A2(KEYINPUT45), .A3(new_n451), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(G469), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n448), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n793), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n448), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n792), .B(new_n674), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n787), .A4(new_n788), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n791), .A2(new_n803), .A3(new_n765), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  AOI21_X1  g620(.A(new_n792), .B1(new_n801), .B2(new_n802), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(KEYINPUT105), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n763), .A2(new_n764), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n310), .A2(new_n812), .A3(new_n755), .A4(new_n385), .ZN(new_n813));
  XNOR2_X1  g627(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n811), .B(new_n813), .C1(new_n807), .C2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  NAND2_X1  g630(.A1(new_n707), .A2(new_n710), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n455), .B(new_n792), .C1(new_n817), .C2(KEYINPUT49), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n619), .A2(new_n818), .A3(new_n636), .A4(new_n683), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n691), .A2(new_n696), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n817), .A2(KEYINPUT49), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT106), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n819), .A2(new_n385), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n788), .A2(new_n787), .A3(new_n578), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT111), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n812), .A2(new_n792), .A3(new_n817), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n750), .A2(new_n660), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n385), .A2(new_n820), .A3(new_n578), .A4(new_n827), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n619), .A2(new_n637), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n828), .A2(new_n829), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n750), .A2(new_n385), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n683), .A2(new_n455), .A3(new_n711), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n826), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n811), .B1(new_n807), .B2(new_n814), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n817), .A2(new_n508), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n826), .A2(new_n834), .A3(new_n765), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n841), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n826), .A2(new_n834), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n842), .B1(new_n508), .B2(new_n817), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT112), .A4(new_n765), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n824), .B1(new_n840), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n760), .B1(KEYINPUT114), .B2(KEYINPUT48), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n826), .A2(new_n827), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n826), .A2(new_n506), .A3(new_n711), .A4(new_n834), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n684), .A2(new_n636), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n577), .B1(new_n830), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n857), .A2(KEYINPUT113), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT113), .B1(new_n857), .B2(new_n860), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n856), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT51), .B1(new_n845), .B2(new_n846), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n852), .B(new_n863), .C1(new_n840), .C2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n750), .A2(new_n660), .A3(new_n770), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n785), .B1(new_n691), .B2(new_n295), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT109), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n615), .A2(new_n685), .A3(new_n666), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n644), .A2(new_n870), .A3(new_n646), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n769), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n871), .A2(new_n869), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n783), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n772), .A3(new_n775), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n547), .B(new_n685), .C1(new_n602), .C2(new_n603), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n622), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n609), .A3(new_n385), .A4(new_n611), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n606), .A2(new_n661), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT108), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n684), .A2(new_n883), .A3(new_n636), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n881), .A2(new_n882), .A3(new_n738), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n738), .A3(new_n884), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n612), .B1(new_n886), .B2(KEYINPUT108), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n880), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n712), .B1(new_n734), .B2(new_n730), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n717), .A3(new_n751), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n876), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n757), .A2(new_n670), .A3(new_n701), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n642), .B1(new_n741), .B2(new_n742), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n610), .A2(new_n666), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n894), .A2(new_n697), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n892), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n670), .A2(new_n701), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n894), .A2(new_n697), .A3(new_n895), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT52), .A4(new_n757), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n773), .A2(KEYINPUT103), .A3(new_n774), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT103), .B1(new_n773), .B2(new_n774), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n783), .A2(new_n867), .A3(new_n874), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n716), .A2(new_n638), .A3(new_n711), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n717), .A2(new_n735), .A3(new_n907), .A4(new_n751), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n886), .A2(KEYINPUT108), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n613), .A3(new_n885), .ZN(new_n910));
  INV_X1    g724(.A(new_n880), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n906), .A2(new_n901), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n866), .B1(new_n902), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n735), .A2(new_n907), .A3(new_n751), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n773), .A2(new_n774), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n918), .A2(KEYINPUT110), .A3(new_n717), .A4(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT110), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n768), .A2(new_n771), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n908), .B2(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n912), .A2(new_n905), .A3(new_n915), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n920), .A2(new_n923), .A3(new_n924), .A4(new_n901), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n916), .A2(new_n866), .A3(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n865), .A2(new_n917), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(G952), .A2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n823), .B1(new_n927), .B2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n312), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n283), .B1(new_n916), .B2(new_n925), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT56), .B1(new_n932), .B2(G210), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n500), .A2(new_n501), .A3(new_n462), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n485), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT55), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n931), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n932), .A2(G210), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT117), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n937), .A2(KEYINPUT116), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(KEYINPUT116), .ZN(new_n942));
  XOR2_X1   g756(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n939), .A2(new_n940), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n932), .A2(G210), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT117), .B1(new_n947), .B2(new_n944), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n938), .B1(new_n946), .B2(new_n948), .ZN(G51));
  XOR2_X1   g763(.A(new_n448), .B(KEYINPUT57), .Z(new_n950));
  AOI21_X1  g764(.A(new_n866), .B1(new_n916), .B2(new_n925), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n926), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n705), .ZN(new_n953));
  INV_X1    g767(.A(new_n932), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(new_n798), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n930), .B1(new_n953), .B2(new_n955), .ZN(G54));
  INV_X1    g770(.A(new_n599), .ZN(new_n957));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .A4(new_n599), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n959), .A2(new_n931), .A3(new_n960), .ZN(G60));
  XNOR2_X1  g775(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n574), .A2(new_n283), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(new_n964));
  NOR2_X1   g778(.A1(new_n633), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT53), .B1(new_n891), .B2(new_n901), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n901), .A2(new_n920), .A3(new_n923), .A4(new_n924), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT54), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n916), .A2(new_n866), .A3(new_n925), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT119), .B1(new_n971), .B2(new_n930), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n965), .B1(new_n926), .B2(new_n951), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT119), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n974), .A3(new_n931), .ZN(new_n975));
  INV_X1    g789(.A(new_n964), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n926), .B2(new_n917), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n633), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n972), .A2(new_n975), .A3(new_n978), .ZN(G63));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n916), .B2(new_n925), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n366), .A2(new_n368), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n658), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n931), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n985), .A2(KEYINPUT61), .A3(new_n931), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G66));
  NAND2_X1  g805(.A1(new_n890), .A2(new_n312), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT120), .ZN(new_n993));
  INV_X1    g807(.A(G224), .ZN(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n580), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n480), .B(new_n484), .C1(G898), .C2(new_n312), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT121), .Z(new_n998));
  XNOR2_X1  g812(.A(new_n996), .B(new_n998), .ZN(G69));
  NAND3_X1  g813(.A1(new_n803), .A2(new_n716), .A3(new_n894), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n783), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n772), .A3(new_n775), .A4(new_n815), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g818(.A(new_n893), .ZN(new_n1005));
  AOI21_X1  g819(.A(KEYINPUT124), .B1(new_n805), .B2(new_n1005), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n805), .A2(KEYINPUT124), .A3(new_n1005), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1003), .B(new_n1004), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g823(.A(KEYINPUT125), .B1(new_n1009), .B2(new_n1002), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1008), .A2(new_n1010), .A3(new_n312), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n275), .A2(new_n277), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1012), .B(new_n1013), .Z(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(G900), .B2(G953), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(G953), .B1(new_n435), .B2(new_n665), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT123), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n698), .A2(new_n898), .A3(new_n757), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n881), .A2(new_n884), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n674), .B1(new_n1023), .B2(new_n877), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n716), .A3(new_n779), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n805), .A2(new_n815), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(KEYINPUT122), .B1(new_n1021), .B2(KEYINPUT62), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1021), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1027), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n312), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1020), .B1(new_n1032), .B2(new_n1014), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n1016), .A2(new_n1019), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1019), .B1(new_n1016), .B2(new_n1033), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1034), .A2(new_n1035), .ZN(G72));
  NOR2_X1   g850(.A1(new_n279), .A2(new_n254), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1008), .A2(new_n1010), .A3(new_n913), .ZN(new_n1039));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  AOI21_X1  g855(.A(new_n1038), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n279), .A2(new_n254), .ZN(new_n1044));
  OAI211_X1 g858(.A(new_n1027), .B(new_n913), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1044), .B1(new_n1045), .B2(new_n1041), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1038), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1047), .B1(new_n902), .B2(new_n916), .ZN(new_n1048));
  NOR3_X1   g862(.A1(new_n1046), .A2(new_n1048), .A3(new_n930), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1043), .A2(KEYINPUT127), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT127), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n1048), .A2(new_n930), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1046), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1051), .B1(new_n1054), .B2(new_n1042), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1050), .A2(new_n1055), .ZN(G57));
endmodule


