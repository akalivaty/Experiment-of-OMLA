//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n634, new_n637, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT68), .B(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  OR3_X1    g047(.A1(new_n471), .A2(KEYINPUT69), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT69), .B1(new_n471), .B2(new_n472), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n464), .A2(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n464), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n467), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n464), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n467), .A2(new_n464), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(KEYINPUT70), .A3(G124), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n486), .B1(new_n491), .B2(new_n492), .ZN(G162));
  OR2_X1    g068(.A1(new_n470), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n467), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G138), .B1(new_n465), .B2(new_n466), .ZN(new_n500));
  OAI211_X1 g075(.A(KEYINPUT71), .B(KEYINPUT4), .C1(new_n479), .C2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n467), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n502), .A2(G138), .A3(new_n464), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n499), .B1(new_n501), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n506), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(new_n510), .B1(new_n506), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n511), .A2(G88), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n511), .A2(G50), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n520), .A2(new_n522), .B1(G651), .B2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(new_n511), .A2(G51), .A3(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT74), .B1(new_n524), .B2(new_n525), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n514), .A2(new_n532), .A3(new_n515), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n531), .A2(new_n533), .A3(G63), .A4(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n507), .A2(new_n510), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n506), .A2(G651), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n535), .A2(G89), .A3(new_n516), .A4(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  AND4_X1   g114(.A1(new_n530), .A2(new_n534), .A3(new_n537), .A4(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n531), .A2(new_n533), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n535), .A2(G52), .A3(G543), .A4(new_n536), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n535), .A2(G90), .A3(new_n516), .A4(new_n536), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT75), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT75), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND4_X1  g126(.A1(new_n535), .A2(G43), .A3(G543), .A4(new_n536), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n535), .A2(G81), .A3(new_n516), .A4(new_n536), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n531), .A2(new_n533), .A3(G56), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n509), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  NAND4_X1  g141(.A1(new_n535), .A2(G53), .A3(G543), .A4(new_n536), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n511), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n514), .B2(new_n515), .ZN(new_n574));
  AND2_X1   g149(.A1(G78), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n535), .A2(G91), .A3(new_n516), .A4(new_n536), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n571), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n572), .B1(new_n571), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G168), .ZN(G286));
  NAND2_X1  g157(.A1(new_n520), .A2(new_n522), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n528), .A2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G303));
  AOI21_X1  g160(.A(G74), .B1(new_n531), .B2(new_n533), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n586), .A2(KEYINPUT79), .A3(new_n509), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT79), .B1(new_n586), .B2(new_n509), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n511), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n587), .A2(new_n588), .B1(G49), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n511), .A2(G87), .A3(new_n516), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT78), .Z(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(KEYINPUT80), .A3(new_n593), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n526), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g176(.A1(G48), .A2(G543), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n601), .A2(G651), .B1(new_n511), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n511), .A2(G86), .A3(new_n516), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G305));
  NAND3_X1  g180(.A1(new_n511), .A2(G47), .A3(G543), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n511), .A2(G85), .A3(new_n516), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT81), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G72), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G60), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n542), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G651), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n526), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G651), .ZN(new_n622));
  INV_X1    g197(.A(G54), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n589), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n535), .A2(G92), .A3(new_n516), .A4(new_n536), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n618), .B1(G868), .B2(new_n629), .ZN(G284));
  OAI21_X1  g205(.A(new_n618), .B1(G868), .B2(new_n629), .ZN(G321));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  NOR2_X1   g207(.A1(G286), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G299), .B(KEYINPUT82), .Z(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(new_n632), .ZN(G297));
  AOI21_X1  g210(.A(new_n633), .B1(new_n634), .B2(new_n632), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n629), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n629), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g217(.A1(new_n467), .A2(new_n471), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G2100), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  INV_X1    g225(.A(G111), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n653));
  AOI22_X1  g228(.A1(new_n479), .A2(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n652), .B2(new_n653), .ZN(new_n655));
  AOI22_X1  g230(.A1(G123), .A2(new_n488), .B1(new_n482), .B2(G135), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(G2096), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n649), .A2(new_n650), .A3(new_n658), .ZN(G156));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT86), .Z(new_n661));
  XOR2_X1   g236(.A(G2451), .B(G2454), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT14), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2427), .B(G2438), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2430), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT15), .B(G2435), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n668), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n664), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  AND3_X1   g249(.A1(new_n673), .A2(G14), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g251(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2072), .B(G2078), .Z(new_n684));
  INV_X1    g259(.A(new_n677), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n693), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n691), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(new_n594), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT33), .B(G1976), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(G166), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G16), .B2(G22), .ZN(new_n715));
  INV_X1    g290(.A(G1971), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n710), .A2(new_n712), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n707), .A2(G6), .ZN(new_n718));
  INV_X1    g293(.A(G305), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n707), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT32), .B(G1981), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n715), .A2(new_n716), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n713), .A2(new_n717), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  OAI221_X1 g304(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT89), .Z(new_n731));
  AOI22_X1  g306(.A1(G119), .A2(new_n488), .B1(new_n482), .B2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n729), .B1(new_n733), .B2(G29), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT35), .B(G1991), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G1986), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n609), .A2(new_n611), .B1(G651), .B2(new_n615), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(new_n707), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n707), .B2(G24), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n737), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n738), .B2(new_n741), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n726), .A2(new_n727), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT36), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n561), .A2(new_n707), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n707), .B2(G19), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G1341), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(G1341), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n707), .A2(G5), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G301), .B2(G16), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n749), .B(new_n750), .C1(G1961), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G168), .A2(new_n707), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n707), .B2(G21), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n728), .A2(G26), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT28), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n482), .A2(G140), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT92), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n488), .A2(G128), .ZN(new_n763));
  OAI221_X1 g338(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n760), .B1(new_n766), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n757), .B2(new_n756), .ZN(new_n770));
  NOR2_X1   g345(.A1(G4), .A2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT91), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n628), .A2(new_n627), .ZN(new_n773));
  INV_X1    g348(.A(new_n624), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n772), .B1(new_n775), .B2(new_n707), .ZN(new_n776));
  INV_X1    g351(.A(G1348), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT30), .B(G28), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n779), .A2(new_n728), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(G164), .A2(G29), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G27), .B2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n782), .B1(new_n728), .B2(new_n657), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  AND4_X1   g362(.A1(new_n758), .A2(new_n770), .A3(new_n778), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n728), .A2(G35), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n728), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2090), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n777), .B2(new_n776), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n754), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT93), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT25), .ZN(new_n797));
  NAND2_X1  g372(.A1(G115), .A2(G2104), .ZN(new_n798));
  INV_X1    g373(.A(G127), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n467), .B2(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT94), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n464), .B1(new_n800), .B2(KEYINPUT94), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n801), .A2(new_n802), .B1(G139), .B2(new_n482), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G33), .B(new_n804), .S(G29), .Z(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(G2072), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(G2072), .ZN(new_n807));
  INV_X1    g382(.A(G34), .ZN(new_n808));
  AOI21_X1  g383(.A(G29), .B1(new_n808), .B2(KEYINPUT24), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT95), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n808), .A2(KEYINPUT24), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n809), .B2(KEYINPUT95), .ZN(new_n812));
  AOI22_X1  g387(.A1(G160), .A2(G29), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G2084), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n728), .A2(G32), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n816));
  NAND3_X1  g391(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n488), .A2(G129), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n482), .A2(G141), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n821));
  AND4_X1   g396(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n815), .B1(new_n822), .B2(new_n728), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT27), .B(G1996), .Z(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT97), .Z(new_n826));
  NAND4_X1  g401(.A1(new_n806), .A2(new_n807), .A3(new_n814), .A4(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT98), .ZN(new_n828));
  NAND2_X1  g403(.A1(G299), .A2(G16), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n707), .A2(G20), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT23), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1956), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n813), .A2(G2084), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n753), .A2(G1961), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n834), .B(new_n835), .C1(new_n823), .C2(new_n824), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n794), .A2(new_n828), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n745), .A2(new_n840), .ZN(G150));
  INV_X1    g416(.A(G150), .ZN(G311));
  NAND2_X1  g417(.A1(new_n629), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n535), .A2(G55), .A3(G543), .A4(new_n536), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n535), .A2(new_n516), .A3(new_n536), .ZN(new_n846));
  INV_X1    g421(.A(G93), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n531), .A2(new_n533), .A3(G67), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n509), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n559), .B2(new_n560), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n555), .A2(new_n556), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT76), .B1(new_n854), .B2(new_n509), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n848), .A2(new_n851), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n557), .A2(new_n558), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n554), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n844), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT100), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n852), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  XNOR2_X1  g442(.A(new_n804), .B(new_n822), .ZN(new_n868));
  AOI22_X1  g443(.A1(G130), .A2(new_n488), .B1(new_n482), .B2(G142), .ZN(new_n869));
  OAI221_X1 g444(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n733), .B(new_n871), .Z(new_n872));
  OR2_X1    g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G164), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n766), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n645), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n873), .A2(new_n878), .A3(new_n874), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G160), .B(new_n657), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G162), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  INV_X1    g461(.A(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(new_n887), .A3(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g465(.A(new_n859), .B(new_n639), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n775), .B1(new_n579), .B2(new_n580), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n571), .A2(new_n578), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT77), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n571), .A2(new_n572), .A3(new_n578), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n629), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT41), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(new_n892), .B2(new_n896), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n898), .B1(new_n891), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n594), .A2(new_n719), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n591), .A2(new_n593), .A3(G305), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(G290), .A2(G166), .ZN(new_n908));
  NAND2_X1  g483(.A1(G303), .A2(new_n739), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n905), .A2(new_n908), .A3(new_n909), .A4(new_n906), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n903), .A2(new_n904), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(G868), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n903), .B2(new_n904), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT101), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n919), .A2(new_n920), .A3(G868), .A4(new_n915), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n918), .B(new_n921), .C1(G868), .C2(new_n856), .ZN(G295));
  OAI211_X1 g497(.A(new_n918), .B(new_n921), .C1(G868), .C2(new_n856), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n853), .A2(new_n858), .ZN(new_n925));
  NAND2_X1  g500(.A1(G301), .A2(G286), .ZN(new_n926));
  OAI211_X1 g501(.A(G168), .B(new_n545), .C1(new_n549), .C2(new_n548), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n925), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n853), .A2(new_n926), .A3(new_n858), .A4(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n926), .A2(new_n927), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n859), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT104), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n853), .A2(new_n858), .B1(new_n926), .B2(new_n927), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n933), .A2(new_n897), .A3(new_n936), .A4(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n859), .A2(new_n934), .ZN(new_n941));
  OAI22_X1  g516(.A1(new_n899), .A2(new_n900), .B1(new_n941), .B2(new_n937), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n935), .A2(new_n931), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n945), .B(KEYINPUT103), .C1(new_n899), .C2(new_n900), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n940), .A2(new_n944), .A3(new_n913), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n886), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n911), .A2(KEYINPUT106), .A3(new_n912), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT106), .B1(new_n911), .B2(new_n912), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n936), .A2(new_n939), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n901), .B1(new_n954), .B2(new_n933), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n935), .A2(new_n897), .A3(new_n931), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n951), .B(new_n952), .C1(new_n955), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n929), .B1(new_n925), .B2(new_n928), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n936), .B(new_n939), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n899), .A2(new_n900), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n957), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  INV_X1    g539(.A(new_n912), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n905), .A2(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n911), .A2(KEYINPUT106), .A3(new_n912), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT107), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n948), .B1(new_n958), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n924), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n947), .A2(new_n886), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n959), .A2(new_n960), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n962), .B1(new_n975), .B2(new_n953), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n956), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n952), .B1(new_n977), .B2(new_n951), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n963), .A2(new_n969), .A3(KEYINPUT107), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n940), .A2(new_n944), .A3(new_n946), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n983), .A2(new_n951), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(new_n948), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n985), .B2(new_n972), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n973), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT43), .B1(new_n984), .B2(new_n948), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n980), .B2(KEYINPUT43), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(G397));
  XOR2_X1   g567(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n993));
  NAND3_X1  g568(.A1(G303), .A2(G8), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  NOR2_X1   g570(.A1(G166), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(KEYINPUT112), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n994), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(G164), .B2(G1384), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n475), .A2(G40), .A3(new_n480), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(KEYINPUT111), .A3(new_n716), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n876), .A2(new_n1008), .A3(new_n1000), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1010));
  INV_X1    g585(.A(G2090), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1005), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n1006), .B2(new_n716), .ZN(new_n1014));
  OAI211_X1 g589(.A(G8), .B(new_n999), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT113), .B(G8), .Z(new_n1016));
  NOR2_X1   g591(.A1(G164), .A2(G1384), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n1005), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT115), .B1(G305), .B2(G1981), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n603), .A2(new_n1021), .A3(new_n1022), .A4(new_n604), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT116), .B(G86), .Z(new_n1025));
  OAI21_X1  g600(.A(new_n603), .B1(new_n846), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G1981), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT117), .B(KEYINPUT49), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1019), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1024), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n596), .A2(new_n1032), .A3(new_n597), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n591), .A2(G1976), .A3(new_n593), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1034), .A2(new_n1018), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1030), .A2(new_n1031), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1018), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT114), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1041), .A3(KEYINPUT52), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(G303), .A2(G8), .A3(new_n993), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n998), .B1(G303), .B2(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1009), .A2(new_n1005), .A3(new_n1010), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1047), .A2(new_n1011), .B1(new_n1006), .B2(new_n716), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1046), .B1(new_n1048), .B2(new_n1016), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1015), .A2(new_n1037), .A3(new_n1043), .A4(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1001), .A2(new_n1003), .A3(new_n785), .A4(new_n1005), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(G2078), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n475), .A2(new_n480), .A3(G40), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1003), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1009), .A2(new_n1005), .A3(new_n1010), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT125), .B(G1961), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1053), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G171), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1050), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1016), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT120), .B(G2084), .Z(new_n1065));
  NAND4_X1  g640(.A1(new_n1009), .A2(new_n1010), .A3(new_n1005), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1004), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1966), .B1(new_n1068), .B2(new_n1003), .ZN(new_n1069));
  OAI211_X1 g644(.A(G286), .B(new_n1064), .C1(new_n1067), .C2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G168), .A2(new_n1016), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1006), .A2(new_n757), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n995), .B1(new_n1072), .B2(new_n1066), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1070), .B(KEYINPUT51), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1066), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1064), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1071), .A2(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1063), .A2(new_n1081), .A3(KEYINPUT126), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1018), .A3(new_n1031), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1041), .B1(new_n1038), .B2(KEYINPUT52), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT114), .B(new_n1035), .C1(new_n1034), .C2(new_n1018), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1062), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1015), .A3(new_n1049), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT62), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1083), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1074), .A2(KEYINPUT62), .A3(new_n1078), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1082), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1075), .A2(G168), .A3(new_n1064), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1050), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT121), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1102), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1046), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1015), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(new_n1098), .C1(new_n1050), .C2(new_n1099), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1101), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1024), .B(KEYINPUT119), .ZN(new_n1110));
  NOR2_X1   g685(.A1(G288), .A2(G1976), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1111), .B2(new_n1086), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n1018), .B(KEYINPUT118), .Z(new_n1113));
  OAI22_X1  g688(.A1(new_n1102), .A2(new_n1015), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1053), .A2(new_n1060), .A3(G301), .A4(new_n1057), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n876), .A2(KEYINPUT109), .A3(new_n1000), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT109), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(G164), .B2(G1384), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1002), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1056), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1053), .A2(new_n1060), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT54), .B(new_n1115), .C1(new_n1121), .C2(G301), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1124));
  NAND4_X1  g699(.A1(new_n1053), .A2(new_n1060), .A3(new_n1120), .A4(G301), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1062), .B2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1123), .A2(new_n1050), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1956), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1058), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1068), .A2(new_n1003), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1132), .A2(KEYINPUT122), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n893), .B(KEYINPUT57), .Z(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1132), .B2(KEYINPUT122), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1129), .A2(new_n1134), .A3(new_n1131), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1004), .A2(G164), .A3(G1384), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1058), .A2(new_n777), .B1(new_n768), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n775), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1133), .A2(new_n1135), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1058), .A2(new_n777), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n768), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1141), .A2(new_n1142), .A3(KEYINPUT60), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT58), .B(G1341), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1006), .A2(G1996), .B1(new_n1137), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n561), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1143), .A2(new_n775), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1129), .A2(new_n1134), .A3(new_n1131), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1134), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n775), .B1(new_n1138), .B2(KEYINPUT60), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1149), .A2(new_n1153), .A3(new_n1154), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1136), .A2(KEYINPUT61), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1140), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1114), .B1(new_n1127), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1097), .A2(new_n1109), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n766), .B(new_n768), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n822), .B(G1996), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1119), .A2(new_n1004), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1170), .A2(KEYINPUT110), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(KEYINPUT110), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n735), .B1(new_n731), .B2(new_n732), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n733), .A2(new_n736), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1169), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1169), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n739), .A2(new_n738), .ZN(new_n1178));
  NAND2_X1  g753(.A1(G290), .A2(G1986), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1165), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n762), .A2(new_n768), .A3(new_n765), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1177), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT48), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1176), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1177), .B1(new_n1166), .B2(new_n822), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT127), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1177), .A2(G1996), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT46), .ZN(new_n1192));
  OR3_X1    g767(.A1(new_n1190), .A2(new_n1192), .A3(KEYINPUT47), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT47), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n1185), .B(new_n1188), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1182), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g771(.A1(G229), .A2(new_n462), .A3(new_n675), .A4(G227), .ZN(new_n1198));
  NAND3_X1  g772(.A1(new_n989), .A2(new_n1198), .A3(new_n889), .ZN(G225));
  INV_X1    g773(.A(G225), .ZN(G308));
endmodule


