//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  XNOR2_X1  g0008(.A(KEYINPUT65), .B(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n202), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n216), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n215), .B(new_n219), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  AND2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G223), .A3(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  INV_X1    g0053(.A(G222), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT70), .B(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(new_n248), .A3(new_n250), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n252), .B1(new_n253), .B2(new_n251), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(new_n264), .A3(G274), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  AND2_X1   g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n263), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(new_n262), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n266), .A2(new_n271), .B1(G226), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n259), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G200), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT75), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n259), .A2(G190), .A3(new_n276), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(KEYINPUT75), .A3(G200), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n210), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT71), .ZN(new_n287));
  INV_X1    g0087(.A(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(new_n247), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n209), .A2(G33), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n203), .A2(G20), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(KEYINPUT72), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G1), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n285), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n272), .A2(G20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G50), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n307), .A2(new_n309), .B1(G50), .B2(new_n304), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n301), .A2(KEYINPUT9), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT9), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n300), .B2(new_n310), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n283), .B(new_n315), .C1(new_n316), .C2(KEYINPUT10), .ZN(new_n317));
  INV_X1    g0117(.A(G238), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT70), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n251), .B1(new_n318), .B2(new_n319), .C1(new_n230), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n248), .A2(new_n250), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n264), .B1(new_n325), .B2(new_n206), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n324), .A2(new_n326), .B1(G244), .B2(new_n275), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n266), .A2(new_n271), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n306), .A2(G77), .A3(new_n308), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G77), .B2(new_n304), .ZN(new_n333));
  XOR2_X1   g0133(.A(KEYINPUT8), .B(G58), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT65), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G20), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n334), .A2(new_n291), .B1(new_n338), .B2(G77), .ZN(new_n339));
  XOR2_X1   g0139(.A(KEYINPUT15), .B(G87), .Z(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(G33), .A3(new_n209), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n286), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n333), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n327), .A2(new_n328), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n331), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n349), .B2(new_n345), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(KEYINPUT73), .B1(new_n351), .B2(new_n329), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT73), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n329), .A2(G169), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(new_n343), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n348), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n280), .A2(new_n281), .A3(new_n316), .A4(new_n282), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT10), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n312), .A2(new_n314), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n301), .A2(new_n311), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n277), .A2(new_n349), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n363), .C1(G179), .C2(new_n277), .ZN(new_n364));
  AND4_X1   g0164(.A1(new_n317), .A2(new_n356), .A3(new_n361), .A4(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT79), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n249), .B2(G33), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n247), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n250), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n367), .B1(new_n371), .B2(new_n209), .ZN(new_n372));
  INV_X1    g0172(.A(G68), .ZN(new_n373));
  NOR2_X1   g0173(.A1(KEYINPUT7), .A2(G20), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n325), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n289), .B2(new_n290), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G58), .A2(G68), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n288), .B1(new_n212), .B2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n366), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n249), .A2(KEYINPUT78), .A3(G33), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT78), .B1(new_n249), .B2(G33), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n248), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n335), .A2(new_n337), .A3(new_n367), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n373), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n249), .A2(G33), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT78), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n247), .B2(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n249), .A2(KEYINPUT78), .A3(G33), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT7), .B1(new_n393), .B2(G20), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n378), .A2(new_n380), .A3(new_n366), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n286), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n382), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n320), .A2(new_n322), .A3(G223), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G226), .A2(G1698), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n393), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n264), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n264), .A2(G232), .A3(new_n273), .ZN(new_n405));
  AND4_X1   g0205(.A1(new_n270), .A2(new_n262), .A3(new_n264), .A4(G274), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n270), .B1(new_n269), .B2(new_n262), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n330), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n405), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n266), .B2(new_n271), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n401), .A2(new_n393), .B1(G33), .B2(G87), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n346), .C1(new_n264), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n295), .B1(new_n272), .B2(G20), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n306), .A2(new_n415), .B1(new_n305), .B2(new_n295), .ZN(new_n416));
  NAND2_X1  g0216(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n417));
  AND4_X1   g0217(.A1(new_n398), .A2(new_n414), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n419));
  INV_X1    g0219(.A(new_n416), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n382), .B2(new_n397), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(new_n421), .B2(new_n414), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n375), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n371), .A2(new_n209), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(G68), .C1(new_n425), .C2(new_n367), .ZN(new_n426));
  INV_X1    g0226(.A(new_n381), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT16), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n367), .B1(new_n385), .B2(new_n288), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n393), .B2(new_n386), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n396), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n285), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n416), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n404), .B2(new_n408), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n411), .B(G179), .C1(new_n264), .C2(new_n412), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g0236(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n398), .A2(new_n416), .B1(new_n434), .B2(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(KEYINPUT80), .A2(KEYINPUT18), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT82), .ZN(new_n442));
  OR3_X1    g0242(.A1(new_n423), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n423), .B2(new_n441), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n294), .A2(new_n253), .B1(new_n288), .B2(G68), .ZN(new_n445));
  INV_X1    g0245(.A(G50), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n292), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n285), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT11), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OR3_X1    g0250(.A1(new_n304), .A2(KEYINPUT12), .A3(G68), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT12), .B1(new_n304), .B2(G68), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n373), .B1(new_n272), .B2(G20), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n451), .A2(new_n452), .B1(new_n306), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n448), .B2(new_n449), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n266), .A2(new_n271), .B1(G238), .B2(new_n275), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n320), .A2(new_n322), .A3(G226), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G232), .A2(G1698), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n325), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G97), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n258), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT13), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n457), .B2(new_n463), .ZN(new_n467));
  OAI21_X1  g0267(.A(G169), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT14), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT14), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(G169), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n458), .A2(new_n459), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n251), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n264), .B1(new_n474), .B2(new_n461), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n406), .A2(new_n407), .B1(new_n318), .B2(new_n274), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT76), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT76), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n457), .A2(new_n463), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(KEYINPUT13), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n465), .A2(G179), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT77), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT77), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n456), .B1(new_n472), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(G200), .B1(new_n466), .B2(new_n467), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n456), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n465), .A2(G190), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n457), .A2(new_n463), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n464), .B1(new_n491), .B2(KEYINPUT76), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n479), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  AND4_X1   g0295(.A1(new_n365), .A2(new_n443), .A3(new_n444), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT86), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n320), .A2(new_n322), .A3(G257), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G264), .A2(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(new_n393), .B1(G303), .B2(new_n325), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n502), .B2(new_n264), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n325), .A2(G303), .ZN(new_n504));
  INV_X1    g0304(.A(new_n500), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n255), .B2(G257), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n506), .B2(new_n385), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(KEYINPUT86), .A3(new_n258), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n261), .A2(G1), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G270), .A3(new_n264), .ZN(new_n514));
  XNOR2_X1  g0314(.A(KEYINPUT5), .B(G41), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n269), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n517), .B1(new_n514), .B2(new_n516), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(G200), .B1(new_n509), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n247), .A2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n335), .A2(new_n337), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT20), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n284), .A2(new_n210), .B1(G20), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(KEYINPUT88), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n272), .A2(new_n527), .A3(G13), .A4(G20), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n272), .A2(G33), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n286), .A2(new_n304), .A3(G116), .A4(new_n532), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT88), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n525), .A2(new_n528), .B1(new_n535), .B2(KEYINPUT20), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n535), .B2(KEYINPUT20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n514), .A2(new_n516), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT85), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n518), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(new_n503), .A3(G190), .A4(new_n508), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n522), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n508), .A3(new_n503), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n349), .B1(new_n534), .B2(new_n537), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT21), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(KEYINPUT21), .A3(new_n546), .ZN(new_n550));
  INV_X1    g0350(.A(new_n509), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n551), .A2(G179), .A3(new_n542), .A4(new_n538), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n544), .A2(new_n549), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  INV_X1    g0354(.A(G87), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n393), .A2(new_n209), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n554), .B1(new_n325), .B2(new_n555), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G116), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n288), .B1(new_n560), .B2(KEYINPUT23), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n338), .A2(new_n562), .B1(KEYINPUT23), .B2(G107), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n557), .A2(new_n558), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n564), .A2(KEYINPUT24), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(KEYINPUT24), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n285), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT25), .B1(new_n305), .B2(new_n206), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n286), .A2(new_n304), .A3(new_n532), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n569), .A2(new_n570), .B1(new_n571), .B2(new_n206), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G257), .A2(G1698), .ZN(new_n574));
  INV_X1    g0374(.A(G250), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n323), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n393), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G294), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n264), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n513), .A2(G264), .A3(new_n264), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n516), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n579), .A2(G190), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n255), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n578), .B1(new_n583), .B2(new_n385), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT89), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n513), .A2(KEYINPUT89), .A3(G264), .A4(new_n264), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n584), .A2(new_n258), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(G200), .B1(new_n588), .B2(new_n516), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n567), .B(new_n573), .C1(new_n582), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n258), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n586), .A2(new_n587), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(G179), .A3(new_n592), .A4(new_n516), .ZN(new_n593));
  OAI21_X1  g0393(.A(G169), .B1(new_n579), .B2(new_n581), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n563), .A2(new_n561), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT24), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n597), .A3(new_n557), .A4(new_n558), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n564), .A2(KEYINPUT24), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n286), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n595), .B1(new_n600), .B2(new_n572), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n248), .A2(new_n250), .A3(G250), .A4(G1698), .ZN(new_n603));
  NAND2_X1  g0403(.A1(KEYINPUT4), .A2(G244), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n524), .B(new_n603), .C1(new_n256), .C2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n320), .A2(new_n322), .A3(G244), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT4), .B1(new_n393), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n258), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n516), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n258), .B1(new_n510), .B2(new_n515), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(G257), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(G190), .A3(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n372), .A2(new_n206), .A3(new_n375), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n205), .A3(G107), .ZN(new_n615));
  XNOR2_X1  g0415(.A(G97), .B(G107), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n617), .A2(new_n209), .B1(new_n253), .B2(new_n292), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n285), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  MUX2_X1   g0419(.A(new_n304), .B(new_n571), .S(G97), .Z(new_n620));
  AND3_X1   g0420(.A1(new_n612), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n608), .A2(new_n611), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G200), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT83), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n330), .B1(new_n608), .B2(new_n611), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT83), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n621), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n340), .A2(new_n304), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n393), .A2(G68), .A3(new_n209), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT19), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n461), .A2(new_n631), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n338), .A2(new_n632), .B1(G87), .B2(new_n207), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n335), .A2(new_n337), .A3(G33), .A4(G97), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n631), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n629), .B1(new_n636), .B2(new_n285), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n306), .A2(new_n532), .A3(new_n340), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n269), .A2(new_n510), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n264), .B(G250), .C1(G1), .C2(new_n261), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(G244), .A2(G1698), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n323), .B2(new_n318), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n560), .B1(new_n645), .B2(new_n393), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n643), .B1(new_n646), .B2(new_n264), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n349), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n255), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n559), .B1(new_n649), .B2(new_n385), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n642), .B1(new_n650), .B2(new_n258), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n351), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n639), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n571), .A2(new_n555), .ZN(new_n654));
  AOI211_X1 g0454(.A(new_n629), .B(new_n654), .C1(new_n636), .C2(new_n285), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(G190), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n647), .A2(G200), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n608), .A2(new_n351), .A3(new_n611), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT84), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT84), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n608), .A2(new_n662), .A3(new_n351), .A4(new_n611), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n349), .A2(new_n622), .B1(new_n619), .B2(new_n620), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n628), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  NOR4_X1   g0467(.A1(new_n497), .A2(new_n553), .A3(new_n602), .A4(new_n667), .ZN(G372));
  INV_X1    g0468(.A(new_n364), .ZN(new_n669));
  INV_X1    g0469(.A(new_n423), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n344), .B(KEYINPUT73), .C1(G169), .C2(new_n329), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n329), .A2(new_n351), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n355), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n494), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n670), .B1(new_n487), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n434), .A2(new_n435), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n421), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n433), .A2(KEYINPUT90), .A3(new_n436), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT18), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(KEYINPUT18), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n317), .A2(new_n361), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n669), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n626), .B(new_n624), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n688), .A2(new_n621), .B1(new_n664), .B2(new_n665), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n549), .A2(new_n601), .A3(new_n550), .A4(new_n552), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n590), .A4(new_n659), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n659), .A2(KEYINPUT26), .A3(new_n664), .A4(new_n665), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n664), .A2(new_n665), .A3(new_n653), .A4(new_n658), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT26), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n691), .A2(new_n696), .A3(new_n653), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n687), .B1(new_n497), .B2(new_n698), .ZN(G369));
  NAND2_X1  g0499(.A1(new_n209), .A2(new_n303), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n539), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n553), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n552), .A2(new_n550), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n549), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n707), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G330), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n602), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n705), .B1(new_n600), .B2(new_n572), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n601), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n705), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n705), .B1(new_n709), .B2(new_n549), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n725), .A2(new_n717), .B1(new_n720), .B2(new_n706), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n217), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G41), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G1), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n555), .A2(new_n205), .A3(new_n206), .A4(new_n527), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(new_n213), .B2(new_n730), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT92), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n696), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n628), .A2(new_n659), .A3(new_n666), .A4(new_n590), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n549), .A2(new_n601), .A3(new_n550), .A4(new_n552), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n653), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(KEYINPUT29), .B(new_n706), .C1(new_n737), .C2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT91), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n697), .A2(new_n706), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(KEYINPUT91), .B(KEYINPUT29), .C1(new_n697), .C2(new_n706), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n588), .A2(new_n651), .A3(new_n608), .A4(new_n611), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n542), .A2(new_n503), .A3(G179), .A4(new_n508), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n651), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n588), .A2(new_n516), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n545), .A2(new_n752), .A3(new_n753), .A4(new_n622), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n749), .A2(new_n750), .A3(new_n748), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n705), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(KEYINPUT31), .B(new_n705), .C1(new_n755), .C2(new_n756), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR4_X1   g0561(.A1(new_n667), .A2(new_n553), .A3(new_n602), .A4(new_n705), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n714), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n747), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n734), .B1(new_n767), .B2(G1), .ZN(G364));
  NOR2_X1   g0568(.A1(new_n338), .A2(new_n302), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n731), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n713), .A2(new_n714), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n716), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT93), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n351), .A2(new_n330), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n338), .A2(G190), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n351), .A2(G200), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n338), .A2(G190), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G50), .A2(new_n779), .B1(new_n782), .B2(G58), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n209), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n780), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n785), .A2(KEYINPUT97), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(KEYINPUT97), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n783), .B1(new_n788), .B2(new_n253), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT98), .Z(new_n790));
  INV_X1    g0590(.A(new_n784), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n791), .A2(G179), .A3(new_n330), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G107), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G179), .A2(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT99), .B(G159), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT32), .Z(new_n804));
  NOR4_X1   g0604(.A1(new_n288), .A2(new_n346), .A3(new_n330), .A4(G179), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n251), .B1(new_n806), .B2(new_n555), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n338), .B1(new_n346), .B2(new_n799), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n205), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n784), .A2(new_n777), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n807), .B(new_n810), .C1(G68), .C2(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n790), .A2(new_n797), .A3(new_n804), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n800), .B(KEYINPUT102), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n796), .A2(G283), .B1(new_n815), .B2(G329), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT103), .Z(new_n817));
  AOI22_X1  g0617(.A1(new_n779), .A2(G326), .B1(G294), .B2(new_n808), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT101), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n782), .A2(G322), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n251), .B1(new_n805), .B2(G303), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n785), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G311), .A2(new_n825), .B1(new_n812), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n820), .A2(new_n821), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n814), .B1(new_n817), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n349), .A2(KEYINPUT95), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n288), .B1(KEYINPUT95), .B2(new_n349), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n210), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT96), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(G13), .A2(G33), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(G20), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n728), .A2(new_n325), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT94), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G355), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(G116), .B2(new_n217), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n393), .A2(new_n728), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(G45), .B2(new_n213), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G45), .B2(new_n244), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n839), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n835), .A2(new_n772), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n713), .B2(new_n838), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n776), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  NAND2_X1  g0651(.A1(new_n796), .A2(G68), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n393), .B1(new_n806), .B2(new_n446), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G58), .B2(new_n808), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n811), .A2(new_n293), .B1(new_n856), .B2(new_n778), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT104), .Z(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n859), .B2(new_n781), .C1(new_n788), .C2(new_n801), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT34), .Z(new_n861));
  AOI211_X1 g0661(.A(new_n855), .B(new_n861), .C1(G132), .C2(new_n815), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n251), .B(new_n810), .C1(G107), .C2(new_n805), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n812), .A2(G283), .B1(G294), .B2(new_n782), .ZN(new_n864));
  INV_X1    g0664(.A(G303), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n778), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n796), .A2(G87), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n527), .B2(new_n788), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n866), .B(new_n868), .C1(G311), .C2(new_n815), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n834), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n348), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n344), .A2(new_n705), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n673), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n673), .B2(new_n872), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(new_n837), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n834), .A2(new_n836), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n773), .B1(new_n876), .B2(new_n253), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n870), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n673), .A2(new_n871), .A3(new_n706), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n692), .A2(new_n695), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n879), .B1(new_n740), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n743), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n882), .B2(new_n874), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(new_n765), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n772), .B1(new_n883), .B2(new_n765), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n878), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(G384));
  NOR2_X1   g0687(.A1(new_n769), .A2(new_n272), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n381), .B1(new_n388), .B2(new_n394), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n285), .B(new_n431), .C1(new_n891), .C2(KEYINPUT16), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n703), .B1(new_n892), .B2(new_n416), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n423), .B2(new_n441), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n677), .A2(new_n703), .B1(new_n416), .B2(new_n892), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n398), .A2(new_n414), .A3(new_n416), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n433), .A2(new_n436), .ZN(new_n898));
  INV_X1    g0698(.A(new_n703), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n433), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n421), .A2(new_n414), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n898), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n897), .A2(KEYINPUT106), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n894), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT106), .B1(new_n897), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n890), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n906), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n894), .A4(new_n904), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n667), .ZN(new_n911));
  INV_X1    g0711(.A(new_n553), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n911), .A2(new_n717), .A3(new_n912), .A4(new_n706), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n759), .A3(new_n760), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n480), .A2(new_n484), .A3(new_n481), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n484), .B1(new_n480), .B2(new_n481), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n469), .B(new_n471), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n456), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n494), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT105), .B1(new_n456), .B2(new_n706), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n922), .B(new_n705), .C1(new_n450), .C2(new_n455), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n487), .B2(new_n494), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n914), .A2(new_n874), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n889), .B1(new_n910), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT107), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n874), .B1(new_n761), .B2(new_n762), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(new_n926), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n907), .A2(new_n909), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(KEYINPUT107), .A3(new_n889), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n678), .A2(KEYINPUT18), .A3(new_n679), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT18), .B1(new_n678), .B2(new_n679), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n670), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n900), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n900), .A2(new_n901), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n678), .B2(new_n679), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n903), .B1(new_n945), .B2(new_n902), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT38), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n905), .A2(new_n890), .A3(new_n906), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n925), .B1(new_n919), .B2(new_n920), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n494), .B(new_n924), .C1(new_n917), .C2(new_n918), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n952), .A2(new_n914), .A3(KEYINPUT40), .A4(new_n874), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n938), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n496), .A2(new_n914), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n956), .A2(new_n957), .A3(new_n714), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n673), .A2(new_n705), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n881), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n952), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n910), .ZN(new_n964));
  INV_X1    g0764(.A(new_n684), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n965), .B2(new_n703), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT39), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n947), .B2(new_n948), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n919), .A2(new_n705), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT39), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n496), .B(new_n741), .C1(new_n745), .C2(new_n746), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n687), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n888), .B1(new_n959), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n975), .B2(new_n959), .ZN(new_n977));
  INV_X1    g0777(.A(new_n617), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT35), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(KEYINPUT35), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n979), .A2(G116), .A3(new_n211), .A4(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT36), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n214), .A2(G77), .A3(new_n379), .ZN(new_n983));
  INV_X1    g0783(.A(new_n201), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n373), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(G1), .A3(new_n302), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n977), .A2(new_n982), .A3(new_n986), .ZN(G367));
  NAND2_X1  g0787(.A1(new_n796), .A2(G97), .ZN(new_n988));
  INV_X1    g0788(.A(new_n800), .ZN(new_n989));
  INV_X1    g0789(.A(G317), .ZN(new_n990));
  INV_X1    g0790(.A(G294), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n989), .A2(new_n990), .B1(new_n991), .B2(new_n811), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G107), .B2(new_n808), .ZN(new_n993));
  INV_X1    g0793(.A(G311), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n865), .A2(new_n781), .B1(new_n778), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT46), .B1(new_n805), .B2(G116), .ZN(new_n997));
  NOR4_X1   g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n393), .ZN(new_n998));
  INV_X1    g0798(.A(new_n788), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(G283), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n988), .A2(new_n993), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n800), .A2(G137), .B1(G68), .B2(new_n808), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n779), .A2(G143), .B1(G58), .B2(new_n805), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n812), .A2(new_n802), .B1(G150), .B2(new_n782), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n796), .A2(G77), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n251), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1005), .B1(new_n201), .B2(new_n788), .C1(new_n1007), .C2(KEYINPUT113), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(KEYINPUT113), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1001), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT47), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n834), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n236), .A2(new_n844), .B1(new_n728), .B2(new_n340), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n773), .B1(new_n839), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n706), .A2(new_n655), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n659), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n653), .B2(new_n1016), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n838), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1013), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n771), .A2(new_n272), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n619), .A2(new_n620), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n628), .B(new_n666), .C1(new_n1024), .C2(new_n706), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n664), .A2(new_n665), .A3(new_n705), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT109), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1025), .A2(KEYINPUT109), .A3(new_n1026), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n726), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(KEYINPUT45), .A3(new_n726), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT44), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1031), .B2(new_n726), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n726), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1039), .A2(new_n1029), .A3(KEYINPUT44), .A4(new_n1030), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1042), .A2(KEYINPUT110), .A3(new_n724), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1034), .A2(new_n1035), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT110), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n723), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n722), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT111), .B1(new_n1048), .B2(new_n725), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT111), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n725), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n722), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1049), .B(new_n1052), .C1(new_n602), .C2(new_n1051), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(new_n715), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n766), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n729), .B(KEYINPUT41), .Z(new_n1056));
  OAI21_X1  g0856(.A(new_n1023), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1018), .A2(KEYINPUT43), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1051), .A2(new_n602), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1031), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT42), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT42), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1031), .A2(new_n1062), .A3(new_n1059), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1031), .A2(new_n720), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n705), .B1(new_n1065), .B2(new_n666), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1058), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1018), .A2(KEYINPUT43), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT108), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n723), .A2(new_n1031), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1069), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1072), .B(new_n1058), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1071), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1057), .A2(KEYINPUT112), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT112), .B1(new_n1057), .B2(new_n1076), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1022), .B1(new_n1078), .B2(new_n1079), .ZN(G387));
  NAND2_X1  g0880(.A1(new_n233), .A2(G45), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1081), .A2(new_n844), .B1(new_n732), .B2(new_n841), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT50), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n334), .B2(new_n446), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n295), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n261), .B1(new_n373), .B2(new_n253), .ZN(new_n1086));
  NOR4_X1   g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n732), .A4(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1082), .A2(new_n1087), .B1(G107), .B2(new_n217), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n773), .B1(new_n1088), .B2(new_n839), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1048), .B2(new_n1019), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n989), .A2(new_n293), .B1(new_n446), .B2(new_n781), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n334), .B2(new_n812), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n393), .B1(new_n806), .B2(new_n253), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G68), .B2(new_n825), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n340), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n809), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G159), .B2(new_n779), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n988), .A2(new_n1092), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n393), .B1(new_n800), .B2(G326), .ZN(new_n1099));
  INV_X1    g0899(.A(G283), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n809), .A2(new_n1100), .B1(new_n806), .B2(new_n991), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n811), .A2(new_n994), .B1(new_n990), .B2(new_n781), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G322), .B2(new_n779), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n788), .B2(new_n865), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT48), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1101), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1105), .B2(new_n1104), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT49), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1099), .B1(new_n527), .B2(new_n795), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1098), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1090), .B1(new_n834), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1023), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1054), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1054), .A2(new_n767), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n729), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1054), .A2(new_n767), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(G393));
  XNOR2_X1  g0918(.A(new_n724), .B(new_n1044), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1116), .B2(new_n1023), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n241), .A2(new_n844), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n839), .B1(new_n205), .B2(new_n217), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n772), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n812), .A2(G303), .B1(G116), .B2(new_n808), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n991), .B2(new_n785), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT114), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n994), .A2(new_n781), .B1(new_n778), .B2(new_n990), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT52), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n325), .B1(new_n806), .B2(new_n1100), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n800), .B2(G322), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1126), .A2(new_n797), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT115), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n393), .B1(new_n806), .B2(new_n373), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n989), .A2(new_n859), .B1(new_n201), .B2(new_n811), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(G77), .C2(new_n808), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n293), .A2(new_n778), .B1(new_n781), .B2(new_n377), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT51), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n999), .A2(new_n334), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n867), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1131), .A2(KEYINPUT115), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1132), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1123), .B1(new_n1141), .B2(new_n834), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1031), .B2(new_n1019), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1043), .A2(new_n1046), .A3(new_n729), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n1115), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1120), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G390));
  INV_X1    g0947(.A(KEYINPUT116), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n914), .A2(G330), .A3(new_n874), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n933), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n969), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n947), .B2(new_n948), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n706), .B(new_n874), .C1(new_n737), .C2(new_n740), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n961), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1152), .B1(new_n1154), .B2(new_n952), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n968), .A2(new_n970), .B1(new_n963), .B2(new_n1151), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1150), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n900), .B1(new_n684), .B2(new_n670), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n946), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n890), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n969), .B1(new_n1160), .B2(new_n909), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n880), .B2(KEYINPUT92), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n740), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n705), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n960), .B1(new_n1165), .B2(new_n874), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1161), .B1(new_n1166), .B2(new_n933), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n960), .B1(new_n697), .B2(new_n879), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1151), .B1(new_n1168), .B2(new_n933), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT39), .B1(new_n1160), .B2(new_n909), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n970), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n764), .A2(new_n952), .A3(new_n874), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1167), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1157), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1148), .B1(new_n1175), .B2(new_n1023), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1157), .A2(new_n1174), .A3(KEYINPUT116), .A4(new_n1113), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n496), .A2(new_n764), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n973), .A2(new_n687), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n952), .B1(new_n764), .B2(new_n874), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n962), .B1(new_n1181), .B2(new_n1150), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1149), .A2(new_n933), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1166), .A2(new_n1173), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1175), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1157), .A2(new_n1174), .A3(new_n1180), .A4(new_n1185), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n729), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n836), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT54), .B(G143), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n999), .A2(new_n1192), .B1(G137), .B2(new_n812), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1194), .A2(KEYINPUT117), .B1(G159), .B2(new_n808), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(KEYINPUT117), .B2(new_n1194), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT118), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT53), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n806), .B2(new_n293), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n805), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1199), .A2(new_n1200), .B1(new_n782), .B2(G132), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n325), .B1(new_n779), .B2(G128), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G125), .B2(new_n815), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n201), .B2(new_n795), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1197), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n815), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n852), .B1(new_n991), .B2(new_n1207), .C1(new_n205), .C2(new_n788), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n325), .B1(new_n806), .B2(new_n555), .C1(new_n809), .C2(new_n253), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G116), .A2(new_n782), .B1(new_n779), .B2(G283), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n206), .B2(new_n811), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT119), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n834), .B1(new_n1206), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n773), .B1(new_n876), .B2(new_n295), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1190), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1178), .A2(new_n1189), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT120), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1178), .A2(new_n1189), .A3(KEYINPUT120), .A4(new_n1216), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(G378));
  INV_X1    g1021(.A(KEYINPUT57), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1188), .B2(new_n1180), .ZN(new_n1223));
  OAI21_X1  g1023(.A(G330), .B1(new_n949), .B2(new_n953), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT107), .B1(new_n936), .B2(new_n889), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n930), .B(KEYINPUT40), .C1(new_n934), .C2(new_n935), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n362), .A2(new_n899), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n686), .A2(new_n364), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n317), .A2(new_n361), .A3(new_n364), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n362), .A3(new_n899), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1228), .A2(new_n1236), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n966), .A2(new_n971), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1236), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n938), .A2(new_n1225), .A3(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1238), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1223), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1239), .B1(new_n938), .B2(new_n1225), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1224), .B(new_n1236), .C1(new_n931), .C2(new_n937), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n972), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1246), .A2(new_n1247), .B1(new_n1180), .B2(new_n1188), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n729), .B(new_n1243), .C1(new_n1248), .C2(KEYINPUT57), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1236), .A2(new_n836), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n834), .A2(new_n984), .A3(new_n836), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n796), .A2(G58), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1100), .B2(new_n1207), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n393), .A2(G41), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n527), .B2(new_n778), .C1(new_n811), .C2(new_n205), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n808), .A2(G68), .B1(new_n805), .B2(G77), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1257), .B1(new_n206), .B2(new_n781), .C1(new_n1095), .C2(new_n785), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1254), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1259), .A2(KEYINPUT58), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n796), .A2(new_n802), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n812), .A2(G132), .B1(G128), .B2(new_n782), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n825), .A2(G137), .B1(G125), .B2(new_n779), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n808), .A2(G150), .B1(new_n805), .B2(new_n1192), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(KEYINPUT59), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(KEYINPUT59), .ZN(new_n1267));
  AOI211_X1 g1067(.A(G33), .B(G41), .C1(new_n800), .C2(G124), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1261), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1259), .A2(KEYINPUT58), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1255), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1271), .B(new_n446), .C1(G33), .C2(G41), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1260), .A2(new_n1269), .A3(new_n1270), .A4(new_n1272), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n773), .B(new_n1252), .C1(new_n1273), .C2(new_n834), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1250), .A2(new_n1113), .B1(new_n1251), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1249), .A2(new_n1275), .ZN(G375));
  INV_X1    g1076(.A(new_n1185), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n952), .A2(new_n837), .ZN(new_n1278));
  OAI221_X1 g1078(.A(new_n1006), .B1(new_n865), .B2(new_n1207), .C1(new_n206), .C2(new_n788), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n251), .B(new_n1096), .C1(G97), .C2(new_n805), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n812), .A2(G116), .B1(G283), .B2(new_n782), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(new_n991), .C2(new_n778), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G150), .A2(new_n825), .B1(new_n812), .B2(new_n1192), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n393), .B1(new_n806), .B2(new_n377), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(G50), .B2(new_n808), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G132), .A2(new_n779), .B1(new_n782), .B2(G137), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1283), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G128), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1253), .B1(new_n1288), .B2(new_n1207), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n1279), .A2(new_n1282), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n834), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n773), .B1(new_n876), .B2(new_n373), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n1277), .A2(new_n1023), .B1(new_n1278), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n973), .A2(new_n687), .A3(new_n1179), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1277), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1056), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1186), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1295), .A2(new_n1299), .ZN(G381));
  AND2_X1   g1100(.A1(new_n1249), .A2(new_n1275), .ZN(new_n1301));
  INV_X1    g1101(.A(G387), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1217), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1146), .A2(new_n886), .ZN(new_n1304));
  NOR4_X1   g1104(.A1(new_n1304), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .A4(new_n1305), .ZN(G407));
  NAND3_X1  g1106(.A1(new_n1301), .A2(new_n704), .A3(new_n1303), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(G407), .A2(G213), .A3(new_n1307), .ZN(G409));
  NAND4_X1  g1108(.A1(new_n1249), .A2(new_n1219), .A3(new_n1220), .A4(new_n1275), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1188), .A2(new_n1180), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1250), .A2(new_n1298), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1275), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1303), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1186), .A2(KEYINPUT60), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1297), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1296), .A2(KEYINPUT60), .A3(new_n1182), .A4(new_n1184), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n729), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G384), .B1(new_n1318), .B2(new_n1295), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n729), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1320), .B1(new_n1315), .B2(new_n1297), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1321), .A2(new_n886), .A3(new_n1294), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1319), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(G213), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(G343), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1314), .A2(new_n1323), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(KEYINPUT121), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1325), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT121), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n1323), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1328), .A2(new_n1329), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT122), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1325), .A2(G2897), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1337), .B1(new_n1319), .B2(new_n1322), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1318), .A2(G384), .A3(new_n1295), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n886), .B1(new_n1321), .B2(new_n1294), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(G2897), .A4(new_n1325), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1338), .A2(KEYINPUT123), .A3(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT123), .B1(new_n1338), .B2(new_n1341), .ZN(new_n1343));
  NOR3_X1   g1143(.A1(new_n1330), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(G393), .B(new_n850), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1057), .A2(new_n1076), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT112), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1077), .ZN(new_n1350));
  AOI21_X1  g1150(.A(G390), .B1(new_n1350), .B2(new_n1022), .ZN(new_n1351));
  AOI211_X1 g1151(.A(new_n1021), .B(new_n1146), .C1(new_n1349), .C2(new_n1077), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1346), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT61), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G387), .A2(new_n1146), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1350), .A2(new_n1022), .A3(G390), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1355), .A2(new_n1345), .A3(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1353), .A2(new_n1354), .A3(new_n1357), .ZN(new_n1358));
  NOR3_X1   g1158(.A1(new_n1336), .A2(new_n1344), .A3(new_n1358), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1328), .A2(KEYINPUT122), .A3(new_n1329), .A4(new_n1332), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1335), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1353), .A2(KEYINPUT125), .A3(new_n1357), .ZN(new_n1362));
  AOI21_X1  g1162(.A(KEYINPUT125), .B1(new_n1353), .B2(new_n1357), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  AND2_X1   g1164(.A1(new_n1338), .A2(new_n1341), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1354), .B1(new_n1330), .B2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(KEYINPUT124), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT124), .ZN(new_n1368));
  OAI211_X1 g1168(.A(new_n1368), .B(new_n1354), .C1(new_n1330), .C2(new_n1365), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1327), .A2(KEYINPUT62), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1367), .A2(new_n1369), .A3(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(KEYINPUT62), .B1(new_n1328), .B2(new_n1332), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1364), .B1(new_n1371), .B2(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1361), .A2(new_n1373), .ZN(G405));
  NAND2_X1  g1174(.A1(G375), .A2(new_n1303), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT126), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1309), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1377));
  INV_X1    g1177(.A(new_n1377), .ZN(new_n1378));
  INV_X1    g1178(.A(KEYINPUT127), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1375), .A2(new_n1376), .ZN(new_n1380));
  NAND4_X1  g1180(.A1(new_n1378), .A2(new_n1379), .A3(new_n1323), .A4(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1323), .A2(new_n1379), .ZN(new_n1382));
  OAI21_X1  g1182(.A(KEYINPUT127), .B1(new_n1319), .B2(new_n1322), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1380), .ZN(new_n1384));
  OAI211_X1 g1184(.A(new_n1382), .B(new_n1383), .C1(new_n1384), .C2(new_n1377), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1381), .A2(new_n1385), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1386), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1364), .A2(new_n1381), .A3(new_n1385), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1387), .A2(new_n1388), .ZN(G402));
endmodule


