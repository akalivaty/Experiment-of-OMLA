//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n215));
  AND3_X1   g0015(.A1(new_n214), .A2(G50), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n211), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT66), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT1), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n217), .A2(new_n227), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n212), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n246), .B1(new_n205), .B2(G20), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n248), .B1(G50), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  OR3_X1    g0059(.A1(new_n259), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT68), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(new_n263), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n206), .A2(G33), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n253), .B1(new_n254), .B2(new_n256), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n252), .B1(new_n268), .B2(new_n246), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G41), .A2(G45), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n279), .A2(new_n212), .B1(new_n280), .B2(G1), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(G226), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n288), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G1698), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n292), .B1(G222), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n283), .B1(new_n297), .B2(new_n276), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT72), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(G200), .B2(new_n298), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n271), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(G232), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G226), .B2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G97), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n306), .A2(new_n295), .B1(new_n285), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n276), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n276), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G238), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n276), .B2(new_n312), .ZN(new_n315));
  OAI211_X1 g0115(.A(KEYINPUT74), .B(new_n277), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n281), .A2(KEYINPUT73), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(G238), .A3(new_n313), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT74), .B1(new_n319), .B2(new_n277), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n310), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(new_n310), .C1(new_n317), .C2(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(new_n299), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n251), .A2(KEYINPUT70), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n249), .A2(new_n206), .A3(G1), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n246), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(G68), .C1(G1), .C2(new_n206), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT12), .B1(new_n331), .B2(G68), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G20), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(KEYINPUT12), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n250), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G50), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n337), .B1(new_n267), .B2(new_n291), .C1(new_n256), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n246), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT11), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n334), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n326), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n325), .A2(G200), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n296), .A2(G232), .ZN(new_n349));
  INV_X1    g0149(.A(G107), .ZN(new_n350));
  INV_X1    g0150(.A(G238), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n349), .B1(new_n350), .B2(new_n288), .C1(new_n351), .C2(new_n289), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n309), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n278), .B1(G244), .B2(new_n282), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G190), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n333), .B(G77), .C1(G1), .C2(new_n206), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT8), .B(G58), .Z(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n267), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n246), .B1(new_n332), .B2(new_n291), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT71), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n357), .A2(new_n365), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n353), .A2(new_n354), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G200), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n356), .A2(new_n364), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n363), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n298), .A2(new_n372), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G179), .B2(new_n298), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n269), .A2(new_n377), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(KEYINPUT69), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(KEYINPUT69), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n303), .A2(new_n348), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n322), .A2(G179), .A3(new_n324), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(new_n372), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n383), .A2(new_n384), .B1(new_n325), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n386), .ZN(new_n388));
  AOI211_X1 g0188(.A(KEYINPUT14), .B(new_n388), .C1(new_n322), .C2(new_n324), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n345), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G200), .ZN(new_n392));
  OAI211_X1 g0192(.A(G223), .B(new_n304), .C1(new_n293), .C2(new_n294), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT77), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n288), .A2(KEYINPUT77), .A3(G223), .A4(new_n304), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(G226), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n276), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n276), .A2(G232), .A3(new_n312), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n277), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT78), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT78), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n277), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n392), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n277), .A2(new_n403), .A3(new_n406), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n406), .B1(new_n277), .B2(new_n403), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n400), .B1(new_n395), .B2(new_n396), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n299), .C1(new_n276), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n286), .A2(new_n206), .A3(new_n287), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n287), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n336), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n259), .A2(new_n336), .ZN(new_n421));
  OAI21_X1  g0221(.A(G20), .B1(new_n421), .B2(new_n201), .ZN(new_n422));
  INV_X1    g0222(.A(G159), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n256), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT76), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT16), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  OAI211_X1 g0227(.A(KEYINPUT76), .B(new_n427), .C1(new_n420), .C2(new_n424), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n246), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n264), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n263), .B1(new_n258), .B2(new_n260), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n247), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n262), .A2(new_n328), .A3(new_n264), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n415), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n429), .A2(new_n435), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n372), .B1(new_n402), .B2(new_n408), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n412), .B(new_n370), .C1(new_n276), .C2(new_n413), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n246), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n425), .B2(KEYINPUT16), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n434), .B1(new_n446), .B2(new_n428), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(new_n442), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT18), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(KEYINPUT17), .A3(new_n415), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n438), .A2(new_n444), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n382), .A2(new_n391), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n445), .B(new_n251), .C1(G1), .C2(new_n285), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G97), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n328), .A2(new_n307), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT80), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n255), .A2(G77), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n350), .A2(KEYINPUT6), .A3(G97), .ZN(new_n462));
  XNOR2_X1  g0262(.A(G97), .B(G107), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n461), .B1(new_n465), .B2(new_n206), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n350), .B1(new_n418), .B2(new_n419), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n246), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT79), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(KEYINPUT79), .B(new_n246), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n205), .B(G45), .C1(new_n272), .C2(KEYINPUT5), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(new_n276), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G244), .B(new_n304), .C1(new_n293), .C2(new_n294), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT4), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n304), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n480), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n477), .B1(new_n484), .B2(new_n309), .ZN(new_n485));
  INV_X1    g0285(.A(G274), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n309), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n273), .A2(G1), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(KEYINPUT5), .C2(new_n272), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n475), .A2(KEYINPUT81), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n487), .A2(new_n473), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n485), .A2(new_n370), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n472), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(G169), .B1(new_n485), .B2(new_n492), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT82), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NOR4_X1   g0298(.A1(new_n472), .A2(new_n493), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n328), .A2(new_n350), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT25), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n454), .A2(new_n350), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n206), .B(G87), .C1(new_n293), .C2(new_n294), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT22), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n285), .A2(new_n508), .A3(G20), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n206), .B2(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n350), .A2(KEYINPUT23), .A3(G20), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT24), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT24), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n507), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n505), .B1(new_n518), .B2(new_n246), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n288), .A2(new_n304), .ZN(new_n520));
  INV_X1    g0320(.A(G250), .ZN(new_n521));
  INV_X1    g0321(.A(G294), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n520), .A2(new_n521), .B1(new_n285), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n288), .A2(G257), .A3(G1698), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n309), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(G264), .B(new_n276), .C1(new_n474), .C2(new_n475), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n492), .A3(new_n527), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n528), .A2(new_n299), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(G200), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n519), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n488), .A2(new_n486), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(new_n276), .C1(G250), .C2(new_n488), .ZN(new_n533));
  MUX2_X1   g0333(.A(G238), .B(G244), .S(G1698), .Z(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n288), .B1(G33), .B2(G116), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n535), .B2(new_n276), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n372), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G179), .B2(new_n536), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n206), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n307), .A3(new_n350), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n206), .B(G68), .C1(new_n293), .C2(new_n294), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n267), .B2(new_n307), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT83), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n445), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT83), .A4(new_n547), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n551), .B1(new_n332), .B2(new_n360), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT84), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n360), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n455), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT85), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n548), .A2(new_n549), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n246), .A3(new_n551), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n332), .A2(new_n360), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n558), .A2(KEYINPUT85), .A3(new_n555), .A4(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n539), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n455), .A2(G87), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n552), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n536), .A2(G200), .ZN(new_n565));
  INV_X1    g0365(.A(new_n536), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G190), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n531), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n485), .A2(new_n492), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n472), .B(new_n572), .C1(new_n299), .C2(new_n571), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n500), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n288), .A2(G264), .A3(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n288), .A2(G257), .A3(new_n304), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n295), .A2(G303), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n578), .A2(new_n309), .ZN(new_n579));
  OAI211_X1 g0379(.A(G270), .B(new_n276), .C1(new_n474), .C2(new_n475), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n492), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT21), .B(G169), .C1(new_n579), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n309), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n583), .A2(G179), .A3(new_n492), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n332), .A2(new_n508), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n245), .A2(new_n212), .B1(G20), .B2(new_n508), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n482), .B(new_n206), .C1(G33), .C2(new_n307), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT86), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n587), .A2(new_n588), .B1(new_n589), .B2(KEYINPUT20), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n589), .B2(KEYINPUT20), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n508), .B1(new_n205), .B2(G33), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n331), .A2(new_n445), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT20), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n587), .A2(KEYINPUT86), .A3(new_n588), .A4(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n586), .A2(new_n591), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n585), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n583), .A2(new_n492), .A3(new_n580), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(G200), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n299), .B2(new_n599), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n599), .A3(G169), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n517), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n516), .B1(new_n507), .B2(new_n513), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n246), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n504), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n296), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n276), .B1(new_n609), .B2(new_n524), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n492), .A2(new_n527), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n372), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n526), .A2(new_n370), .A3(new_n492), .A4(new_n527), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n598), .A2(new_n601), .A3(new_n604), .A4(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n453), .A2(new_n574), .A3(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n444), .A2(new_n449), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n374), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n391), .B1(new_n348), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n438), .A2(new_n450), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n303), .B1(new_n379), .B2(new_n380), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n472), .A2(new_n495), .A3(new_n493), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n562), .A4(new_n568), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT89), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n558), .A2(new_n555), .A3(new_n559), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n560), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n629), .B1(new_n633), .B2(new_n539), .ZN(new_n634));
  AOI211_X1 g0434(.A(KEYINPUT89), .B(new_n538), .C1(new_n632), .C2(new_n560), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n562), .A2(new_n568), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n470), .A2(new_n471), .ZN(new_n638));
  INV_X1    g0438(.A(new_n460), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n493), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n496), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n498), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n494), .A2(KEYINPUT82), .A3(new_n496), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n628), .B(new_n636), .C1(new_n645), .C2(new_n627), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n644), .A3(new_n573), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n597), .A2(new_n604), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT88), .B1(new_n519), .B2(new_n614), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT88), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n608), .A2(new_n615), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n647), .A2(new_n652), .A3(new_n569), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n625), .B1(new_n453), .B2(new_n654), .ZN(G369));
  NAND2_X1  g0455(.A1(new_n598), .A2(new_n604), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n601), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT92), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n250), .A2(new_n206), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT90), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT91), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  INV_X1    g0465(.A(G213), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n664), .A2(G343), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n596), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n658), .A2(KEYINPUT92), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n659), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n669), .A2(new_n648), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n608), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n531), .A3(new_n616), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n668), .A2(new_n608), .A3(new_n615), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n671), .A2(G330), .A3(new_n672), .A4(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n674), .ZN(new_n678));
  INV_X1    g0478(.A(new_n668), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n656), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n649), .A2(new_n651), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n668), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n209), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n543), .A2(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n216), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n688), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n679), .B1(new_n646), .B2(new_n653), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT93), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT93), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n697), .B(new_n679), .C1(new_n646), .C2(new_n653), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT94), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n597), .A2(KEYINPUT87), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n597), .A2(KEYINPUT87), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n604), .B(new_n616), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n574), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT26), .B1(new_n637), .B2(new_n642), .ZN(new_n706));
  INV_X1    g0506(.A(new_n637), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n497), .B2(new_n499), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n636), .B(new_n706), .C1(new_n708), .C2(KEYINPUT26), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT29), .B(new_n679), .C1(new_n705), .C2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT94), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n695), .A2(new_n711), .A3(new_n696), .A4(new_n698), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n700), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n574), .A2(new_n617), .A3(new_n668), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n528), .A2(new_n536), .ZN(new_n715));
  INV_X1    g0515(.A(new_n584), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n485), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT30), .A4(new_n485), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n566), .A2(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n571), .A2(new_n721), .A3(new_n528), .A4(new_n599), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n723), .B2(new_n668), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(G330), .B1(new_n714), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n713), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n693), .B1(new_n730), .B2(G1), .ZN(G364));
  AND2_X1   g0531(.A1(new_n671), .A2(new_n672), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n671), .A2(G330), .A3(new_n672), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n249), .A2(G20), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G45), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT95), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(KEYINPUT95), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n687), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n733), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT96), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n732), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n212), .B1(G20), .B2(new_n372), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n206), .A2(new_n370), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G200), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT97), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n299), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(G190), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G50), .A2(new_n755), .B1(new_n756), .B2(G68), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n206), .A2(G179), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G190), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G159), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT98), .B(KEYINPUT32), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n758), .A2(new_n299), .A3(G200), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n762), .A2(new_n763), .B1(new_n350), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n299), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n206), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n307), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n751), .A2(new_n759), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n288), .B1(new_n770), .B2(new_n291), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n751), .A2(G190), .A3(new_n392), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n771), .B1(G58), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n542), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n762), .B2(new_n763), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n757), .A2(new_n769), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n755), .A2(G326), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n756), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n295), .B1(new_n770), .B2(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(G329), .C2(new_n761), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  INV_X1    g0587(.A(G303), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n764), .B1(new_n775), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n767), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G294), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n779), .A2(new_n781), .A3(new_n786), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n750), .B1(new_n778), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n686), .A2(new_n295), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G355), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G116), .B2(new_n209), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n686), .A2(new_n288), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n216), .B2(new_n273), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n240), .A2(new_n273), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n746), .A2(new_n749), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n740), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n793), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n743), .B1(new_n748), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  NAND2_X1  g0607(.A1(new_n621), .A2(new_n679), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT100), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n368), .A2(new_n366), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G190), .A2(new_n355), .B1(new_n363), .B2(KEYINPUT71), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n810), .A2(new_n811), .B1(new_n363), .B2(new_n668), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n808), .B(new_n809), .C1(new_n812), .C2(new_n621), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n668), .A2(new_n363), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n373), .A2(new_n363), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n369), .A2(new_n814), .B1(new_n815), .B2(new_n371), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n374), .A2(new_n668), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT100), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n695), .A2(new_n698), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n636), .A2(new_n628), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(KEYINPUT26), .B2(new_n708), .ZN(new_n823));
  INV_X1    g0623(.A(new_n648), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n682), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n825), .A2(new_n500), .A3(new_n570), .A4(new_n573), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n668), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n819), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n740), .B1(new_n829), .B2(new_n728), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n728), .B2(new_n829), .ZN(new_n831));
  INV_X1    g0631(.A(new_n770), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n773), .A2(G143), .B1(new_n832), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(new_n755), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(new_n756), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n833), .B1(new_n834), .B2(new_n835), .C1(new_n254), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT99), .Z(new_n838));
  INV_X1    g0638(.A(KEYINPUT34), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n764), .A2(new_n336), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n295), .B(new_n842), .C1(G132), .C2(new_n761), .ZN(new_n843));
  INV_X1    g0643(.A(new_n775), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n790), .A2(G58), .B1(new_n844), .B2(G50), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n840), .A2(new_n841), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G283), .A2(new_n756), .B1(new_n755), .B2(G303), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n772), .A2(new_n522), .B1(new_n770), .B2(new_n508), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n288), .B(new_n848), .C1(G311), .C2(new_n761), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n764), .A2(new_n542), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n850), .B(new_n768), .C1(G107), .C2(new_n844), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n847), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n750), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n749), .A2(new_n744), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n741), .B(new_n853), .C1(new_n291), .C2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n745), .B2(new_n819), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n831), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  INV_X1    g0658(.A(new_n465), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n859), .A2(KEYINPUT35), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(KEYINPUT35), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n860), .A2(new_n861), .A3(G116), .A4(new_n213), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT36), .Z(new_n863));
  OAI211_X1 g0663(.A(new_n216), .B(G77), .C1(new_n259), .C2(new_n336), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n341), .A2(G68), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n205), .B(G13), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n436), .B1(new_n447), .B2(new_n448), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n664), .A2(new_n667), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n447), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n869), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n439), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n439), .A2(new_n443), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n436), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n871), .A2(new_n876), .B1(new_n451), .B2(new_n870), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT103), .B1(new_n877), .B2(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n871), .A2(new_n876), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n451), .A2(new_n870), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n881), .A2(KEYINPUT103), .A3(new_n882), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT104), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n387), .A2(new_n389), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n348), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n668), .A2(new_n345), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n390), .A2(KEYINPUT101), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT101), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n345), .C1(new_n387), .C2(new_n389), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n891), .B1(new_n346), .B2(new_n347), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n894), .A2(KEYINPUT102), .A3(new_n896), .A4(new_n897), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n893), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n817), .B1(new_n827), .B2(new_n819), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n888), .A2(new_n904), .B1(new_n619), .B2(new_n869), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n894), .ZN(new_n907));
  INV_X1    g0707(.A(new_n896), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n679), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n879), .B2(new_n880), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n877), .A2(new_n913), .A3(KEYINPUT38), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(KEYINPUT106), .B(new_n910), .C1(new_n914), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n910), .B1(new_n914), .B2(new_n916), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n909), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n906), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n700), .A2(new_n452), .A3(new_n710), .A4(new_n712), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(new_n625), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n925), .B(new_n927), .Z(new_n928));
  NAND2_X1  g0728(.A1(new_n884), .A2(new_n885), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n900), .A2(new_n901), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n892), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n885), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n726), .B1(new_n724), .B2(KEYINPUT107), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT107), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n723), .A2(new_n936), .A3(KEYINPUT31), .A4(new_n668), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n819), .B1(new_n938), .B2(new_n714), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n931), .A2(new_n933), .A3(new_n934), .A4(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n877), .A2(KEYINPUT38), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n883), .A2(KEYINPUT105), .A3(new_n944), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n945), .A2(new_n915), .A3(KEYINPUT40), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(new_n933), .A3(new_n940), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n938), .ZN(new_n949));
  INV_X1    g0749(.A(new_n714), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n452), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n948), .A2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(G330), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n928), .A2(new_n956), .B1(new_n205), .B2(new_n735), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n928), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n867), .B1(new_n957), .B2(new_n958), .ZN(G367));
  NOR2_X1   g0759(.A1(new_n798), .A2(new_n236), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n802), .B1(new_n209), .B2(new_n360), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n740), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G143), .A2(new_n755), .B1(new_n756), .B2(G159), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT110), .B(G137), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n770), .A2(new_n341), .B1(new_n760), .B2(new_n964), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n295), .B(new_n965), .C1(G150), .C2(new_n773), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n775), .A2(new_n259), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n764), .A2(new_n291), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(G68), .C2(new_n790), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n963), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n844), .A2(G116), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT46), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n288), .B1(new_n761), .B2(G317), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n773), .A2(G303), .B1(new_n832), .B2(G283), .ZN(new_n974));
  INV_X1    g0774(.A(new_n764), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n790), .A2(G107), .B1(new_n975), .B2(G97), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n522), .A2(new_n836), .B1(new_n834), .B2(new_n784), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n970), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT47), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n962), .B1(new_n980), .B2(new_n749), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n679), .A2(new_n564), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n634), .B2(new_n635), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n637), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n981), .B1(new_n984), .B2(new_n747), .ZN(new_n985));
  INV_X1    g0785(.A(new_n677), .ZN(new_n986));
  INV_X1    g0786(.A(new_n684), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n500), .B(new_n573), .C1(new_n472), .C2(new_n679), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n626), .A2(new_n668), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT108), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT108), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n684), .A2(new_n993), .A3(new_n990), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(KEYINPUT45), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n987), .A2(KEYINPUT44), .A3(new_n991), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n684), .B2(new_n990), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT45), .B1(new_n992), .B2(new_n994), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n986), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n992), .A2(new_n994), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1005), .A2(new_n677), .A3(new_n999), .A4(new_n995), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n676), .B1(new_n656), .B2(new_n679), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT109), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n681), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n1009), .B2(new_n1008), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n734), .B(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n730), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n687), .B(KEYINPUT41), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n739), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n990), .A2(new_n681), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT42), .Z(new_n1017));
  OAI21_X1  g0817(.A(new_n500), .B1(new_n991), .B2(new_n616), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n679), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1017), .A2(new_n1019), .B1(KEYINPUT43), .B2(new_n984), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n677), .A2(new_n991), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1022), .B(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n985), .B1(new_n1015), .B2(new_n1025), .ZN(G387));
  INV_X1    g0826(.A(new_n1012), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n730), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1012), .A2(new_n729), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1028), .A2(new_n272), .A3(new_n209), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n689), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n794), .A2(new_n1031), .B1(new_n350), .B2(new_n686), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n233), .A2(new_n273), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n358), .A2(new_n341), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT50), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n689), .B(new_n273), .C1(new_n336), .C2(new_n291), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n797), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1032), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n741), .B1(new_n1038), .B2(new_n802), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n676), .B2(new_n747), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n554), .A2(new_n790), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n341), .B2(new_n772), .C1(new_n336), .C2(new_n770), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G159), .B2(new_n755), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n295), .B1(new_n761), .B2(G150), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n844), .A2(G77), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n307), .C2(new_n764), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT111), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1043), .B(new_n1047), .C1(new_n266), .C2(new_n836), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n773), .A2(G317), .B1(new_n832), .B2(G303), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n834), .B2(new_n782), .C1(new_n784), .C2(new_n836), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n790), .A2(G283), .B1(new_n844), .B2(G294), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT49), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT112), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n764), .A2(new_n508), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n288), .B(new_n1059), .C1(G326), .C2(new_n761), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1057), .A2(KEYINPUT112), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1048), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1040), .B1(new_n1063), .B2(new_n749), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n1027), .B2(new_n739), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1030), .A2(new_n1065), .ZN(G393));
  NAND3_X1  g0866(.A1(new_n1002), .A2(KEYINPUT113), .A3(new_n1006), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT113), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n1069), .A3(new_n677), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n739), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n802), .B1(new_n307), .B2(new_n209), .C1(new_n798), .C2(new_n243), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n741), .B1(new_n1073), .B2(KEYINPUT114), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(KEYINPUT114), .B2(new_n1073), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n755), .A2(G150), .B1(G159), .B2(new_n773), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n836), .A2(new_n341), .ZN(new_n1078));
  INV_X1    g0878(.A(G143), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n288), .B1(new_n760), .B2(new_n1079), .C1(new_n257), .C2(new_n770), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n850), .B1(G68), .B2(new_n844), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n291), .B2(new_n767), .ZN(new_n1082));
  NOR4_X1   g0882(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n755), .A2(G317), .B1(G311), .B2(new_n773), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT52), .Z(new_n1087));
  OAI22_X1  g0887(.A1(new_n350), .A2(new_n764), .B1(new_n775), .B2(new_n787), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n295), .B1(new_n760), .B2(new_n782), .C1(new_n522), .C2(new_n770), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G116), .C2(new_n790), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1087), .B(new_n1090), .C1(new_n788), .C2(new_n836), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1084), .A2(new_n1085), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1075), .B1(new_n1092), .B2(new_n749), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n990), .B2(new_n747), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1028), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n687), .B1(new_n1028), .B2(new_n1007), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1072), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(G390));
  OAI21_X1  g0897(.A(new_n909), .B1(new_n902), .B2(new_n903), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n923), .A2(new_n1098), .A3(new_n918), .A4(new_n917), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n819), .B(new_n679), .C1(new_n705), .C2(new_n709), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n808), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n933), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1102), .A2(new_n909), .A3(new_n915), .A4(new_n945), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(G330), .B(new_n819), .C1(new_n938), .C2(new_n714), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n902), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(G330), .B(new_n819), .C1(new_n714), .C2(new_n727), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n902), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1099), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n739), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT116), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n452), .A2(G330), .A3(new_n951), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n926), .A2(new_n625), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n902), .A2(new_n1108), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n902), .B2(new_n1105), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n903), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1101), .B1(new_n902), .B2(new_n1105), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1116), .A2(new_n1117), .B1(new_n1118), .B2(new_n1109), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n1110), .A3(new_n1107), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1099), .A2(new_n1109), .A3(new_n1103), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1106), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1122), .A2(new_n1124), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(new_n1125), .A3(new_n687), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n741), .B1(new_n266), .B2(new_n854), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n964), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G128), .A2(new_n755), .B1(new_n756), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G132), .ZN(new_n1130));
  INV_X1    g0930(.A(G125), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n772), .A2(new_n1130), .B1(new_n760), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  AOI211_X1 g0933(.A(new_n295), .B(new_n1132), .C1(new_n832), .C2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n790), .A2(G159), .B1(new_n975), .B2(G50), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n775), .A2(new_n254), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1129), .A2(new_n1134), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G107), .A2(new_n756), .B1(new_n755), .B2(G283), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n772), .A2(new_n508), .B1(new_n760), .B2(new_n522), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n288), .B(new_n1140), .C1(G97), .C2(new_n832), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n776), .B(new_n842), .C1(G77), .C2(new_n790), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n920), .A2(new_n923), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1127), .B1(new_n750), .B2(new_n1144), .C1(new_n1145), .C2(new_n745), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1112), .A2(new_n1126), .A3(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1114), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1121), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n378), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n303), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n269), .A2(new_n869), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1154), .B(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n902), .A2(new_n939), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT40), .B1(new_n888), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n947), .A2(G330), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT119), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT119), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n955), .B1(new_n1158), .B2(new_n946), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n943), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1157), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1162), .B1(new_n943), .B2(new_n1163), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1154), .B(new_n1155), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(KEYINPUT121), .B(new_n925), .C1(new_n1165), .C2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1159), .A2(new_n1160), .A3(KEYINPUT119), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1167), .B1(new_n1170), .B2(new_n1166), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n924), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(new_n905), .A3(KEYINPUT121), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1161), .A2(new_n1157), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT121), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n906), .B2(new_n924), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1150), .A2(new_n1169), .A3(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1114), .B1(new_n1179), .B2(new_n1120), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT120), .B1(new_n906), .B2(new_n924), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1171), .A2(new_n1174), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT120), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1172), .B2(new_n905), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1180), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n687), .B(new_n1178), .C1(new_n1186), .C2(KEYINPUT57), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1157), .A2(new_n745), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n288), .A2(G41), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n787), .B2(new_n760), .C1(new_n350), .C2(new_n772), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1045), .B1(new_n259), .B2(new_n764), .C1(new_n336), .C2(new_n767), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n554), .C2(new_n832), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n307), .B2(new_n836), .C1(new_n508), .C2(new_n834), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT117), .Z(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1189), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G50), .B1(new_n285), .B2(new_n272), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1194), .A2(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n767), .A2(new_n254), .ZN(new_n1199));
  INV_X1    g0999(.A(G128), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n772), .A2(new_n1200), .B1(new_n770), .B2(new_n835), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(new_n844), .C2(new_n1133), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n834), .B2(new_n1131), .C1(new_n1130), .C2(new_n836), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n975), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1198), .B1(new_n1195), .B2(new_n1194), .C1(new_n1204), .C2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT118), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n750), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n1210), .B2(new_n1209), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n854), .A2(new_n341), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1188), .A2(new_n740), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1185), .A2(new_n1182), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n739), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1187), .A2(new_n1217), .ZN(G375));
  INV_X1    g1018(.A(new_n1119), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n902), .A2(new_n744), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT123), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n749), .A2(G68), .A3(new_n744), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G132), .A2(new_n755), .B1(new_n756), .B2(new_n1133), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n770), .A2(new_n254), .B1(new_n760), .B2(new_n1200), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n295), .B(new_n1224), .C1(new_n773), .C2(new_n1128), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n767), .A2(new_n341), .B1(new_n764), .B2(new_n259), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G159), .B2(new_n844), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n968), .B1(G97), .B2(new_n844), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n288), .B1(new_n773), .B2(G283), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G107), .A2(new_n832), .B1(new_n761), .B2(G303), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1041), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n508), .A2(new_n836), .B1(new_n834), .B2(new_n522), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1228), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT124), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n750), .B1(new_n1234), .B2(KEYINPUT124), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n741), .B(new_n1222), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1219), .A2(new_n739), .B1(new_n1221), .B2(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1014), .B(KEYINPUT122), .Z(new_n1239));
  OR2_X1    g1039(.A1(new_n1120), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1238), .B1(new_n1240), .B2(new_n1242), .ZN(G381));
  NAND3_X1  g1043(.A1(new_n1030), .A2(new_n806), .A3(new_n1065), .ZN(new_n1244));
  OR4_X1    g1044(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1244), .ZN(new_n1245));
  OR4_X1    g1045(.A1(G387), .A2(new_n1245), .A3(G375), .A4(G378), .ZN(G407));
  AND3_X1   g1046(.A1(new_n1112), .A2(new_n1126), .A3(new_n1146), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n666), .A2(G343), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G375), .C2(new_n1249), .ZN(G409));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1187), .A2(G378), .A3(new_n1217), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1239), .B(new_n1180), .C1(new_n1182), .C2(new_n1185), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1169), .A2(new_n1177), .A3(new_n739), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1214), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1247), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1248), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1242), .A2(KEYINPUT60), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT60), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1241), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1120), .A2(new_n688), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1258), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1238), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n857), .A2(KEYINPUT125), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n857), .A2(KEYINPUT125), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1248), .A2(G2897), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1262), .A2(KEYINPUT125), .A3(new_n857), .A4(new_n1238), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1267), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1251), .B1(new_n1257), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT127), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(KEYINPUT127), .B(new_n1251), .C1(new_n1257), .C2(new_n1271), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1257), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1257), .A2(new_n1279), .A3(new_n1276), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1274), .A2(new_n1275), .A3(new_n1278), .A4(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1022), .B(new_n1023), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n739), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n985), .A3(G390), .ZN(new_n1285));
  INV_X1    g1085(.A(G390), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(G387), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1244), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n806), .B1(new_n1030), .B2(new_n1065), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1285), .A2(new_n1287), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1281), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1251), .A3(new_n1294), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1297), .B(KEYINPUT126), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1257), .A2(new_n1271), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1257), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT63), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1277), .A2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .A4(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1296), .A2(new_n1303), .ZN(G405));
  XNOR2_X1  g1104(.A(G375), .B(G378), .ZN(new_n1305));
  OR2_X1    g1105(.A1(new_n1305), .A2(new_n1276), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1295), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1276), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1307), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


